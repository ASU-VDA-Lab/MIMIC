module fake_jpeg_20580_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_28),
.B(n_1),
.Y(n_44)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_33),
.Y(n_38)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

AO22x1_ASAP7_75t_L g34 ( 
.A1(n_19),
.A2(n_24),
.B1(n_26),
.B2(n_23),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_26),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_48),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_28),
.B1(n_15),
.B2(n_14),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_20),
.Y(n_46)
);

A2O1A1O1Ixp25_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_34),
.B(n_14),
.C(n_15),
.D(n_13),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_33),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_19),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

XOR2x2_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_35),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_45),
.C(n_34),
.Y(n_75)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_54),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_61),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_60),
.C(n_44),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_36),
.B1(n_33),
.B2(n_31),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_45),
.B1(n_48),
.B2(n_30),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_38),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_67),
.B(n_70),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_43),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_72),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_38),
.B(n_45),
.C(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_13),
.Y(n_74)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_77),
.C(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_41),
.C(n_34),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_86),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_60),
.B1(n_30),
.B2(n_32),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_91),
.B1(n_63),
.B2(n_71),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_23),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_77),
.C(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_18),
.B1(n_17),
.B2(n_26),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_42),
.B1(n_49),
.B2(n_39),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_63),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_103),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_67),
.C(n_73),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_84),
.C(n_90),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_65),
.B1(n_66),
.B2(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_98),
.B(n_99),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_91),
.C(n_81),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_85),
.B(n_90),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_18),
.C(n_17),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_88),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_110),
.C(n_111),
.Y(n_114)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_11),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_98),
.B1(n_101),
.B2(n_94),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_87),
.Y(n_111)
);

MAJx2_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_104),
.C(n_53),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_117),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_102),
.B1(n_96),
.B2(n_82),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_115),
.A2(n_116),
.B(n_55),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_112),
.B1(n_111),
.B2(n_108),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_27),
.B1(n_23),
.B2(n_55),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_2),
.C(n_3),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_119),
.B(n_9),
.Y(n_121)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_123),
.C(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_4),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_27),
.Y(n_122)
);

OAI31xp33_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_10),
.A3(n_116),
.B(n_6),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_126),
.A3(n_122),
.B1(n_5),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_127),
.B(n_128),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_114),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_130),
.A2(n_129),
.B(n_5),
.C(n_7),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_114),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_4),
.B(n_7),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_132),
.Y(n_135)
);


endmodule