module real_jpeg_25838_n_5 (n_4, n_0, n_1, n_2, n_3, n_5);

input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_5;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_6;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g8 ( 
.A1(n_1),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_8)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx8_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_3),
.A2(n_9),
.B1(n_11),
.B2(n_18),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_3),
.B(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_4),
.A2(n_8),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g5 ( 
.A(n_6),
.B(n_22),
.Y(n_5)
);

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_7),
.B(n_19),
.Y(n_6)
);

AOI21xp5_ASAP7_75t_SL g7 ( 
.A1(n_8),
.A2(n_12),
.B(n_14),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_9),
.B(n_20),
.Y(n_19)
);

OA22x2_ASAP7_75t_L g26 ( 
.A1(n_9),
.A2(n_11),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_17),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_32),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);


endmodule