module fake_jpeg_11578_n_649 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_649);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_649;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_3),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_5),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_1),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_63),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_66),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_18),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_67),
.B(n_72),
.Y(n_136)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_69),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_71),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_21),
.B(n_18),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_75),
.Y(n_175)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_77),
.A2(n_29),
.B1(n_55),
.B2(n_28),
.Y(n_150)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_85),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_86),
.Y(n_190)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

BUFx12f_ASAP7_75t_SL g88 ( 
.A(n_42),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_88),
.A2(n_40),
.B(n_49),
.Y(n_163)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_93),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_94),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_96),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_46),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_98),
.B(n_110),
.Y(n_203)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_18),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_101),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_27),
.B(n_18),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_102),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g209 ( 
.A(n_103),
.Y(n_209)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_105),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_54),
.Y(n_107)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_27),
.B(n_17),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_123),
.Y(n_144)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_33),
.B(n_16),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_21),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_111),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_21),
.Y(n_114)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_21),
.B(n_16),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_115),
.B(n_120),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_33),
.B(n_16),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_30),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_125),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_126),
.Y(n_214)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_48),
.Y(n_128)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_48),
.Y(n_129)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_129),
.Y(n_187)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_42),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_19),
.B1(n_50),
.B2(n_57),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_132),
.A2(n_156),
.B1(n_159),
.B2(n_168),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_63),
.B(n_49),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_149),
.B(n_123),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_150),
.A2(n_158),
.B1(n_160),
.B2(n_188),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_70),
.A2(n_19),
.B1(n_50),
.B2(n_57),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g158 ( 
.A1(n_77),
.A2(n_79),
.B1(n_103),
.B2(n_95),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_65),
.A2(n_39),
.B1(n_44),
.B2(n_30),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_67),
.A2(n_50),
.B1(n_19),
.B2(n_40),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_163),
.B(n_127),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_72),
.B(n_28),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_167),
.B(n_202),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_88),
.A2(n_39),
.B1(n_44),
.B2(n_57),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_80),
.A2(n_39),
.B1(n_44),
.B2(n_54),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_177),
.A2(n_179),
.B1(n_216),
.B2(n_102),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_69),
.A2(n_48),
.B1(n_41),
.B2(n_36),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_83),
.A2(n_55),
.B1(n_45),
.B2(n_43),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g289 ( 
.A1(n_180),
.A2(n_192),
.B1(n_207),
.B2(n_208),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_L g188 ( 
.A1(n_71),
.A2(n_45),
.B1(n_43),
.B2(n_20),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_73),
.A2(n_20),
.B1(n_38),
.B2(n_29),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_64),
.B(n_38),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_85),
.A2(n_86),
.B1(n_94),
.B2(n_105),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_204),
.A2(n_119),
.B1(n_126),
.B2(n_124),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_112),
.A2(n_35),
.B1(n_31),
.B2(n_36),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_115),
.A2(n_35),
.B1(n_31),
.B2(n_34),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_111),
.A2(n_41),
.B1(n_23),
.B2(n_34),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_93),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_107),
.Y(n_213)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_92),
.A2(n_23),
.B1(n_15),
.B2(n_14),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_217),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_218),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

INVx5_ASAP7_75t_L g353 ( 
.A(n_219),
.Y(n_353)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_221),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_222),
.Y(n_309)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_224),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_203),
.B(n_113),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_225),
.B(n_237),
.Y(n_300)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_170),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_227),
.Y(n_318)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_228),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_134),
.B(n_130),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_229),
.B(n_231),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_183),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_232),
.B(n_242),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_233),
.Y(n_305)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_234),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_133),
.B(n_129),
.Y(n_237)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_165),
.Y(n_238)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_238),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_157),
.Y(n_239)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_178),
.B(n_128),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_240),
.B(n_244),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_241),
.Y(n_324)
);

AND2x4_ASAP7_75t_SL g242 ( 
.A(n_136),
.B(n_66),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_243),
.B(n_259),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_144),
.B(n_123),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_245),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_178),
.B(n_13),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_246),
.B(n_254),
.Y(n_347)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_248),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_249),
.A2(n_268),
.B1(n_279),
.B2(n_286),
.Y(n_312)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_250),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_163),
.A2(n_122),
.B1(n_114),
.B2(n_131),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_251),
.Y(n_327)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_169),
.Y(n_252)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_252),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_165),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_253),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_141),
.B(n_15),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_182),
.Y(n_255)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_255),
.Y(n_321)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_183),
.Y(n_256)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_256),
.Y(n_330)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_173),
.Y(n_257)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_257),
.Y(n_322)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_258),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_183),
.Y(n_259)
);

INVx3_ASAP7_75t_SL g260 ( 
.A(n_142),
.Y(n_260)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_260),
.Y(n_331)
);

NOR2x1_ASAP7_75t_L g261 ( 
.A(n_136),
.B(n_149),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_261),
.A2(n_285),
.B(n_292),
.Y(n_340)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_187),
.Y(n_262)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_262),
.Y(n_336)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_263),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_143),
.B(n_14),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_264),
.B(n_265),
.Y(n_338)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_137),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_139),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_266),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_145),
.B(n_0),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_288),
.C(n_185),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_180),
.A2(n_116),
.B1(n_37),
.B2(n_14),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_172),
.Y(n_269)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_269),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_175),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_274),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_146),
.B(n_13),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_147),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_180),
.B(n_13),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_273),
.B(n_275),
.Y(n_316)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_151),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_188),
.B(n_12),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_192),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_277),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_146),
.B(n_12),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_168),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_278),
.B(n_280),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_158),
.A2(n_37),
.B1(n_1),
.B2(n_2),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_186),
.B(n_0),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_152),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_281),
.B(n_283),
.Y(n_351)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_195),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_282),
.B(n_284),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_164),
.B(n_2),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_140),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_176),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_148),
.A2(n_37),
.B1(n_3),
.B2(n_5),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_142),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g315 ( 
.A(n_287),
.B(n_185),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_212),
.B(n_196),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_138),
.B(n_2),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_216),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_166),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_291),
.A2(n_200),
.B(n_193),
.Y(n_326)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_155),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_232),
.A2(n_179),
.B(n_177),
.C(n_159),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_297),
.B(n_328),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_235),
.A2(n_204),
.B1(n_205),
.B2(n_140),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_301),
.A2(n_304),
.B1(n_311),
.B2(n_333),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_303),
.B(n_239),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_263),
.A2(n_171),
.B1(n_161),
.B2(n_190),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_242),
.B(n_232),
.C(n_288),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_308),
.B(n_10),
.C(n_8),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_278),
.A2(n_171),
.B1(n_161),
.B2(n_190),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_314),
.B(n_303),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_315),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_223),
.A2(n_156),
.B1(n_132),
.B2(n_194),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_320),
.A2(n_341),
.B1(n_342),
.B2(n_287),
.Y(n_370)
);

AOI32xp33_ASAP7_75t_L g325 ( 
.A1(n_242),
.A2(n_174),
.A3(n_198),
.B1(n_135),
.B2(n_215),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_325),
.A2(n_298),
.B(n_305),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_326),
.A2(n_270),
.B(n_218),
.Y(n_373)
);

A2O1A1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_261),
.A2(n_209),
.B(n_184),
.C(n_154),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_223),
.A2(n_247),
.B1(n_289),
.B2(n_249),
.Y(n_333)
);

OA22x2_ASAP7_75t_L g337 ( 
.A1(n_289),
.A2(n_209),
.B1(n_194),
.B2(n_37),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_269),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_289),
.A2(n_37),
.B1(n_6),
.B2(n_7),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_289),
.A2(n_229),
.B1(n_236),
.B2(n_266),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_267),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_343),
.A2(n_222),
.B1(n_253),
.B2(n_291),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_309),
.Y(n_354)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_354),
.Y(n_403)
);

O2A1O1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_297),
.A2(n_288),
.B(n_230),
.C(n_267),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_355),
.A2(n_313),
.B(n_346),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_349),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_356),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_357),
.B(n_374),
.Y(n_409)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_306),
.Y(n_358)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_358),
.Y(n_406)
);

OAI22x1_ASAP7_75t_SL g359 ( 
.A1(n_333),
.A2(n_260),
.B1(n_234),
.B2(n_227),
.Y(n_359)
);

AOI22x1_ASAP7_75t_L g423 ( 
.A1(n_359),
.A2(n_376),
.B1(n_339),
.B2(n_302),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_300),
.B(n_220),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_360),
.B(n_378),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_256),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_361),
.B(n_399),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_301),
.A2(n_265),
.B1(n_274),
.B2(n_272),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_362),
.A2(n_365),
.B1(n_368),
.B2(n_375),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_317),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_364),
.B(n_385),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_324),
.A2(n_284),
.B1(n_217),
.B2(n_250),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_309),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_366),
.Y(n_428)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_349),
.Y(n_367)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_324),
.A2(n_258),
.B1(n_238),
.B2(n_226),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_370),
.A2(n_371),
.B1(n_377),
.B2(n_389),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_341),
.A2(n_312),
.B1(n_334),
.B2(n_314),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_373),
.A2(n_396),
.B(n_352),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_334),
.A2(n_228),
.B1(n_245),
.B2(n_224),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_323),
.A2(n_316),
.B1(n_337),
.B2(n_350),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_248),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_379),
.A2(n_382),
.B1(n_395),
.B2(n_387),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_327),
.A2(n_282),
.B(n_221),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_380),
.A2(n_298),
.B(n_353),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_8),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_381),
.B(n_386),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_316),
.A2(n_252),
.B1(n_219),
.B2(n_10),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_319),
.C(n_352),
.Y(n_424)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_307),
.Y(n_384)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_295),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_8),
.Y(n_386)
);

AO22x2_ASAP7_75t_L g388 ( 
.A1(n_337),
.A2(n_9),
.B1(n_328),
.B2(n_323),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_390),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_337),
.A2(n_9),
.B1(n_327),
.B2(n_294),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_347),
.B(n_338),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_338),
.B(n_340),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_391),
.B(n_401),
.Y(n_425)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_329),
.Y(n_392)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_392),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_294),
.A2(n_308),
.B1(n_338),
.B2(n_315),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_393),
.A2(n_394),
.B1(n_397),
.B2(n_387),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_294),
.A2(n_315),
.B1(n_340),
.B2(n_311),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_304),
.A2(n_335),
.B1(n_326),
.B2(n_343),
.Y(n_395)
);

OAI21xp33_ASAP7_75t_L g396 ( 
.A1(n_299),
.A2(n_344),
.B(n_331),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_322),
.A2(n_336),
.B1(n_321),
.B2(n_306),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_305),
.B(n_318),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_398),
.B(n_400),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_296),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_313),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_402),
.A2(n_376),
.B(n_388),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_357),
.B(n_318),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_404),
.B(n_430),
.C(n_383),
.Y(n_452)
);

OAI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_361),
.A2(n_330),
.B1(n_348),
.B2(n_310),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_407),
.A2(n_419),
.B1(n_439),
.B2(n_359),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_SL g466 ( 
.A(n_411),
.B(n_438),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_374),
.B(n_319),
.Y(n_413)
);

XOR2x2_ASAP7_75t_L g460 ( 
.A(n_413),
.B(n_376),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_397),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_414),
.B(n_415),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_356),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_418),
.A2(n_380),
.B(n_373),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_371),
.A2(n_293),
.B1(n_332),
.B2(n_346),
.Y(n_419)
);

OA22x2_ASAP7_75t_L g465 ( 
.A1(n_423),
.A2(n_414),
.B1(n_420),
.B2(n_405),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_424),
.B(n_413),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_396),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_426),
.B(n_429),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_398),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_393),
.B(n_302),
.C(n_310),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_367),
.B(n_339),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_401),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_381),
.B(n_330),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_433),
.B(n_440),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_435),
.A2(n_442),
.B1(n_408),
.B2(n_411),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_437),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_372),
.A2(n_296),
.B(n_353),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_370),
.A2(n_293),
.B1(n_332),
.B2(n_361),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_386),
.B(n_390),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_378),
.B(n_360),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_441),
.B(n_442),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_391),
.Y(n_442)
);

OAI21xp33_ASAP7_75t_L g443 ( 
.A1(n_410),
.A2(n_355),
.B(n_372),
.Y(n_443)
);

MAJx2_ASAP7_75t_L g506 ( 
.A(n_443),
.B(n_444),
.C(n_424),
.Y(n_506)
);

OAI21xp33_ASAP7_75t_L g444 ( 
.A1(n_410),
.A2(n_355),
.B(n_399),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_445),
.B(n_474),
.C(n_476),
.Y(n_492)
);

AOI322xp5_ASAP7_75t_L g446 ( 
.A1(n_427),
.A2(n_363),
.A3(n_395),
.B1(n_388),
.B2(n_377),
.C1(n_359),
.C2(n_382),
.Y(n_446)
);

OAI31xp33_ASAP7_75t_L g491 ( 
.A1(n_446),
.A2(n_448),
.A3(n_455),
.B(n_426),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_435),
.A2(n_389),
.B1(n_394),
.B2(n_388),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_449),
.A2(n_456),
.B1(n_461),
.B2(n_427),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_421),
.B(n_388),
.Y(n_450)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_450),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_431),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_451),
.B(n_458),
.Y(n_485)
);

XNOR2x1_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_430),
.Y(n_482)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_416),
.Y(n_453)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_453),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_454),
.A2(n_425),
.B1(n_420),
.B2(n_438),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_421),
.A2(n_388),
.B1(n_363),
.B2(n_376),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_409),
.B(n_383),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_457),
.B(n_477),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_434),
.Y(n_458)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_459),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_460),
.B(n_437),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_422),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_462),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_418),
.B(n_411),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_463),
.Y(n_494)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_416),
.Y(n_464)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_464),
.Y(n_509)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_465),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_405),
.B(n_375),
.Y(n_467)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_467),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_422),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_468),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_415),
.B(n_392),
.Y(n_470)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_470),
.Y(n_511)
);

INVxp33_ASAP7_75t_L g471 ( 
.A(n_434),
.Y(n_471)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_471),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_408),
.B(n_384),
.Y(n_473)
);

XOR2x1_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_479),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_409),
.B(n_404),
.C(n_413),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_409),
.B(n_404),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_440),
.B(n_362),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_429),
.B(n_412),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_475),
.A2(n_450),
.B1(n_472),
.B2(n_454),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_480),
.A2(n_484),
.B1(n_499),
.B2(n_501),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_481),
.A2(n_488),
.B1(n_478),
.B2(n_447),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_482),
.B(n_512),
.C(n_460),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_487),
.B(n_498),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_456),
.A2(n_439),
.B1(n_419),
.B2(n_438),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_458),
.A2(n_462),
.B1(n_468),
.B2(n_432),
.Y(n_490)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_490),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_491),
.A2(n_466),
.B(n_463),
.Y(n_520)
);

XNOR2x2_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_425),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_506),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_476),
.B(n_430),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_472),
.A2(n_402),
.B1(n_423),
.B2(n_433),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_470),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_508),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_451),
.A2(n_423),
.B1(n_432),
.B2(n_441),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_465),
.Y(n_505)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_505),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_445),
.B(n_424),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_455),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_473),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_452),
.B(n_412),
.C(n_417),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_453),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_513),
.B(n_406),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_447),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_515),
.B(n_530),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_499),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_517),
.B(n_536),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_520),
.A2(n_529),
.B(n_494),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_521),
.A2(n_525),
.B1(n_543),
.B2(n_489),
.Y(n_552)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_485),
.Y(n_523)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_523),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_504),
.B(n_459),
.Y(n_524)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_524),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_481),
.A2(n_479),
.B1(n_448),
.B2(n_461),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_482),
.B(n_457),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_526),
.B(n_532),
.Y(n_553)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_485),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_527),
.B(n_528),
.Y(n_564)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_501),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_491),
.A2(n_466),
.B(n_463),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_469),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_492),
.B(n_478),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_533),
.B(n_541),
.C(n_406),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_534),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_480),
.A2(n_449),
.B1(n_460),
.B2(n_446),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_535),
.A2(n_497),
.B1(n_493),
.B2(n_511),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_502),
.Y(n_536)
);

XOR2x2_ASAP7_75t_L g537 ( 
.A(n_495),
.B(n_477),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_537),
.B(n_539),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_SL g546 ( 
.A(n_538),
.B(n_495),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_492),
.B(n_469),
.Y(n_539)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_488),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_540),
.B(n_542),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_507),
.B(n_465),
.C(n_464),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_513),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_493),
.A2(n_465),
.B1(n_467),
.B2(n_423),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_506),
.B(n_498),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_544),
.B(n_496),
.Y(n_559)
);

XNOR2x1_ASAP7_75t_L g545 ( 
.A(n_538),
.B(n_487),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_545),
.B(n_546),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_548),
.B(n_559),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_520),
.A2(n_494),
.B(n_505),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_549),
.A2(n_563),
.B(n_569),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_519),
.A2(n_510),
.B1(n_489),
.B2(n_483),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_551),
.B(n_555),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_552),
.A2(n_561),
.B1(n_543),
.B2(n_536),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_535),
.A2(n_522),
.B1(n_517),
.B2(n_516),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_529),
.A2(n_483),
.B(n_511),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_557),
.B(n_365),
.Y(n_587)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_560),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_521),
.A2(n_510),
.B1(n_465),
.B2(n_486),
.Y(n_561)
);

A2O1A1Ixp33_ASAP7_75t_SL g563 ( 
.A1(n_531),
.A2(n_486),
.B(n_407),
.C(n_509),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_544),
.B(n_417),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_565),
.B(n_566),
.Y(n_575)
);

A2O1A1Ixp33_ASAP7_75t_L g568 ( 
.A1(n_524),
.A2(n_541),
.B(n_522),
.C(n_525),
.Y(n_568)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_568),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_531),
.A2(n_436),
.B(n_428),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_556),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_571),
.B(n_573),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_547),
.B(n_539),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_566),
.B(n_532),
.C(n_533),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_577),
.B(n_581),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_549),
.A2(n_556),
.B(n_561),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_578),
.A2(n_584),
.B(n_587),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_579),
.A2(n_588),
.B1(n_550),
.B2(n_563),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_547),
.B(n_358),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_553),
.B(n_526),
.C(n_518),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_582),
.B(n_583),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_553),
.B(n_518),
.C(n_514),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g584 ( 
.A1(n_548),
.A2(n_514),
.B(n_537),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_567),
.Y(n_585)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_585),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_564),
.B(n_354),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_586),
.B(n_354),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_552),
.A2(n_403),
.B1(n_366),
.B2(n_369),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_565),
.B(n_554),
.C(n_545),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_590),
.B(n_554),
.C(n_559),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_575),
.B(n_577),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_591),
.B(n_595),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_592),
.B(n_605),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_580),
.B(n_558),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_596),
.B(n_598),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_576),
.A2(n_567),
.B1(n_558),
.B2(n_550),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_575),
.B(n_562),
.C(n_560),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_599),
.B(n_602),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_SL g601 ( 
.A(n_589),
.B(n_546),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_SL g618 ( 
.A(n_601),
.B(n_608),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_576),
.B(n_562),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_604),
.A2(n_563),
.B1(n_571),
.B2(n_588),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_572),
.B(n_557),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_590),
.B(n_563),
.C(n_568),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_606),
.B(n_570),
.C(n_578),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_572),
.B(n_579),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_607),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_570),
.B(n_569),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_610),
.B(n_611),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_594),
.B(n_574),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_591),
.B(n_582),
.C(n_583),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_613),
.B(n_615),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_600),
.A2(n_593),
.B(n_608),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_606),
.B(n_574),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_616),
.B(n_592),
.C(n_601),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_600),
.A2(n_608),
.B(n_585),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_617),
.B(n_622),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_621),
.B(n_604),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_599),
.B(n_589),
.C(n_563),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g635 ( 
.A1(n_623),
.A2(n_631),
.B1(n_610),
.B2(n_622),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_620),
.B(n_603),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_625),
.A2(n_630),
.B(n_632),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_614),
.B(n_597),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_628),
.B(n_629),
.Y(n_637)
);

NOR2xp67_ASAP7_75t_L g630 ( 
.A(n_611),
.B(n_584),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_613),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_609),
.B(n_619),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_626),
.B(n_615),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_634),
.B(n_635),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_627),
.B(n_616),
.C(n_617),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_636),
.A2(n_638),
.B(n_618),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_624),
.B(n_621),
.C(n_618),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_625),
.B(n_612),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_639),
.B(n_623),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_641),
.A2(n_643),
.B(n_636),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_642),
.A2(n_637),
.B(n_638),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_633),
.A2(n_403),
.B(n_369),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_644),
.B(n_645),
.C(n_634),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_639),
.C(n_640),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_368),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_648),
.A2(n_366),
.B(n_379),
.Y(n_649)
);


endmodule