module fake_jpeg_28933_n_249 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_13),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_35),
.B(n_44),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g72 ( 
.A(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_37),
.B(n_26),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_17),
.C(n_19),
.Y(n_48)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_41),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_42),
.A2(n_31),
.B1(n_27),
.B2(n_24),
.Y(n_77)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_15),
.B(n_5),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_48),
.B(n_73),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_28),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_32),
.Y(n_92)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_52),
.Y(n_119)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_61),
.Y(n_105)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_69),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_37),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_79),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_16),
.B1(n_31),
.B2(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_29),
.B1(n_66),
.B2(n_68),
.Y(n_104)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_36),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_36),
.B(n_24),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_32),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g116 ( 
.A(n_83),
.B(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_45),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_35),
.B(n_21),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_88),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_37),
.B(n_29),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_35),
.B(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_90),
.Y(n_113)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_91),
.B(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_49),
.B(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_107),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_87),
.C(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_110),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_85),
.B1(n_75),
.B2(n_55),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_32),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_117),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_25),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_21),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_120),
.B(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_71),
.B1(n_68),
.B2(n_50),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_124),
.A2(n_128),
.B1(n_138),
.B2(n_142),
.Y(n_171)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_50),
.B1(n_25),
.B2(n_22),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_98),
.B(n_25),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_32),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_139),
.Y(n_154)
);

OAI21x1_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_116),
.B(n_94),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_147),
.Y(n_153)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_23),
.B(n_57),
.C(n_84),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_137),
.A2(n_106),
.B(n_76),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_60),
.B1(n_55),
.B2(n_65),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_23),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_112),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_141),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_65),
.B1(n_59),
.B2(n_51),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_51),
.B1(n_57),
.B2(n_23),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_23),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_25),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_104),
.A2(n_23),
.B1(n_22),
.B2(n_82),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_76),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_102),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_121),
.C(n_127),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_142),
.B1(n_126),
.B2(n_137),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_113),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_158),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_107),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_160),
.B(n_161),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_119),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_119),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_169),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_116),
.B(n_110),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

BUFx12_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_99),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_174),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_123),
.B(n_94),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_175),
.A2(n_160),
.B(n_162),
.Y(n_185)
);

OAI22x1_ASAP7_75t_SL g176 ( 
.A1(n_155),
.A2(n_144),
.B1(n_128),
.B2(n_129),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_193),
.B1(n_173),
.B2(n_166),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_129),
.A3(n_133),
.B1(n_124),
.B2(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_181),
.B1(n_188),
.B2(n_174),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_136),
.B1(n_132),
.B2(n_143),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_153),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_183),
.B(n_22),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_186),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_185),
.B(n_192),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_125),
.C(n_106),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_170),
.B1(n_159),
.B2(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_190),
.Y(n_197)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_117),
.B(n_115),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_101),
.C(n_115),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_101),
.B1(n_22),
.B2(n_115),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_198),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_168),
.B(n_159),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_207),
.B(n_209),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_200),
.B1(n_190),
.B2(n_177),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_179),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_164),
.B1(n_157),
.B2(n_172),
.Y(n_200)
);

OAI322xp33_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_154),
.A3(n_164),
.B1(n_157),
.B2(n_172),
.C1(n_150),
.C2(n_166),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_187),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_203),
.Y(n_220)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_167),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_194),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_169),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_210),
.B(n_211),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_186),
.C(n_184),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_219),
.C(n_169),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_197),
.B1(n_195),
.B2(n_205),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_192),
.C(n_185),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_226),
.B1(n_220),
.B2(n_213),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_212),
.A2(n_197),
.B(n_199),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_210),
.Y(n_231)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_203),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_228),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_200),
.B1(n_206),
.B2(n_169),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_224),
.C(n_222),
.Y(n_234)
);

NOR3xp33_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_6),
.C(n_7),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_217),
.B(n_216),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_232),
.Y(n_238)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_231),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_223),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_226),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_235),
.C(n_221),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_221),
.A2(n_220),
.B(n_211),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_6),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_240),
.Y(n_242)
);

AOI31xp67_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_213),
.A3(n_7),
.B(n_8),
.Y(n_240)
);

AOI21x1_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_234),
.B(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_232),
.C(n_8),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_243),
.B(n_244),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_242),
.C(n_8),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_246),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_6),
.Y(n_249)
);


endmodule