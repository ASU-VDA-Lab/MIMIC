module fake_netlist_6_3664_n_886 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_886);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_886;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_796;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_386;
wire n_201;
wire n_249;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

BUFx2_ASAP7_75t_L g201 ( 
.A(n_15),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_15),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_109),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_63),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_140),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_193),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_28),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_196),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_93),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_9),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_53),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_58),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_101),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_29),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_130),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_111),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_195),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_164),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_65),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_143),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_16),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_110),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_70),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_6),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_117),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_52),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_151),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_38),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_L g235 ( 
.A(n_35),
.B(n_121),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_190),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_112),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_32),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_181),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_5),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_20),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_45),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_167),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_98),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_44),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_136),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_34),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_152),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_126),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_128),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_80),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_6),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_142),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_188),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_36),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_165),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_55),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_137),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_156),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_166),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_177),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_174),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_89),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_10),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_182),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_27),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_5),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_123),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_41),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_106),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_16),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_157),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_77),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_79),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_122),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_14),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_40),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_57),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_94),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_0),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_213),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_0),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_213),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_210),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_213),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_206),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_210),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_202),
.Y(n_288)
);

CKINVDCx6p67_ASAP7_75t_R g289 ( 
.A(n_229),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_202),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_206),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_206),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_202),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_206),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_204),
.Y(n_295)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_18),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_217),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_226),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_205),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_201),
.B(n_1),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_217),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_240),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_217),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_203),
.Y(n_304)
);

BUFx12f_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_252),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_207),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_224),
.B(n_242),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_208),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_215),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_269),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_220),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_244),
.B(n_2),
.Y(n_314)
);

BUFx12f_ASAP7_75t_L g315 ( 
.A(n_271),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_230),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_232),
.Y(n_317)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_243),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_234),
.B(n_3),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_276),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_206),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_231),
.B(n_4),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_261),
.B(n_4),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_245),
.B(n_256),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_257),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_258),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_260),
.Y(n_327)
);

AND2x4_ASAP7_75t_L g328 ( 
.A(n_262),
.B(n_7),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_219),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_329)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_211),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_221),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_310),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_304),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_305),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_315),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_320),
.Y(n_338)
);

NOR2x1p5_ASAP7_75t_L g339 ( 
.A(n_284),
.B(n_209),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_281),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_R g341 ( 
.A(n_330),
.B(n_266),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_331),
.Y(n_342)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_330),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_R g344 ( 
.A(n_330),
.B(n_278),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_283),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_288),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_289),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_284),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_318),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_287),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_287),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_R g352 ( 
.A(n_330),
.B(n_212),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_318),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_288),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_318),
.B(n_293),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_318),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_295),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_R g359 ( 
.A(n_323),
.B(n_214),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_295),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_299),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_299),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_324),
.Y(n_363)
);

INVxp33_ASAP7_75t_L g364 ( 
.A(n_300),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_285),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_290),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_R g367 ( 
.A(n_323),
.B(n_216),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_290),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_290),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_307),
.Y(n_370)
);

NAND2xp33_ASAP7_75t_R g371 ( 
.A(n_314),
.B(n_8),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_307),
.Y(n_372)
);

NOR2x1p5_ASAP7_75t_L g373 ( 
.A(n_314),
.B(n_218),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_317),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_317),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_322),
.Y(n_376)
);

NAND2xp33_ASAP7_75t_R g377 ( 
.A(n_280),
.B(n_10),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_312),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_312),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_322),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_297),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_312),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_297),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_297),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_301),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_301),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_280),
.B(n_265),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_346),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_308),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_366),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_368),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_383),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_363),
.B(n_319),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_384),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_308),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_354),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_354),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_364),
.B(n_319),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

NOR3xp33_ASAP7_75t_L g401 ( 
.A(n_338),
.B(n_302),
.C(n_282),
.Y(n_401)
);

OAI221xp5_ASAP7_75t_L g402 ( 
.A1(n_377),
.A2(n_282),
.B1(n_324),
.B2(n_302),
.C(n_311),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_359),
.B(n_328),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_293),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_360),
.B(n_296),
.Y(n_405)
);

NOR3xp33_ASAP7_75t_L g406 ( 
.A(n_338),
.B(n_329),
.C(n_274),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_367),
.B(n_328),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_372),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_354),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_286),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_291),
.Y(n_412)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_358),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_385),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_361),
.B(n_222),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_382),
.B(n_313),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_354),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

INVx8_ASAP7_75t_L g420 ( 
.A(n_349),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_362),
.B(n_296),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_370),
.B(n_223),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_374),
.B(n_225),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_345),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_365),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_296),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_L g427 ( 
.A(n_373),
.B(n_296),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_333),
.B(n_316),
.Y(n_428)
);

OR2x6_ASAP7_75t_L g429 ( 
.A(n_339),
.B(n_298),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_356),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_348),
.Y(n_431)
);

INVxp33_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_343),
.B(n_301),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_344),
.B(n_227),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_350),
.B(n_228),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_376),
.B(n_235),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_353),
.B(n_303),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_357),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_SL g440 ( 
.A(n_377),
.B(n_233),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_L g441 ( 
.A(n_335),
.B(n_206),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_351),
.B(n_236),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_380),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_334),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_352),
.B(n_292),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_342),
.Y(n_446)
);

NOR3xp33_ASAP7_75t_L g447 ( 
.A(n_347),
.B(n_329),
.C(n_309),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_334),
.B(n_294),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_336),
.B(n_237),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_337),
.B(n_238),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_371),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_371),
.Y(n_452)
);

INVx8_ASAP7_75t_L g453 ( 
.A(n_349),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_346),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_346),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_346),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_363),
.B(n_303),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_399),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_306),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_409),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_389),
.B(n_457),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_425),
.Y(n_462)
);

NOR2x1p5_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_239),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_390),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_452),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_391),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_443),
.Y(n_467)
);

AND2x6_ASAP7_75t_SL g468 ( 
.A(n_429),
.B(n_272),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_411),
.B(n_273),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_420),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_411),
.B(n_279),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_SL g472 ( 
.A(n_437),
.B(n_246),
.C(n_241),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_403),
.A2(n_270),
.B1(n_248),
.B2(n_249),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_393),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_454),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_412),
.B(n_332),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_429),
.B(n_332),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_394),
.B(n_247),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_437),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_444),
.B(n_253),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_402),
.A2(n_275),
.B1(n_255),
.B2(n_259),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_SL g482 ( 
.A1(n_394),
.A2(n_254),
.B1(n_268),
.B2(n_277),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_412),
.B(n_325),
.Y(n_483)
);

BUFx8_ASAP7_75t_L g484 ( 
.A(n_431),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_430),
.B(n_325),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_439),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_429),
.B(n_325),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_388),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_418),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_448),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_392),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_401),
.A2(n_321),
.B1(n_326),
.B2(n_327),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_395),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_419),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_438),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_455),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_420),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_408),
.B(n_326),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_446),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_419),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_432),
.B(n_326),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_419),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_396),
.B(n_327),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_456),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_440),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_420),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_428),
.B(n_327),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_439),
.B(n_303),
.Y(n_509)
);

OR2x4_ASAP7_75t_L g510 ( 
.A(n_416),
.B(n_11),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_439),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_453),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_413),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_445),
.B(n_12),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_414),
.B(n_19),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_445),
.B(n_21),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_397),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_427),
.A2(n_115),
.B1(n_199),
.B2(n_198),
.Y(n_519)
);

AND2x2_ASAP7_75t_SL g520 ( 
.A(n_406),
.B(n_13),
.Y(n_520)
);

A2O1A1Ixp33_ASAP7_75t_L g521 ( 
.A1(n_405),
.A2(n_14),
.B(n_17),
.C(n_22),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_441),
.A2(n_116),
.B1(n_23),
.B2(n_24),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_404),
.B(n_25),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_398),
.Y(n_524)
);

NOR2x1p5_ASAP7_75t_L g525 ( 
.A(n_421),
.B(n_17),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_453),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_410),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_415),
.B(n_26),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_447),
.B(n_30),
.Y(n_529)
);

AO21x1_ASAP7_75t_L g530 ( 
.A1(n_478),
.A2(n_528),
.B(n_517),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_458),
.B(n_436),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_461),
.A2(n_426),
.B(n_433),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_465),
.A2(n_423),
.B1(n_422),
.B2(n_442),
.Y(n_533)
);

INVx6_ASAP7_75t_SL g534 ( 
.A(n_487),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_490),
.B(n_433),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_483),
.A2(n_434),
.B(n_435),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_486),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_479),
.B(n_449),
.Y(n_538)
);

A2O1A1Ixp33_ASAP7_75t_L g539 ( 
.A1(n_508),
.A2(n_450),
.B(n_417),
.C(n_453),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_476),
.A2(n_31),
.B(n_33),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_511),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_523),
.A2(n_37),
.B(n_39),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_459),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_498),
.A2(n_42),
.B(n_43),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_495),
.A2(n_46),
.B(n_47),
.Y(n_545)
);

BUFx4f_ASAP7_75t_SL g546 ( 
.A(n_506),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_494),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_494),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_505),
.B(n_48),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_499),
.B(n_49),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_485),
.A2(n_50),
.B(n_51),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_526),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_459),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_469),
.B(n_54),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_471),
.A2(n_56),
.B(n_59),
.Y(n_555)
);

INVx8_ASAP7_75t_L g556 ( 
.A(n_487),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_467),
.B(n_60),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_524),
.Y(n_558)
);

OA22x2_ASAP7_75t_L g559 ( 
.A1(n_514),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_460),
.B(n_66),
.Y(n_560)
);

A2O1A1Ixp33_ASAP7_75t_L g561 ( 
.A1(n_501),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_503),
.B(n_71),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_481),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_529),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_494),
.B(n_81),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_500),
.B(n_82),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_500),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_477),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_529),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_477),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_500),
.B(n_90),
.Y(n_571)
);

A2O1A1Ixp33_ASAP7_75t_L g572 ( 
.A1(n_515),
.A2(n_91),
.B(n_92),
.C(n_95),
.Y(n_572)
);

NOR2x1_ASAP7_75t_SL g573 ( 
.A(n_502),
.B(n_96),
.Y(n_573)
);

OAI21xp33_ASAP7_75t_SL g574 ( 
.A1(n_507),
.A2(n_97),
.B(n_99),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_502),
.B(n_100),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_488),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_513),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_463),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_578)
);

BUFx12f_ASAP7_75t_L g579 ( 
.A(n_470),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_502),
.B(n_105),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_510),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_489),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_462),
.A2(n_107),
.B(n_108),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_464),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_482),
.B(n_113),
.Y(n_585)
);

NOR3xp33_ASAP7_75t_SL g586 ( 
.A(n_472),
.B(n_118),
.C(n_119),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_466),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_516),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_480),
.B(n_120),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_534),
.Y(n_590)
);

AO21x2_ASAP7_75t_L g591 ( 
.A1(n_530),
.A2(n_532),
.B(n_536),
.Y(n_591)
);

CKINVDCx11_ASAP7_75t_R g592 ( 
.A(n_579),
.Y(n_592)
);

BUFx2_ASAP7_75t_SL g593 ( 
.A(n_537),
.Y(n_593)
);

AOI21x1_ASAP7_75t_L g594 ( 
.A1(n_562),
.A2(n_474),
.B(n_475),
.Y(n_594)
);

OAI21x1_ASAP7_75t_L g595 ( 
.A1(n_565),
.A2(n_527),
.B(n_518),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_576),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g597 ( 
.A(n_552),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_558),
.Y(n_598)
);

AOI22x1_ASAP7_75t_L g599 ( 
.A1(n_589),
.A2(n_525),
.B1(n_491),
.B2(n_493),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_534),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_584),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_588),
.B(n_496),
.Y(n_602)
);

BUFx2_ASAP7_75t_SL g603 ( 
.A(n_541),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_556),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_558),
.Y(n_605)
);

BUFx2_ASAP7_75t_R g606 ( 
.A(n_581),
.Y(n_606)
);

BUFx12f_ASAP7_75t_L g607 ( 
.A(n_550),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_584),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_546),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_531),
.B(n_492),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_554),
.A2(n_521),
.B(n_519),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_570),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_535),
.A2(n_516),
.B(n_509),
.Y(n_613)
);

OAI21x1_ASAP7_75t_L g614 ( 
.A1(n_566),
.A2(n_504),
.B(n_522),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_556),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_587),
.Y(n_616)
);

AO21x1_ASAP7_75t_L g617 ( 
.A1(n_585),
.A2(n_473),
.B(n_520),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_587),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_588),
.B(n_512),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_568),
.B(n_497),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_547),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_547),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_L g623 ( 
.A1(n_533),
.A2(n_468),
.B(n_125),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_548),
.Y(n_624)
);

OAI21x1_ASAP7_75t_L g625 ( 
.A1(n_571),
.A2(n_124),
.B(n_127),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_575),
.A2(n_129),
.B(n_131),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_582),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_543),
.B(n_553),
.Y(n_628)
);

AO21x2_ASAP7_75t_L g629 ( 
.A1(n_539),
.A2(n_132),
.B(n_133),
.Y(n_629)
);

CKINVDCx16_ASAP7_75t_R g630 ( 
.A(n_550),
.Y(n_630)
);

BUFx8_ASAP7_75t_SL g631 ( 
.A(n_577),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_557),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_559),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_548),
.B(n_134),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_574),
.A2(n_538),
.B(n_580),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_560),
.Y(n_636)
);

AO21x2_ASAP7_75t_L g637 ( 
.A1(n_545),
.A2(n_135),
.B(n_138),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_542),
.A2(n_139),
.B(n_141),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_636),
.A2(n_564),
.B1(n_569),
.B2(n_563),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_598),
.Y(n_640)
);

BUFx10_ASAP7_75t_L g641 ( 
.A(n_619),
.Y(n_641)
);

CKINVDCx11_ASAP7_75t_R g642 ( 
.A(n_592),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_622),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_623),
.A2(n_549),
.B1(n_578),
.B2(n_567),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_595),
.A2(n_540),
.B(n_583),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_622),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_598),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_610),
.B(n_586),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_597),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_605),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_592),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_605),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_618),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_618),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_636),
.B(n_484),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_604),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_601),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_608),
.Y(n_658)
);

BUFx2_ASAP7_75t_SL g659 ( 
.A(n_604),
.Y(n_659)
);

CKINVDCx12_ASAP7_75t_R g660 ( 
.A(n_628),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_616),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_620),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_610),
.B(n_573),
.Y(n_663)
);

INVx6_ASAP7_75t_L g664 ( 
.A(n_615),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_596),
.Y(n_665)
);

NAND2x1p5_ASAP7_75t_L g666 ( 
.A(n_622),
.B(n_544),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_627),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_620),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_617),
.A2(n_555),
.B1(n_551),
.B2(n_484),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_632),
.B(n_572),
.Y(n_670)
);

OA21x2_ASAP7_75t_L g671 ( 
.A1(n_595),
.A2(n_561),
.B(n_145),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_612),
.Y(n_672)
);

INVx6_ASAP7_75t_L g673 ( 
.A(n_615),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_630),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_617),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_627),
.Y(n_676)
);

NAND2x1p5_ASAP7_75t_L g677 ( 
.A(n_634),
.B(n_153),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_633),
.B(n_154),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_621),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_621),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_635),
.A2(n_155),
.B1(n_158),
.B2(n_159),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_640),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_SL g683 ( 
.A1(n_655),
.A2(n_607),
.B1(n_620),
.B2(n_619),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_652),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_665),
.Y(n_685)
);

CKINVDCx16_ASAP7_75t_R g686 ( 
.A(n_651),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_672),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_643),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_679),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_R g690 ( 
.A(n_660),
.B(n_609),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_647),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_672),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_650),
.Y(n_693)
);

CKINVDCx16_ASAP7_75t_R g694 ( 
.A(n_649),
.Y(n_694)
);

OAI21x1_ASAP7_75t_SL g695 ( 
.A1(n_681),
.A2(n_599),
.B(n_613),
.Y(n_695)
);

INVx11_ASAP7_75t_L g696 ( 
.A(n_659),
.Y(n_696)
);

AO21x2_ASAP7_75t_L g697 ( 
.A1(n_645),
.A2(n_591),
.B(n_611),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_R g698 ( 
.A(n_663),
.B(n_648),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_658),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_648),
.B(n_619),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_661),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_657),
.Y(n_702)
);

NAND3xp33_ASAP7_75t_L g703 ( 
.A(n_644),
.B(n_602),
.C(n_634),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_662),
.B(n_668),
.Y(n_704)
);

CKINVDCx16_ASAP7_75t_R g705 ( 
.A(n_641),
.Y(n_705)
);

OAI21xp33_ASAP7_75t_SL g706 ( 
.A1(n_644),
.A2(n_638),
.B(n_625),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_670),
.B(n_593),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_642),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_680),
.B(n_603),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_678),
.B(n_602),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_R g711 ( 
.A(n_671),
.B(n_602),
.Y(n_711)
);

NAND2x1p5_ASAP7_75t_L g712 ( 
.A(n_643),
.B(n_634),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_678),
.B(n_631),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_667),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_676),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_653),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_639),
.A2(n_607),
.B1(n_629),
.B2(n_637),
.Y(n_717)
);

INVxp67_ASAP7_75t_SL g718 ( 
.A(n_654),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_646),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_641),
.B(n_624),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_639),
.B(n_631),
.Y(n_721)
);

AO31x2_ASAP7_75t_L g722 ( 
.A1(n_681),
.A2(n_591),
.A3(n_629),
.B(n_594),
.Y(n_722)
);

BUFx2_ASAP7_75t_SL g723 ( 
.A(n_656),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_SL g724 ( 
.A1(n_677),
.A2(n_637),
.B1(n_638),
.B2(n_626),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_646),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_679),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_671),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_679),
.B(n_600),
.Y(n_728)
);

NOR3xp33_ASAP7_75t_SL g729 ( 
.A(n_674),
.B(n_606),
.C(n_590),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_699),
.Y(n_730)
);

AND2x4_ASAP7_75t_SL g731 ( 
.A(n_687),
.B(n_656),
.Y(n_731)
);

NOR2x1_ASAP7_75t_SL g732 ( 
.A(n_703),
.B(n_656),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_687),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_710),
.B(n_677),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_700),
.B(n_674),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_701),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_690),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_692),
.B(n_669),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_721),
.B(n_669),
.Y(n_739)
);

INVxp67_ASAP7_75t_SL g740 ( 
.A(n_718),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_707),
.B(n_675),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_691),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_691),
.B(n_693),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_685),
.B(n_702),
.Y(n_744)
);

OR2x6_ASAP7_75t_L g745 ( 
.A(n_695),
.B(n_666),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_693),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_704),
.B(n_675),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_718),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_713),
.B(n_716),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_714),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_715),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_682),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_682),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_684),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_684),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_719),
.B(n_626),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_720),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_727),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_709),
.B(n_624),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_729),
.B(n_673),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_727),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_688),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_697),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_697),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_688),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_722),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_725),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_698),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_743),
.B(n_730),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_733),
.B(n_717),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_743),
.B(n_717),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_736),
.B(n_722),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_737),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_740),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_733),
.B(n_722),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_748),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_768),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_768),
.B(n_722),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_742),
.B(n_724),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_738),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_740),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_742),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_758),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_749),
.B(n_705),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_750),
.B(n_694),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_746),
.B(n_726),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_766),
.B(n_724),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_756),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_746),
.B(n_706),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_751),
.B(n_729),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_731),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_758),
.B(n_761),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_761),
.B(n_625),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_741),
.B(n_725),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_757),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_744),
.B(n_728),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_769),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_780),
.B(n_739),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_795),
.B(n_757),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_777),
.B(n_766),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_778),
.B(n_763),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_769),
.B(n_757),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_791),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_790),
.B(n_757),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_778),
.B(n_763),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_776),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_794),
.B(n_735),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_783),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_782),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_772),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_779),
.B(n_788),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_794),
.B(n_731),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_809),
.Y(n_813)
);

OAI322xp33_ASAP7_75t_L g814 ( 
.A1(n_810),
.A2(n_796),
.A3(n_775),
.B1(n_770),
.B2(n_787),
.C1(n_781),
.C2(n_785),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_808),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_801),
.Y(n_816)
);

NAND2x2_ASAP7_75t_L g817 ( 
.A(n_798),
.B(n_784),
.Y(n_817)
);

NOR2xp67_ASAP7_75t_L g818 ( 
.A(n_808),
.B(n_788),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_804),
.B(n_683),
.C(n_760),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_806),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_803),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_807),
.B(n_779),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_816),
.B(n_811),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_815),
.Y(n_824)
);

OA22x2_ASAP7_75t_L g825 ( 
.A1(n_821),
.A2(n_773),
.B1(n_811),
.B2(n_810),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_822),
.B(n_797),
.Y(n_826)
);

OAI21xp33_ASAP7_75t_L g827 ( 
.A1(n_819),
.A2(n_804),
.B(n_772),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_826),
.B(n_820),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_827),
.A2(n_817),
.B1(n_698),
.B2(n_771),
.Y(n_829)
);

AOI21xp33_ASAP7_75t_L g830 ( 
.A1(n_825),
.A2(n_813),
.B(n_800),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_823),
.A2(n_787),
.B1(n_821),
.B2(n_818),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_824),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_824),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_829),
.B(n_802),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_832),
.B(n_786),
.C(n_759),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_828),
.B(n_708),
.Y(n_836)
);

O2A1O1Ixp5_ASAP7_75t_SL g837 ( 
.A1(n_833),
.A2(n_767),
.B(n_765),
.C(n_762),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_836),
.B(n_831),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_835),
.A2(n_830),
.B1(n_771),
.B2(n_788),
.Y(n_839)
);

AO22x2_ASAP7_75t_L g840 ( 
.A1(n_834),
.A2(n_791),
.B1(n_774),
.B2(n_799),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_839),
.A2(n_686),
.B1(n_805),
.B2(n_791),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_840),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_838),
.B(n_814),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_838),
.B(n_837),
.Y(n_844)
);

NOR3xp33_ASAP7_75t_L g845 ( 
.A(n_844),
.B(n_726),
.C(n_689),
.Y(n_845)
);

NOR2xp67_ASAP7_75t_L g846 ( 
.A(n_842),
.B(n_689),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_843),
.Y(n_847)
);

OAI21xp5_ASAP7_75t_SL g848 ( 
.A1(n_841),
.A2(n_747),
.B(n_734),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_842),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_843),
.A2(n_786),
.B1(n_812),
.B2(n_723),
.Y(n_850)
);

NOR2x1_ASAP7_75t_L g851 ( 
.A(n_842),
.B(n_696),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_847),
.B(n_690),
.Y(n_852)
);

BUFx4f_ASAP7_75t_SL g853 ( 
.A(n_849),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_L g854 ( 
.A(n_845),
.B(n_614),
.C(n_786),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_851),
.B(n_664),
.Y(n_855)
);

OAI222xp33_ASAP7_75t_L g856 ( 
.A1(n_850),
.A2(n_745),
.B1(n_775),
.B2(n_789),
.C1(n_712),
.C2(n_754),
.Y(n_856)
);

NOR4xp75_ASAP7_75t_SL g857 ( 
.A(n_846),
.B(n_673),
.C(n_664),
.D(n_732),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_848),
.B(n_789),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_853),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_852),
.A2(n_745),
.B(n_756),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_855),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_858),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_854),
.B(n_783),
.Y(n_863)
);

CKINVDCx14_ASAP7_75t_R g864 ( 
.A(n_857),
.Y(n_864)
);

CKINVDCx16_ASAP7_75t_R g865 ( 
.A(n_856),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_862),
.Y(n_866)
);

AO22x2_ASAP7_75t_L g867 ( 
.A1(n_859),
.A2(n_664),
.B1(n_673),
.B2(n_764),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_865),
.A2(n_745),
.B1(n_756),
.B2(n_711),
.Y(n_868)
);

AOI22x1_ASAP7_75t_L g869 ( 
.A1(n_861),
.A2(n_712),
.B1(n_666),
.B2(n_764),
.Y(n_869)
);

AOI22x1_ASAP7_75t_L g870 ( 
.A1(n_864),
.A2(n_755),
.B1(n_753),
.B2(n_752),
.Y(n_870)
);

XOR2xp5_ASAP7_75t_L g871 ( 
.A(n_860),
.B(n_160),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_863),
.B(n_161),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_866),
.B(n_792),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_872),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_L g875 ( 
.A1(n_868),
.A2(n_755),
.B1(n_753),
.B2(n_752),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_SL g876 ( 
.A1(n_870),
.A2(n_793),
.B1(n_792),
.B2(n_614),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_871),
.A2(n_867),
.B1(n_869),
.B2(n_711),
.Y(n_877)
);

AND3x1_ASAP7_75t_L g878 ( 
.A(n_874),
.B(n_793),
.C(n_163),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_SL g879 ( 
.A1(n_877),
.A2(n_162),
.B1(n_168),
.B2(n_170),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_SL g880 ( 
.A1(n_873),
.A2(n_200),
.B1(n_172),
.B2(n_173),
.Y(n_880)
);

OAI222xp33_ASAP7_75t_L g881 ( 
.A1(n_880),
.A2(n_876),
.B1(n_875),
.B2(n_179),
.C1(n_180),
.C2(n_183),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_878),
.Y(n_882)
);

XNOR2xp5_ASAP7_75t_L g883 ( 
.A(n_882),
.B(n_879),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_SL g884 ( 
.A1(n_883),
.A2(n_881),
.B1(n_176),
.B2(n_184),
.Y(n_884)
);

AOI221x1_ASAP7_75t_L g885 ( 
.A1(n_884),
.A2(n_171),
.B1(n_185),
.B2(n_186),
.C(n_187),
.Y(n_885)
);

AOI211xp5_ASAP7_75t_L g886 ( 
.A1(n_885),
.A2(n_189),
.B(n_191),
.C(n_192),
.Y(n_886)
);


endmodule