module fake_aes_12067_n_40 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
wire n_39;
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_5), .Y(n_12) );
INVx3_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_2), .Y(n_17) );
OA21x2_ASAP7_75t_L g18 ( .A1(n_9), .A2(n_4), .B(n_3), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_13), .B(n_0), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_16), .B(n_0), .Y(n_21) );
NOR2x1_ASAP7_75t_L g22 ( .A(n_13), .B(n_6), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_19), .B(n_15), .Y(n_23) );
AOI22xp33_ASAP7_75t_SL g24 ( .A1(n_21), .A2(n_12), .B1(n_17), .B2(n_14), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
INVx4_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_20), .B1(n_17), .B2(n_14), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_26), .B(n_23), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_27), .B(n_25), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
CKINVDCx5p33_ASAP7_75t_R g31 ( .A(n_29), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_30), .B(n_25), .Y(n_32) );
A2O1A1Ixp33_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_13), .B(n_15), .C(n_18), .Y(n_33) );
OAI21xp33_ASAP7_75t_SL g34 ( .A1(n_31), .A2(n_13), .B(n_15), .Y(n_34) );
NOR3xp33_ASAP7_75t_SL g35 ( .A(n_34), .B(n_18), .C(n_2), .Y(n_35) );
OR2x2_ASAP7_75t_L g36 ( .A(n_32), .B(n_1), .Y(n_36) );
NAND2xp5_ASAP7_75t_L g37 ( .A(n_33), .B(n_18), .Y(n_37) );
AOI22xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_18), .B1(n_1), .B2(n_8), .Y(n_38) );
HB1xp67_ASAP7_75t_L g39 ( .A(n_36), .Y(n_39) );
AOI222xp33_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_7), .B1(n_11), .B2(n_18), .C1(n_37), .C2(n_38), .Y(n_40) );
endmodule