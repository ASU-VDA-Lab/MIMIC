module fake_jpeg_9516_n_208 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_41),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_28),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_31),
.B1(n_22),
.B2(n_27),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_53),
.B1(n_2),
.B2(n_3),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_31),
.B1(n_22),
.B2(n_34),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_52),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_31),
.B1(n_34),
.B2(n_19),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_27),
.B1(n_33),
.B2(n_25),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_1),
.B(n_2),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_67),
.B(n_1),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_32),
.B1(n_33),
.B2(n_19),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_58),
.B(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_62),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_18),
.C(n_20),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_24),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_68),
.Y(n_95)
);

FAx1_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_21),
.CI(n_27),
.CON(n_67),
.SN(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_24),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_40),
.B1(n_28),
.B2(n_43),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_82),
.B1(n_86),
.B2(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_77),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_75),
.B1(n_83),
.B2(n_66),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_26),
.B1(n_23),
.B2(n_18),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_76),
.A2(n_97),
.B(n_12),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_2),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_81),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_58),
.B1(n_64),
.B2(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_14),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_56),
.B1(n_47),
.B2(n_63),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_87),
.B1(n_94),
.B2(n_66),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_9),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_14),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_60),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_97),
.A2(n_49),
.B1(n_62),
.B2(n_59),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_108),
.B1(n_113),
.B2(n_114),
.Y(n_132)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_118),
.Y(n_136)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_73),
.B(n_72),
.C(n_71),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_112),
.B(n_72),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_71),
.A2(n_59),
.B1(n_69),
.B2(n_47),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_59),
.B1(n_69),
.B2(n_47),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_79),
.A2(n_69),
.B1(n_65),
.B2(n_13),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_115),
.A2(n_116),
.B1(n_89),
.B2(n_76),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_71),
.B(n_11),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_117),
.A2(n_77),
.B(n_91),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_121),
.A2(n_137),
.B1(n_140),
.B2(n_115),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_133),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_103),
.A3(n_12),
.B1(n_111),
.B2(n_70),
.Y(n_158)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_96),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_107),
.C(n_108),
.Y(n_148)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_130),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_89),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

BUFx4f_ASAP7_75t_SL g135 ( 
.A(n_109),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_99),
.B(n_81),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_117),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_80),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_101),
.C(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_114),
.B1(n_112),
.B2(n_110),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_147),
.B1(n_121),
.B2(n_132),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_145),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_101),
.C(n_112),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_148),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_78),
.C(n_94),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_153),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_98),
.C(n_106),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_132),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_156),
.Y(n_171)
);

OA21x2_ASAP7_75t_SL g156 ( 
.A1(n_139),
.A2(n_103),
.B(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_158),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_134),
.B1(n_136),
.B2(n_138),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_159),
.A2(n_142),
.B1(n_136),
.B2(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_131),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_120),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_167),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_170),
.B1(n_70),
.B2(n_84),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_127),
.A3(n_144),
.B1(n_122),
.B2(n_135),
.C1(n_143),
.C2(n_130),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_125),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_135),
.C(n_84),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_160),
.A2(n_145),
.B1(n_149),
.B2(n_152),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_149),
.B1(n_153),
.B2(n_146),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_146),
.B1(n_124),
.B2(n_128),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_166),
.B(n_161),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_163),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_172),
.A2(n_109),
.B1(n_135),
.B2(n_100),
.Y(n_182)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_165),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_185),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_162),
.B(n_164),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_190),
.B(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_178),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_166),
.B(n_163),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_174),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_180),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_197),
.C(n_190),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_194),
.B(n_195),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_188),
.A2(n_176),
.B1(n_182),
.B2(n_183),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_173),
.B1(n_181),
.B2(n_187),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_201),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_192),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_195),
.B(n_187),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.C(n_199),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_185),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_206),
.B(n_203),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_179),
.Y(n_208)
);


endmodule