module fake_jpeg_30847_n_530 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_530);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_530;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_57),
.B(n_64),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_61),
.Y(n_114)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_15),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_65),
.Y(n_171)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_80),
.Y(n_156)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_36),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_82),
.A2(n_53),
.B1(n_51),
.B2(n_17),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

CKINVDCx9p33_ASAP7_75t_R g84 ( 
.A(n_43),
.Y(n_84)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_26),
.B(n_37),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_90),
.B(n_101),
.Y(n_151)
);

BUFx12f_ASAP7_75t_SL g91 ( 
.A(n_21),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g137 ( 
.A(n_91),
.Y(n_137)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_19),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_107),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_105),
.Y(n_164)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_106),
.B(n_108),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_44),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_34),
.C(n_40),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_115),
.B(n_16),
.C(n_20),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_64),
.B(n_54),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_121),
.B(n_125),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_54),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_55),
.B(n_37),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_127),
.B(n_128),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_35),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_61),
.A2(n_46),
.B(n_49),
.C(n_107),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g208 ( 
.A1(n_134),
.A2(n_138),
.B1(n_33),
.B2(n_44),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_29),
.B1(n_52),
.B2(n_45),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_136),
.A2(n_141),
.B1(n_153),
.B2(n_162),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_63),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_107),
.A2(n_29),
.B1(n_52),
.B2(n_45),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_145),
.B1(n_163),
.B2(n_169),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_60),
.A2(n_52),
.B1(n_45),
.B2(n_53),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_52),
.B1(n_34),
.B2(n_40),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_101),
.A2(n_48),
.B1(n_24),
.B2(n_39),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_68),
.A2(n_72),
.B1(n_97),
.B2(n_96),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_89),
.A2(n_48),
.B1(n_39),
.B2(n_38),
.Y(n_163)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_59),
.B1(n_56),
.B2(n_105),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_176),
.A2(n_198),
.B1(n_202),
.B2(n_209),
.Y(n_240)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_117),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_179),
.B(n_191),
.Y(n_234)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_86),
.B1(n_76),
.B2(n_75),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_181),
.A2(n_182),
.B1(n_208),
.B2(n_212),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_131),
.A2(n_94),
.B1(n_16),
.B2(n_17),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_184),
.Y(n_263)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_188),
.B(n_206),
.Y(n_262)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

BUFx2_ASAP7_75t_SL g190 ( 
.A(n_114),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_190),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_155),
.B(n_38),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_192),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_134),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_193),
.B(n_197),
.Y(n_258)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_199),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_20),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_200),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_163),
.A2(n_56),
.B1(n_59),
.B2(n_22),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_196),
.A2(n_154),
.B1(n_149),
.B2(n_166),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_113),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_156),
.A2(n_22),
.B1(n_27),
.B2(n_24),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_132),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_27),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_156),
.A2(n_43),
.B1(n_33),
.B2(n_9),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_205),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_144),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_157),
.A2(n_33),
.B1(n_14),
.B2(n_12),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_119),
.B(n_12),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_219),
.Y(n_238)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_211),
.B(n_216),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_145),
.A2(n_33),
.B1(n_11),
.B2(n_10),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_165),
.B(n_9),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_213),
.B(n_0),
.Y(n_251)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_135),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_215),
.A2(n_123),
.B1(n_157),
.B2(n_158),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_139),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_111),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_140),
.A2(n_33),
.B1(n_44),
.B2(n_3),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_113),
.B1(n_129),
.B2(n_167),
.Y(n_235)
);

BUFx12_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g260 ( 
.A(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_111),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_130),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_223),
.A2(n_172),
.B1(n_133),
.B2(n_148),
.Y(n_261)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_130),
.Y(n_224)
);

BUFx12_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_118),
.B(n_0),
.Y(n_225)
);

AND2x4_ASAP7_75t_SL g226 ( 
.A(n_171),
.B(n_44),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_133),
.C(n_143),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_235),
.A2(n_239),
.B1(n_244),
.B2(n_256),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_183),
.A2(n_118),
.B1(n_167),
.B2(n_150),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_249),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_175),
.A2(n_136),
.B(n_162),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_242),
.A2(n_199),
.B(n_148),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_204),
.A2(n_150),
.B1(n_158),
.B2(n_143),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_218),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_204),
.A2(n_166),
.B1(n_160),
.B2(n_154),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_200),
.B(n_160),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_180),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_261),
.A2(n_194),
.B1(n_197),
.B2(n_223),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_267),
.B(n_277),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_254),
.Y(n_268)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_268),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_187),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_282),
.C(n_292),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_270),
.Y(n_300)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_254),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_275),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_228),
.Y(n_274)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_274),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_231),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_227),
.B(n_207),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_278),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_234),
.B(n_238),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_247),
.B(n_207),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_242),
.A2(n_225),
.B1(n_196),
.B2(n_208),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_279),
.A2(n_284),
.B1(n_295),
.B2(n_287),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_208),
.B1(n_174),
.B2(n_226),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_280),
.A2(n_288),
.B1(n_291),
.B2(n_293),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_228),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_281),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_188),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_233),
.Y(n_283)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_283),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_245),
.A2(n_208),
.B1(n_195),
.B2(n_135),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_285),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_241),
.B(n_226),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_287),
.A2(n_253),
.B(n_264),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_244),
.A2(n_192),
.B1(n_211),
.B2(n_216),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_294),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_243),
.A2(n_205),
.B1(n_206),
.B2(n_201),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_239),
.B1(n_235),
.B2(n_249),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_243),
.A2(n_184),
.B1(n_178),
.B2(n_186),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_247),
.B(n_210),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_258),
.A2(n_149),
.B1(n_172),
.B2(n_123),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_222),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_296),
.A2(n_240),
.B(n_266),
.Y(n_303)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_260),
.Y(n_297)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_258),
.A2(n_173),
.B1(n_215),
.B2(n_219),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_298),
.A2(n_263),
.B1(n_248),
.B2(n_253),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_299),
.Y(n_345)
);

NOR2x1_ASAP7_75t_R g302 ( 
.A(n_274),
.B(n_281),
.Y(n_302)
);

OA21x2_ASAP7_75t_L g354 ( 
.A1(n_302),
.A2(n_314),
.B(n_327),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_303),
.A2(n_317),
.B(n_320),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_279),
.A2(n_245),
.B1(n_231),
.B2(n_234),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_304),
.A2(n_312),
.B1(n_326),
.B2(n_328),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_238),
.B1(n_228),
.B2(n_265),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_305),
.A2(n_293),
.B1(n_298),
.B2(n_283),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_284),
.A2(n_251),
.B1(n_250),
.B2(n_252),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_267),
.B(n_232),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_315),
.B(n_321),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_274),
.A2(n_230),
.B(n_229),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_286),
.A2(n_230),
.B(n_229),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_277),
.B(n_232),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_252),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_324),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_237),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_289),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_263),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_327),
.A2(n_255),
.B(n_236),
.Y(n_353)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_324),
.Y(n_329)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_329),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_305),
.A2(n_286),
.B1(n_278),
.B2(n_276),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_330),
.A2(n_331),
.B1(n_334),
.B2(n_344),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_309),
.A2(n_286),
.B1(n_287),
.B2(n_272),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_309),
.A2(n_286),
.B1(n_287),
.B2(n_272),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_306),
.Y(n_335)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_335),
.Y(n_385)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_306),
.Y(n_336)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_336),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_308),
.Y(n_337)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_337),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_304),
.A2(n_328),
.B1(n_312),
.B2(n_280),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_339),
.A2(n_350),
.B1(n_314),
.B2(n_316),
.Y(n_368)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_301),
.Y(n_340)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_340),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_282),
.C(n_269),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_325),
.C(n_203),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_323),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_271),
.Y(n_343)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_343),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_285),
.Y(n_346)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_346),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_328),
.A2(n_288),
.B1(n_268),
.B2(n_273),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_355),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_315),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_348),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

BUFx8_ASAP7_75t_L g365 ( 
.A(n_349),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_299),
.A2(n_291),
.B1(n_273),
.B2(n_263),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_311),
.B(n_255),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_351),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_353),
.A2(n_317),
.B(n_320),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_354),
.A2(n_319),
.B(n_310),
.Y(n_375)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_301),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_236),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_357),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_318),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_318),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_325),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_313),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_360),
.B(n_363),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_313),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_364),
.B(n_382),
.C(n_386),
.Y(n_404)
);

A2O1A1Ixp33_ASAP7_75t_SL g367 ( 
.A1(n_354),
.A2(n_302),
.B(n_320),
.C(n_317),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_367),
.A2(n_372),
.B(n_380),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_368),
.B(n_347),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_348),
.B(n_307),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_370),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_340),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_338),
.B(n_307),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_351),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_345),
.A2(n_303),
.B1(n_316),
.B2(n_302),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_375),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_352),
.A2(n_319),
.B(n_310),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_377),
.A2(n_388),
.B(n_344),
.Y(n_418)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_379),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_SL g380 ( 
.A(n_352),
.B(n_323),
.C(n_326),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_337),
.B(n_300),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_384),
.A2(n_339),
.B1(n_332),
.B2(n_353),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_330),
.B(n_237),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_354),
.A2(n_300),
.B(n_297),
.Y(n_388)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_373),
.Y(n_391)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_391),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_376),
.A2(n_350),
.B1(n_345),
.B2(n_338),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_393),
.A2(n_405),
.B1(n_408),
.B2(n_410),
.Y(n_424)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_373),
.Y(n_394)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_394),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_396),
.B(n_397),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_389),
.B(n_346),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_379),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_400),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_384),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_372),
.A2(n_354),
.B(n_336),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_407),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_378),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_402),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_380),
.A2(n_335),
.B(n_329),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_367),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_366),
.B(n_343),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_406),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_359),
.A2(n_332),
.B1(n_331),
.B2(n_334),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_366),
.B(n_356),
.Y(n_409)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_409),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_365),
.Y(n_410)
);

OAI32xp33_ASAP7_75t_L g411 ( 
.A1(n_361),
.A2(n_333),
.A3(n_344),
.B1(n_357),
.B2(n_358),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_411),
.B(n_416),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_364),
.B(n_360),
.C(n_382),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_413),
.B(n_363),
.C(n_386),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_365),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_414),
.B(n_365),
.Y(n_438)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_378),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_415),
.A2(n_355),
.B1(n_387),
.B2(n_383),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_383),
.B(n_333),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_361),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_417),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_418),
.A2(n_368),
.B(n_367),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_412),
.B(n_404),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_419),
.B(n_442),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_423),
.C(n_426),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_377),
.C(n_342),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_404),
.C(n_403),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_395),
.B(n_342),
.C(n_388),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_427),
.B(n_434),
.C(n_398),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_395),
.B(n_374),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_432),
.B(n_411),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_398),
.A2(n_385),
.B1(n_381),
.B2(n_362),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_433),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_390),
.B(n_375),
.C(n_362),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_435),
.A2(n_407),
.B(n_433),
.Y(n_456)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_438),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_439),
.B(n_441),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_392),
.A2(n_387),
.B1(n_349),
.B2(n_300),
.Y(n_441)
);

FAx1_ASAP7_75t_SL g444 ( 
.A(n_442),
.B(n_416),
.CI(n_409),
.CON(n_444),
.SN(n_444)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_454),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_451),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_424),
.A2(n_418),
.B1(n_399),
.B2(n_398),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_446),
.A2(n_455),
.B1(n_457),
.B2(n_248),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_420),
.B(n_396),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_448),
.B(n_453),
.Y(n_473)
);

XNOR2x1_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_397),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_426),
.A2(n_392),
.B(n_390),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_425),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_431),
.A2(n_440),
.B1(n_437),
.B2(n_430),
.Y(n_455)
);

AOI221xp5_ASAP7_75t_L g464 ( 
.A1(n_456),
.A2(n_435),
.B1(n_428),
.B2(n_432),
.C(n_436),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_431),
.A2(n_391),
.B1(n_394),
.B2(n_402),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_408),
.C(n_405),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_458),
.B(n_459),
.C(n_460),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_422),
.B(n_401),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_423),
.B(n_406),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_189),
.C(n_185),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_449),
.B(n_410),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_467),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_472),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_459),
.A2(n_428),
.B1(n_421),
.B2(n_417),
.Y(n_465)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_465),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_434),
.C(n_429),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_470),
.C(n_260),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_461),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_SL g468 ( 
.A1(n_456),
.A2(n_414),
.B1(n_349),
.B2(n_415),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_468),
.A2(n_476),
.B1(n_477),
.B2(n_224),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_445),
.C(n_458),
.Y(n_470)
);

NOR2x1_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_421),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_474),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_450),
.A2(n_429),
.B1(n_367),
.B2(n_217),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_450),
.A2(n_270),
.B1(n_248),
.B2(n_177),
.Y(n_474)
);

OAI321xp33_ASAP7_75t_L g476 ( 
.A1(n_447),
.A2(n_270),
.A3(n_237),
.B1(n_230),
.B2(n_197),
.C(n_260),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_478),
.B(n_173),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_454),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_485),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_471),
.A2(n_451),
.B1(n_444),
.B2(n_460),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_482),
.Y(n_507)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_483),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_472),
.A2(n_444),
.B1(n_452),
.B2(n_214),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_462),
.B(n_452),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_490),
.C(n_494),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_230),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_489),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_260),
.Y(n_489)
);

CKINVDCx14_ASAP7_75t_R g491 ( 
.A(n_473),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_491),
.B(n_492),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_469),
.A2(n_257),
.B1(n_1),
.B2(n_3),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_493),
.B(n_0),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_257),
.C(n_221),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_482),
.A2(n_465),
.B(n_462),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_498),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_480),
.A2(n_475),
.B1(n_221),
.B2(n_257),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_499),
.B(n_4),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_257),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_502),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_485),
.A2(n_486),
.B(n_490),
.Y(n_502)
);

OA21x2_ASAP7_75t_SL g504 ( 
.A1(n_487),
.A2(n_494),
.B(n_484),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_504),
.B(n_1),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_484),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_3),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_508),
.A2(n_497),
.B(n_503),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_44),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_510),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_501),
.B(n_4),
.C(n_5),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_513),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_505),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_514),
.B(n_496),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_518),
.B(n_519),
.Y(n_522)
);

AO21x1_ASAP7_75t_L g519 ( 
.A1(n_515),
.A2(n_502),
.B(n_495),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_520),
.B(n_511),
.C(n_507),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_519),
.A2(n_508),
.B(n_507),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_521),
.A2(n_523),
.B(n_517),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_524),
.B(n_525),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_522),
.A2(n_516),
.B(n_498),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_SL g527 ( 
.A1(n_526),
.A2(n_514),
.B(n_7),
.C(n_8),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_527),
.A2(n_5),
.B(n_7),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_7),
.B1(n_8),
.B2(n_376),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_8),
.Y(n_530)
);


endmodule