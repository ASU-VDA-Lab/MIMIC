module fake_ariane_1643_n_2072 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2072);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2072;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_4),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_123),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_89),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_126),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_152),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_18),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_115),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_32),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_201),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_83),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_86),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_19),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_67),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_8),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_91),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_2),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_114),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_147),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_80),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_49),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_129),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_95),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_111),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_104),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_151),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_15),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_64),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_130),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_77),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_96),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_1),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_8),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_63),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_34),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_70),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_142),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_205),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_76),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_165),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_102),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_41),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_145),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_105),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_86),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_71),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_178),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_133),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_184),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_141),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_50),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_103),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_78),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_192),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_28),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_180),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_132),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_190),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_55),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_80),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_79),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_68),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_154),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_16),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_19),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_98),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_166),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_139),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_88),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_128),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_15),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_10),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_200),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_65),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_173),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_32),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_127),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_13),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_117),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_97),
.Y(n_294)
);

BUFx5_ASAP7_75t_L g295 ( 
.A(n_12),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_46),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_76),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_43),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_69),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_198),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_26),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_195),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_16),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_148),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_109),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_183),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_43),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_62),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_72),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_124),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_75),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_167),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_181),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_85),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_77),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_28),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_169),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_99),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_47),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_206),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_189),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_5),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_3),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_9),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_134),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_39),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_45),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_85),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_6),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_137),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_107),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_73),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_75),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_49),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_31),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_140),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_1),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_158),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_74),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_11),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_203),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_65),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_61),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_155),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_161),
.Y(n_345)
);

BUFx10_ASAP7_75t_L g346 ( 
.A(n_177),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_48),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_172),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_125),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_191),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_92),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_83),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_46),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_144),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_143),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_135),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_70),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_81),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_153),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_37),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_82),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_35),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_14),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_10),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_67),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_101),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_58),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_41),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_185),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_199),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_42),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_30),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_156),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_51),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_87),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_29),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_24),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_136),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_149),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_110),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_84),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_34),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_79),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_6),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_17),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_78),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_18),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_100),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_64),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_82),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_193),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_29),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_31),
.Y(n_393)
);

CKINVDCx14_ASAP7_75t_R g394 ( 
.A(n_69),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_44),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_73),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_168),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_66),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_131),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_150),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_56),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_0),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_174),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_93),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_4),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_394),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_326),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_365),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_295),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_235),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_238),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_326),
.B(n_2),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_295),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_295),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_242),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_252),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_261),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_222),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_295),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_295),
.B(n_3),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_295),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_263),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_270),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_295),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_295),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_295),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_326),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_208),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_208),
.B(n_5),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_337),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_310),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_212),
.Y(n_432)
);

BUFx10_ASAP7_75t_L g433 ( 
.A(n_219),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_212),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_221),
.B(n_7),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_221),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_229),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_320),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_229),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_336),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_230),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_337),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_354),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_222),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_230),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_356),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_233),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_285),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_256),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_256),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_233),
.B(n_9),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_334),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_298),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g454 ( 
.A(n_217),
.B(n_11),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_236),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_236),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_223),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_334),
.Y(n_458)
);

BUFx6f_ASAP7_75t_SL g459 ( 
.A(n_247),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_224),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_232),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_234),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_244),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_244),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_403),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_209),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_301),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_240),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_352),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_251),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_251),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_209),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_311),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_255),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_352),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_243),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_322),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_352),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_352),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_403),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g481 ( 
.A(n_217),
.B(n_13),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_254),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_255),
.Y(n_483)
);

BUFx6f_ASAP7_75t_SL g484 ( 
.A(n_247),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_245),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_258),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_257),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_257),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_248),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_L g490 ( 
.A(n_220),
.B(n_14),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_271),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_317),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_253),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_352),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_402),
.Y(n_495)
);

INVxp33_ASAP7_75t_SL g496 ( 
.A(n_260),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_271),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_283),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_283),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_289),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_247),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_269),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_225),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_289),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_402),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_273),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_293),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_274),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_247),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_402),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_293),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_346),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_346),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_302),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_409),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_409),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_469),
.B(n_302),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_428),
.B(n_402),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_478),
.B(n_305),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_421),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_421),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_413),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_413),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_449),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_428),
.B(n_220),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_432),
.B(n_275),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_414),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_414),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_430),
.A2(n_241),
.B1(n_249),
.B2(n_215),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_419),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_424),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_411),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_433),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_461),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_425),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_425),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_432),
.B(n_402),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_426),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_434),
.B(n_275),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_475),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_479),
.B(n_305),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_426),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_433),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_434),
.B(n_276),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_436),
.B(n_276),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_475),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_475),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_433),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_494),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_495),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_436),
.B(n_225),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_476),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_505),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_412),
.B(n_219),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_510),
.B(n_306),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_437),
.B(n_439),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_427),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_427),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_448),
.B(n_286),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_433),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_420),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_437),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_439),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_441),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_441),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_445),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_445),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_407),
.B(n_306),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_447),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_502),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_447),
.B(n_312),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_418),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_455),
.B(n_312),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_455),
.B(n_226),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_456),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_456),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_463),
.B(n_321),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_463),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_464),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_464),
.B(n_470),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_450),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_470),
.Y(n_585)
);

AND2x6_ASAP7_75t_L g586 ( 
.A(n_471),
.B(n_219),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_471),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_474),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_474),
.B(n_321),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_483),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_483),
.B(n_330),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_487),
.B(n_226),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_487),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_488),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_488),
.B(n_346),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_491),
.Y(n_596)
);

INVx6_ASAP7_75t_L g597 ( 
.A(n_418),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_491),
.B(n_497),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_480),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_497),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_453),
.B(n_467),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_442),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_602),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_595),
.A2(n_465),
.B1(n_482),
.B2(n_408),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_597),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_559),
.B(n_465),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_572),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_564),
.B(n_498),
.Y(n_608)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_557),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_570),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_570),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_552),
.B(n_482),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_595),
.B(n_418),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_581),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_601),
.Y(n_615)
);

AND2x6_ASAP7_75t_L g616 ( 
.A(n_595),
.B(n_330),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_597),
.Y(n_617)
);

AND2x2_ASAP7_75t_SL g618 ( 
.A(n_554),
.B(n_451),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_551),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_523),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_572),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_523),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_575),
.B(n_444),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_582),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_535),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_582),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_537),
.A2(n_496),
.B1(n_429),
.B2(n_435),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_525),
.B(n_454),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_523),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_585),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_575),
.B(n_444),
.Y(n_631)
);

AOI21x1_ASAP7_75t_L g632 ( 
.A1(n_515),
.A2(n_499),
.B(n_498),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_552),
.B(n_457),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_572),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_523),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_572),
.Y(n_636)
);

NAND3xp33_ASAP7_75t_L g637 ( 
.A(n_555),
.B(n_462),
.C(n_460),
.Y(n_637)
);

AO22x2_ASAP7_75t_L g638 ( 
.A1(n_530),
.A2(n_500),
.B1(n_504),
.B2(n_499),
.Y(n_638)
);

AND2x6_ASAP7_75t_L g639 ( 
.A(n_564),
.B(n_331),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_529),
.Y(n_640)
);

NAND2x1p5_ASAP7_75t_L g641 ( 
.A(n_564),
.B(n_500),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_553),
.B(n_468),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_529),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_575),
.B(n_444),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_553),
.B(n_485),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_551),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_572),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_602),
.B(n_442),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_585),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_555),
.B(n_489),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_573),
.B(n_493),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_551),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_587),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_557),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_559),
.B(n_598),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_572),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_551),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_573),
.A2(n_508),
.B1(n_506),
.B2(n_484),
.Y(n_658)
);

NOR2x1p5_ASAP7_75t_L g659 ( 
.A(n_535),
.B(n_415),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_529),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_525),
.B(n_584),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_529),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_557),
.A2(n_459),
.B1(n_484),
.B2(n_481),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_587),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_531),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_556),
.B(n_459),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_590),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_525),
.B(n_584),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_597),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_597),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_557),
.A2(n_459),
.B1(n_484),
.B2(n_481),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_559),
.B(n_486),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_531),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_590),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_517),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_531),
.Y(n_676)
);

AOI21x1_ASAP7_75t_L g677 ( 
.A1(n_515),
.A2(n_507),
.B(n_504),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_584),
.B(n_416),
.Y(n_678)
);

XNOR2xp5_ASAP7_75t_L g679 ( 
.A(n_562),
.B(n_473),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_517),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_598),
.B(n_492),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_531),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_530),
.B(n_417),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_556),
.B(n_486),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_572),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_517),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_557),
.A2(n_459),
.B1(n_484),
.B2(n_454),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_598),
.B(n_486),
.Y(n_688)
);

AND2x6_ASAP7_75t_L g689 ( 
.A(n_564),
.B(n_331),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_572),
.Y(n_690)
);

INVx4_ASAP7_75t_L g691 ( 
.A(n_551),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_597),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_533),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_533),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_578),
.Y(n_695)
);

BUFx4f_ASAP7_75t_L g696 ( 
.A(n_564),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_533),
.Y(n_697)
);

INVx5_ASAP7_75t_L g698 ( 
.A(n_557),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_563),
.B(n_507),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_533),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_L g701 ( 
.A(n_557),
.B(n_341),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_571),
.B(n_422),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_594),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_526),
.B(n_511),
.Y(n_704)
);

OAI22xp33_ASAP7_75t_L g705 ( 
.A1(n_571),
.A2(n_324),
.B1(n_340),
.B2(n_314),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_534),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_578),
.Y(n_707)
);

OAI21xp33_ASAP7_75t_L g708 ( 
.A1(n_583),
.A2(n_596),
.B(n_576),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_578),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_597),
.B(n_406),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_578),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_601),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_551),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_596),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_563),
.B(n_569),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_SL g716 ( 
.A(n_599),
.B(n_501),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_578),
.Y(n_717)
);

AND2x6_ASAP7_75t_L g718 ( 
.A(n_564),
.B(n_341),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_534),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_578),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_557),
.A2(n_512),
.B1(n_513),
.B2(n_509),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_560),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_578),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_563),
.B(n_511),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_517),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_563),
.B(n_514),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_557),
.B(n_349),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_534),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_601),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_599),
.B(n_423),
.Y(n_730)
);

NOR2x1p5_ASAP7_75t_L g731 ( 
.A(n_583),
.B(n_438),
.Y(n_731)
);

BUFx10_ASAP7_75t_L g732 ( 
.A(n_554),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_557),
.A2(n_490),
.B1(n_514),
.B2(n_228),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_R g734 ( 
.A(n_599),
.B(n_440),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_551),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_569),
.B(n_443),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_578),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_569),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_562),
.B(n_446),
.Y(n_739)
);

NAND2x1p5_ASAP7_75t_L g740 ( 
.A(n_564),
.B(n_258),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_534),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_563),
.B(n_452),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_569),
.B(n_466),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_569),
.B(n_588),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_588),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_518),
.B(n_458),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_588),
.A2(n_259),
.B1(n_292),
.B2(n_288),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_R g748 ( 
.A(n_588),
.B(n_410),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_516),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_588),
.B(n_250),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_SL g751 ( 
.A(n_557),
.B(n_431),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_593),
.B(n_250),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_620),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_732),
.B(n_546),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_742),
.B(n_593),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_603),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_738),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_738),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_L g759 ( 
.A(n_616),
.B(n_564),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_732),
.B(n_658),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_746),
.B(n_593),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_745),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_732),
.B(n_546),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_633),
.B(n_546),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_616),
.B(n_593),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_616),
.B(n_593),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_642),
.B(n_546),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_616),
.B(n_532),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_616),
.B(n_518),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_645),
.B(n_546),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_638),
.A2(n_554),
.B1(n_592),
.B2(n_577),
.Y(n_771)
);

O2A1O1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_688),
.A2(n_524),
.B(n_528),
.C(n_516),
.Y(n_772)
);

NAND3xp33_ASAP7_75t_L g773 ( 
.A(n_627),
.B(n_544),
.C(n_520),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_745),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_616),
.B(n_520),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_613),
.B(n_544),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_620),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_734),
.Y(n_778)
);

NOR3xp33_ASAP7_75t_L g779 ( 
.A(n_661),
.B(n_668),
.C(n_651),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_702),
.B(n_477),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_613),
.B(n_558),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_622),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_650),
.B(n_736),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_655),
.B(n_554),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_613),
.B(n_536),
.Y(n_785)
);

NOR3xp33_ASAP7_75t_L g786 ( 
.A(n_625),
.B(n_376),
.C(n_362),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_724),
.B(n_558),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_648),
.B(n_562),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_604),
.B(n_536),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_749),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_704),
.B(n_554),
.Y(n_791)
);

NOR2x1_ASAP7_75t_L g792 ( 
.A(n_637),
.B(n_574),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_612),
.B(n_561),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_629),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_704),
.B(n_554),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_655),
.B(n_536),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_672),
.B(n_577),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_655),
.B(n_577),
.Y(n_798)
);

NOR2xp67_ASAP7_75t_L g799 ( 
.A(n_625),
.B(n_576),
.Y(n_799)
);

OAI22x1_ASAP7_75t_SL g800 ( 
.A1(n_615),
.A2(n_297),
.B1(n_299),
.B2(n_296),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_606),
.B(n_577),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_606),
.B(n_577),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_629),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_672),
.B(n_577),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_672),
.B(n_592),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_743),
.B(n_592),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_708),
.B(n_592),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_681),
.B(n_561),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_638),
.A2(n_592),
.B1(n_542),
.B2(n_540),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_635),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_618),
.B(n_638),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_666),
.B(n_618),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_748),
.B(n_551),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_648),
.B(n_524),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_635),
.Y(n_815)
);

INVxp33_ASAP7_75t_L g816 ( 
.A(n_678),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_610),
.B(n_528),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_751),
.B(n_580),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_749),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_696),
.B(n_580),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_744),
.A2(n_545),
.B(n_541),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_696),
.A2(n_591),
.B1(n_589),
.B2(n_566),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_611),
.B(n_545),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_614),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_710),
.B(n_589),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_628),
.B(n_683),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_624),
.B(n_565),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_626),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_630),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_696),
.B(n_591),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_609),
.Y(n_831)
);

AND2x6_ASAP7_75t_L g832 ( 
.A(n_640),
.B(n_526),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_643),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_649),
.B(n_565),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_653),
.B(n_565),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_664),
.B(n_565),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_667),
.B(n_566),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_643),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_608),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_660),
.Y(n_840)
);

BUFx6f_ASAP7_75t_SL g841 ( 
.A(n_628),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_628),
.B(n_526),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_733),
.A2(n_542),
.B1(n_540),
.B2(n_519),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_674),
.B(n_566),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_660),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_730),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_SL g847 ( 
.A1(n_615),
.A2(n_729),
.B1(n_679),
.B2(n_712),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_662),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_703),
.B(n_567),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_730),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_662),
.Y(n_851)
);

AO221x1_ASAP7_75t_L g852 ( 
.A1(n_705),
.A2(n_503),
.B1(n_472),
.B2(n_747),
.C(n_246),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_714),
.B(n_567),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_665),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_721),
.B(n_567),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_722),
.B(n_684),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_665),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_608),
.Y(n_858)
);

NAND3xp33_ASAP7_75t_L g859 ( 
.A(n_701),
.B(n_541),
.C(n_539),
.Y(n_859)
);

NOR2xp67_ASAP7_75t_L g860 ( 
.A(n_683),
.B(n_568),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_699),
.B(n_568),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_609),
.B(n_568),
.Y(n_862)
);

INVx8_ASAP7_75t_L g863 ( 
.A(n_639),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_673),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_673),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_676),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_676),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_726),
.B(n_568),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_628),
.B(n_527),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_609),
.B(n_579),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_750),
.B(n_579),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_752),
.B(n_579),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_682),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_716),
.B(n_579),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_682),
.A2(n_600),
.B(n_539),
.C(n_541),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_641),
.B(n_693),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_693),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_641),
.B(n_600),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_701),
.A2(n_542),
.B1(n_547),
.B2(n_527),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_694),
.B(n_600),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_694),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_697),
.Y(n_882)
);

AOI221xp5_ASAP7_75t_L g883 ( 
.A1(n_727),
.A2(n_246),
.B1(n_265),
.B2(n_228),
.C(n_267),
.Y(n_883)
);

AND2x6_ASAP7_75t_L g884 ( 
.A(n_697),
.B(n_527),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_609),
.B(n_600),
.Y(n_885)
);

NAND2x1p5_ASAP7_75t_L g886 ( 
.A(n_609),
.B(n_522),
.Y(n_886)
);

BUFx8_ASAP7_75t_L g887 ( 
.A(n_739),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_727),
.A2(n_542),
.B1(n_548),
.B2(n_547),
.Y(n_888)
);

NAND2x1_ASAP7_75t_L g889 ( 
.A(n_621),
.B(n_522),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_700),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_731),
.B(n_547),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_700),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_706),
.B(n_548),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_706),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_739),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_719),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_712),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_719),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_728),
.B(n_548),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_605),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_740),
.B(n_542),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_715),
.B(n_539),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_654),
.B(n_519),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_728),
.B(n_741),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_741),
.B(n_522),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_632),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_632),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_677),
.Y(n_908)
);

NAND2xp33_ASAP7_75t_L g909 ( 
.A(n_675),
.B(n_532),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_623),
.B(n_631),
.Y(n_910)
);

AOI22x1_ASAP7_75t_L g911 ( 
.A1(n_621),
.A2(n_541),
.B1(n_539),
.B2(n_521),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_677),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_607),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_644),
.B(n_522),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_SL g915 ( 
.A(n_729),
.B(n_346),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_757),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_787),
.A2(n_646),
.B(n_619),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_850),
.B(n_816),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_793),
.B(n_639),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_910),
.A2(n_646),
.B(n_619),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_839),
.Y(n_921)
);

BUFx4f_ASAP7_75t_L g922 ( 
.A(n_842),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_842),
.B(n_659),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_757),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_816),
.B(n_679),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_811),
.A2(n_639),
.B1(n_718),
.B2(n_689),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_914),
.A2(n_646),
.B(n_619),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_758),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_812),
.B(n_675),
.Y(n_929)
);

NAND2x1_ASAP7_75t_L g930 ( 
.A(n_831),
.B(n_621),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_825),
.A2(n_636),
.B(n_656),
.C(n_634),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_814),
.B(n_639),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_755),
.A2(n_657),
.B(n_652),
.Y(n_933)
);

AOI21xp33_ASAP7_75t_L g934 ( 
.A1(n_874),
.A2(n_671),
.B(n_663),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_765),
.B(n_675),
.Y(n_935)
);

AOI21x1_ASAP7_75t_L g936 ( 
.A1(n_907),
.A2(n_647),
.B(n_607),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_876),
.A2(n_685),
.B(n_647),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_766),
.B(n_675),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_802),
.A2(n_265),
.B(n_278),
.C(n_267),
.Y(n_939)
);

NOR2x1_ASAP7_75t_L g940 ( 
.A(n_799),
.B(n_634),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_826),
.B(n_634),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_773),
.A2(n_490),
.B(n_540),
.C(n_519),
.Y(n_942)
);

BUFx2_ASAP7_75t_SL g943 ( 
.A(n_841),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_758),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_762),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_863),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_820),
.A2(n_657),
.B(n_652),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_902),
.A2(n_690),
.B(n_685),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_846),
.B(n_519),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_839),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_761),
.A2(n_652),
.B1(n_691),
.B2(n_657),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_801),
.B(n_776),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_830),
.A2(n_713),
.B(n_691),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_801),
.B(n_639),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_781),
.B(n_639),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_762),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_887),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_887),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_858),
.Y(n_959)
);

OAI321xp33_ASAP7_75t_L g960 ( 
.A1(n_883),
.A2(n_329),
.A3(n_278),
.B1(n_279),
.B2(n_385),
.C(n_290),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_860),
.B(n_784),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_858),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_811),
.A2(n_689),
.B1(n_718),
.B2(n_687),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_784),
.Y(n_964)
);

AOI21x1_ASAP7_75t_L g965 ( 
.A1(n_907),
.A2(n_711),
.B(n_690),
.Y(n_965)
);

AO21x1_ASAP7_75t_L g966 ( 
.A1(n_818),
.A2(n_740),
.B(n_711),
.Y(n_966)
);

OAI21xp33_ASAP7_75t_L g967 ( 
.A1(n_806),
.A2(n_307),
.B(n_303),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_753),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_804),
.B(n_689),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_783),
.A2(n_718),
.B1(n_689),
.B2(n_656),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_819),
.B(n_675),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_887),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_861),
.A2(n_713),
.B(n_691),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_868),
.A2(n_767),
.B(n_764),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_770),
.A2(n_735),
.B(n_713),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_759),
.A2(n_735),
.B(n_670),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_759),
.A2(n_735),
.B(n_670),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_842),
.B(n_636),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_856),
.A2(n_617),
.B(n_636),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_869),
.B(n_656),
.Y(n_980)
);

NOR2x1p5_ASAP7_75t_L g981 ( 
.A(n_788),
.B(n_279),
.Y(n_981)
);

BUFx4f_ASAP7_75t_L g982 ( 
.A(n_869),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_900),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_769),
.A2(n_695),
.B(n_709),
.C(n_707),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_774),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_909),
.A2(n_617),
.B(n_695),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_804),
.B(n_689),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_791),
.B(n_718),
.Y(n_988)
);

BUFx8_ASAP7_75t_SL g989 ( 
.A(n_841),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_795),
.B(n_718),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_819),
.B(n_680),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_909),
.A2(n_707),
.B(n_695),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_824),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_878),
.A2(n_709),
.B(n_707),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_863),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_775),
.B(n_680),
.Y(n_996)
);

OAI321xp33_ASAP7_75t_L g997 ( 
.A1(n_771),
.A2(n_383),
.A3(n_363),
.B1(n_385),
.B2(n_387),
.C(n_335),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_904),
.A2(n_717),
.B(n_709),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_821),
.A2(n_720),
.B(n_717),
.Y(n_999)
);

NAND2xp33_ASAP7_75t_L g1000 ( 
.A(n_832),
.B(n_884),
.Y(n_1000)
);

AND2x2_ASAP7_75t_SL g1001 ( 
.A(n_768),
.B(n_349),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_753),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_798),
.B(n_519),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_905),
.A2(n_880),
.B(n_763),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_828),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_829),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_754),
.A2(n_720),
.B(n_717),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_808),
.B(n_797),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_900),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_760),
.B(n_680),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_805),
.B(n_519),
.Y(n_1011)
);

BUFx4f_ASAP7_75t_L g1012 ( 
.A(n_869),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_871),
.A2(n_723),
.B(n_737),
.C(n_720),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_756),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_863),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_792),
.B(n_540),
.Y(n_1016)
);

CKINVDCx10_ASAP7_75t_R g1017 ( 
.A(n_841),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_817),
.A2(n_737),
.B1(n_723),
.B2(n_686),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_872),
.A2(n_737),
.B(n_723),
.C(n_698),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_913),
.B(n_680),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_913),
.A2(n_725),
.B(n_686),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_768),
.A2(n_725),
.B(n_686),
.Y(n_1022)
);

O2A1O1Ixp5_ASAP7_75t_L g1023 ( 
.A1(n_822),
.A2(n_540),
.B(n_522),
.C(n_521),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_779),
.A2(n_725),
.B1(n_686),
.B2(n_692),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_908),
.A2(n_912),
.B(n_906),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_879),
.B(n_686),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_895),
.B(n_250),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_908),
.A2(n_725),
.B(n_669),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_823),
.A2(n_315),
.B(n_308),
.Y(n_1029)
);

BUFx4f_ASAP7_75t_L g1030 ( 
.A(n_891),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_831),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_859),
.A2(n_875),
.B(n_906),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_893),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_912),
.A2(n_698),
.B(n_654),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_863),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_827),
.A2(n_725),
.B(n_669),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_899),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_796),
.A2(n_396),
.B(n_328),
.C(n_327),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_834),
.A2(n_692),
.B(n_605),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_780),
.B(n_250),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_777),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_835),
.A2(n_396),
.B(n_328),
.C(n_329),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_888),
.B(n_521),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_891),
.B(n_698),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_789),
.A2(n_654),
.B1(n_698),
.B2(n_370),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_836),
.A2(n_654),
.B(n_698),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_832),
.B(n_521),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_832),
.B(n_654),
.Y(n_1048)
);

OAI21xp33_ASAP7_75t_L g1049 ( 
.A1(n_790),
.A2(n_332),
.B(n_319),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_837),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_844),
.A2(n_363),
.B(n_309),
.C(n_387),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_782),
.B(n_532),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_832),
.B(n_517),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_832),
.B(n_517),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_897),
.B(n_323),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_772),
.A2(n_810),
.B(n_782),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_778),
.B(n_532),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_832),
.B(n_884),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_788),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_884),
.B(n_517),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_849),
.A2(n_538),
.B(n_532),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_853),
.A2(n_538),
.B(n_532),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_889),
.A2(n_538),
.B(n_517),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_847),
.B(n_290),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_889),
.A2(n_538),
.B(n_211),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_807),
.A2(n_379),
.B(n_351),
.C(n_388),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_815),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_884),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_785),
.B(n_538),
.Y(n_1069)
);

BUFx12f_ASAP7_75t_L g1070 ( 
.A(n_884),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_833),
.A2(n_845),
.B(n_848),
.C(n_838),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_884),
.B(n_309),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_901),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_901),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_809),
.A2(n_347),
.B1(n_357),
.B2(n_360),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_845),
.B(n_351),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_848),
.A2(n_399),
.B(n_369),
.C(n_370),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_857),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_843),
.B(n_316),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_857),
.A2(n_399),
.B(n_369),
.C(n_373),
.Y(n_1080)
);

AO21x1_ASAP7_75t_L g1081 ( 
.A1(n_855),
.A2(n_375),
.B(n_373),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_864),
.B(n_375),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_864),
.B(n_316),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_915),
.B(n_333),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_800),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_867),
.A2(n_213),
.B(n_210),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_786),
.B(n_327),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_SL g1088 ( 
.A(n_831),
.B(n_323),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_SL g1089 ( 
.A1(n_867),
.A2(n_388),
.B(n_379),
.C(n_390),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_873),
.B(n_335),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_873),
.A2(n_216),
.B(n_214),
.Y(n_1091)
);

AO21x1_ASAP7_75t_L g1092 ( 
.A1(n_813),
.A2(n_898),
.B(n_881),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_881),
.A2(n_898),
.B(n_911),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_903),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_852),
.B(n_383),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_852),
.B(n_794),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_921),
.Y(n_1097)
);

AOI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1010),
.A2(n_803),
.B(n_794),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_1030),
.B(n_886),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1059),
.B(n_803),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_993),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1064),
.A2(n_882),
.B1(n_896),
.B2(n_894),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_923),
.B(n_862),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_925),
.B(n_840),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_968),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1008),
.B(n_840),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_974),
.A2(n_911),
.B(n_854),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_SL g1108 ( 
.A(n_967),
.B(n_1029),
.C(n_342),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_957),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_917),
.A2(n_854),
.B(n_851),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_1030),
.B(n_886),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_922),
.B(n_886),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1002),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_952),
.B(n_851),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_918),
.B(n_323),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1084),
.A2(n_386),
.B1(n_339),
.B2(n_343),
.Y(n_1116)
);

NAND2x1_ASAP7_75t_L g1117 ( 
.A(n_1068),
.B(n_865),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1042),
.A2(n_390),
.B(n_389),
.C(n_395),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_919),
.A2(n_866),
.B(n_865),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_922),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_936),
.A2(n_965),
.B(n_1025),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1041),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1014),
.Y(n_1123)
);

BUFx8_ASAP7_75t_L g1124 ( 
.A(n_1085),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_964),
.B(n_1033),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_1014),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_941),
.A2(n_896),
.B(n_894),
.C(n_892),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1000),
.A2(n_877),
.B(n_866),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1084),
.A2(n_382),
.B1(n_353),
.B2(n_372),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1040),
.B(n_877),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_920),
.A2(n_890),
.B(n_882),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1051),
.A2(n_389),
.B(n_395),
.C(n_890),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_964),
.B(n_892),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_932),
.A2(n_549),
.B(n_543),
.C(n_870),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_942),
.A2(n_549),
.B(n_543),
.C(n_885),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1037),
.B(n_358),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1005),
.Y(n_1137)
);

NAND2x1p5_ASAP7_75t_L g1138 ( 
.A(n_1068),
.B(n_543),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_942),
.A2(n_549),
.B(n_543),
.C(n_313),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_SL g1140 ( 
.A1(n_923),
.A2(n_361),
.B1(n_364),
.B2(n_367),
.Y(n_1140)
);

OAI21xp33_ASAP7_75t_L g1141 ( 
.A1(n_1075),
.A2(n_393),
.B(n_401),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1073),
.B(n_368),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1093),
.A2(n_550),
.B(n_543),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_933),
.A2(n_300),
.B(n_304),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1021),
.A2(n_300),
.B(n_304),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1094),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_921),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1001),
.A2(n_398),
.B1(n_371),
.B2(n_405),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_982),
.B(n_374),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1001),
.A2(n_392),
.B1(n_384),
.B2(n_381),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1050),
.A2(n_313),
.B(n_550),
.C(n_380),
.Y(n_1151)
);

AOI21xp33_ASAP7_75t_L g1152 ( 
.A1(n_961),
.A2(n_377),
.B(n_397),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_941),
.A2(n_397),
.B(n_550),
.C(n_404),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_SL g1154 ( 
.A1(n_958),
.A2(n_268),
.B1(n_266),
.B2(n_264),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1073),
.B(n_323),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1074),
.B(n_1006),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_949),
.B(n_17),
.Y(n_1157)
);

AOI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1010),
.A2(n_586),
.B(n_219),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_1017),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_948),
.A2(n_219),
.B(n_366),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_981),
.B(n_20),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1032),
.A2(n_586),
.B(n_366),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1027),
.B(n_218),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_916),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1011),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_978),
.A2(n_294),
.B1(n_400),
.B2(n_391),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_989),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_924),
.B(n_21),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_982),
.B(n_227),
.Y(n_1169)
);

AOI21x1_ASAP7_75t_L g1170 ( 
.A1(n_929),
.A2(n_586),
.B(n_366),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_921),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1012),
.B(n_231),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_928),
.B(n_22),
.Y(n_1173)
);

BUFx12f_ASAP7_75t_L g1174 ( 
.A(n_972),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1012),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_973),
.A2(n_366),
.B(n_378),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_943),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_978),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1057),
.A2(n_287),
.B(n_239),
.C(n_359),
.Y(n_1179)
);

OR2x6_ASAP7_75t_L g1180 ( 
.A(n_1070),
.B(n_366),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_944),
.B(n_23),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_945),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_956),
.Y(n_1183)
);

OR2x6_ASAP7_75t_SL g1184 ( 
.A(n_1087),
.B(n_237),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_SL g1185 ( 
.A1(n_1020),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_1185)
);

O2A1O1Ixp5_ASAP7_75t_L g1186 ( 
.A1(n_1023),
.A2(n_586),
.B(n_26),
.C(n_27),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1055),
.B(n_25),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1057),
.A2(n_318),
.B(n_355),
.C(n_350),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1015),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_SL g1190 ( 
.A(n_939),
.B(n_1088),
.C(n_1095),
.Y(n_1190)
);

AOI22x1_ASAP7_75t_L g1191 ( 
.A1(n_947),
.A2(n_262),
.B1(n_272),
.B2(n_277),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1015),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_983),
.B(n_280),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_927),
.A2(n_1004),
.B(n_931),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_SL g1195 ( 
.A1(n_1079),
.A2(n_281),
.B1(n_282),
.B2(n_284),
.Y(n_1195)
);

NOR2xp67_ASAP7_75t_L g1196 ( 
.A(n_1009),
.B(n_291),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_983),
.B(n_325),
.Y(n_1197)
);

INVx4_ASAP7_75t_L g1198 ( 
.A(n_983),
.Y(n_1198)
);

BUFx8_ASAP7_75t_L g1199 ( 
.A(n_983),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1028),
.A2(n_586),
.B(n_160),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_921),
.Y(n_1201)
);

BUFx10_ASAP7_75t_L g1202 ( 
.A(n_980),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_980),
.B(n_338),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1044),
.B(n_348),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_1072),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_951),
.A2(n_345),
.B(n_344),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1023),
.A2(n_586),
.B(n_33),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_985),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_SL g1209 ( 
.A1(n_1056),
.A2(n_1065),
.B(n_1069),
.C(n_999),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_950),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_950),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1003),
.B(n_36),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1044),
.A2(n_586),
.B1(n_37),
.B2(n_38),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_976),
.A2(n_977),
.B(n_1013),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_934),
.A2(n_586),
.B(n_38),
.C(n_39),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1066),
.A2(n_36),
.B(n_40),
.C(n_42),
.Y(n_1216)
);

OAI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1049),
.A2(n_40),
.B(n_44),
.Y(n_1217)
);

CKINVDCx16_ASAP7_75t_R g1218 ( 
.A(n_946),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1015),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_950),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_997),
.A2(n_586),
.B(n_47),
.C(n_48),
.Y(n_1221)
);

AO32x1_ASAP7_75t_L g1222 ( 
.A1(n_1018),
.A2(n_45),
.A3(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_954),
.A2(n_1077),
.B(n_1080),
.C(n_990),
.Y(n_1223)
);

INVx8_ASAP7_75t_L g1224 ( 
.A(n_950),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_959),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1058),
.B(n_52),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1026),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_R g1228 ( 
.A(n_959),
.B(n_116),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_984),
.A2(n_53),
.B(n_54),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1067),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1078),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_963),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_1232)
);

INVxp67_ASAP7_75t_L g1233 ( 
.A(n_1096),
.Y(n_1233)
);

CKINVDCx16_ASAP7_75t_R g1234 ( 
.A(n_946),
.Y(n_1234)
);

BUFx12f_ASAP7_75t_L g1235 ( 
.A(n_1015),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_962),
.B(n_57),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_962),
.B(n_59),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1022),
.A2(n_59),
.B(n_60),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1083),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1009),
.B(n_60),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1090),
.B(n_61),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_960),
.A2(n_62),
.B(n_63),
.C(n_66),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1035),
.B(n_68),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1016),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_955),
.A2(n_1069),
.B(n_988),
.C(n_1038),
.Y(n_1245)
);

NAND2x1_ASAP7_75t_L g1246 ( 
.A(n_995),
.B(n_1031),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_969),
.B(n_71),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1071),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1076),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_987),
.B(n_72),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1035),
.Y(n_1251)
);

AND2x6_ASAP7_75t_SL g1252 ( 
.A(n_1047),
.B(n_74),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1076),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_1007),
.A2(n_81),
.B(n_90),
.C(n_94),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1167),
.Y(n_1255)
);

INVx5_ASAP7_75t_SL g1256 ( 
.A(n_1180),
.Y(n_1256)
);

BUFx2_ASAP7_75t_R g1257 ( 
.A(n_1184),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1214),
.A2(n_1019),
.B(n_986),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1244),
.B(n_1043),
.Y(n_1259)
);

AOI21xp33_ASAP7_75t_L g1260 ( 
.A1(n_1151),
.A2(n_963),
.B(n_1081),
.Y(n_1260)
);

BUFx12f_ASAP7_75t_L g1261 ( 
.A(n_1124),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1239),
.B(n_1082),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1214),
.A2(n_992),
.B(n_1036),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1124),
.Y(n_1264)
);

INVx6_ASAP7_75t_SL g1265 ( 
.A(n_1180),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_SL g1266 ( 
.A1(n_1209),
.A2(n_1020),
.B(n_991),
.C(n_971),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1174),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1194),
.A2(n_1062),
.B(n_1061),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1101),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1109),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1150),
.A2(n_1089),
.B(n_991),
.C(n_971),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1114),
.B(n_1082),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1235),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1120),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1216),
.A2(n_1089),
.B(n_1091),
.C(n_1086),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1233),
.B(n_937),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1137),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1123),
.B(n_1126),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1245),
.A2(n_979),
.B(n_1039),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1146),
.B(n_1156),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1163),
.A2(n_926),
.B1(n_970),
.B2(n_1024),
.Y(n_1281)
);

AOI31xp67_ASAP7_75t_L g1282 ( 
.A1(n_1226),
.A2(n_996),
.A3(n_935),
.B(n_938),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1178),
.B(n_940),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1104),
.B(n_926),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1160),
.A2(n_1053),
.B(n_1060),
.Y(n_1285)
);

AOI221xp5_ASAP7_75t_SL g1286 ( 
.A1(n_1165),
.A2(n_994),
.B1(n_998),
.B2(n_953),
.C(n_1052),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1164),
.Y(n_1287)
);

O2A1O1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1216),
.A2(n_938),
.B(n_935),
.C(n_1052),
.Y(n_1288)
);

INVxp67_ASAP7_75t_SL g1289 ( 
.A(n_1100),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1115),
.B(n_1054),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1159),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1223),
.A2(n_996),
.B(n_975),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1182),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1160),
.A2(n_1092),
.A3(n_1063),
.B(n_1046),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1232),
.A2(n_995),
.B1(n_1035),
.B2(n_1045),
.Y(n_1295)
);

AO31x2_ASAP7_75t_L g1296 ( 
.A1(n_1119),
.A2(n_1048),
.A3(n_1034),
.B(n_930),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1110),
.A2(n_1031),
.B(n_1035),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1183),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1208),
.Y(n_1299)
);

O2A1O1Ixp5_ASAP7_75t_L g1300 ( 
.A1(n_1207),
.A2(n_106),
.B(n_108),
.C(n_112),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1233),
.B(n_118),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1125),
.A2(n_1242),
.B1(n_1212),
.B2(n_1247),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1107),
.A2(n_119),
.B(n_120),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1202),
.B(n_121),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1231),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1120),
.B(n_122),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1203),
.A2(n_138),
.B1(n_146),
.B2(n_157),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1107),
.A2(n_159),
.B(n_162),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1118),
.A2(n_164),
.B(n_170),
.C(n_171),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1106),
.B(n_176),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1110),
.A2(n_179),
.B(n_186),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1227),
.A2(n_194),
.B(n_197),
.C(n_204),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1202),
.B(n_207),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1131),
.A2(n_1162),
.B(n_1098),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1131),
.A2(n_1119),
.B(n_1143),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1217),
.B(n_1165),
.C(n_1215),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_SL g1317 ( 
.A1(n_1246),
.A2(n_1179),
.B(n_1188),
.C(n_1254),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1127),
.A2(n_1176),
.A3(n_1248),
.B(n_1128),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1199),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1218),
.B(n_1234),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1118),
.A2(n_1130),
.B(n_1151),
.C(n_1108),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1223),
.A2(n_1186),
.B(n_1139),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1205),
.B(n_1142),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1175),
.B(n_1220),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1176),
.A2(n_1128),
.A3(n_1145),
.B(n_1144),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1108),
.B(n_1169),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1199),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1105),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1221),
.A2(n_1173),
.B1(n_1168),
.B2(n_1181),
.Y(n_1329)
);

AOI31xp67_ASAP7_75t_L g1330 ( 
.A1(n_1250),
.A2(n_1243),
.A3(n_1237),
.B(n_1236),
.Y(n_1330)
);

NOR2x1_ASAP7_75t_SL g1331 ( 
.A(n_1097),
.B(n_1147),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1139),
.A2(n_1180),
.B(n_1190),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1172),
.B(n_1155),
.Y(n_1333)
);

NAND3xp33_ASAP7_75t_L g1334 ( 
.A(n_1238),
.B(n_1229),
.C(n_1132),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1230),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1132),
.A2(n_1190),
.B(n_1241),
.C(n_1152),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1103),
.B(n_1099),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1141),
.A2(n_1136),
.B(n_1149),
.C(n_1185),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1113),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1103),
.B(n_1111),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1122),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1133),
.B(n_1253),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1186),
.A2(n_1229),
.B(n_1135),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1144),
.A2(n_1206),
.B(n_1117),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1200),
.A2(n_1170),
.B(n_1158),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1153),
.A2(n_1249),
.B(n_1148),
.C(n_1206),
.Y(n_1346)
);

O2A1O1Ixp5_ASAP7_75t_SL g1347 ( 
.A1(n_1193),
.A2(n_1197),
.B(n_1211),
.C(n_1240),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1140),
.B(n_1154),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1196),
.A2(n_1238),
.B(n_1187),
.C(n_1157),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1210),
.B(n_1112),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1177),
.B(n_1225),
.Y(n_1351)
);

AO31x2_ASAP7_75t_L g1352 ( 
.A1(n_1198),
.A2(n_1222),
.A3(n_1135),
.B(n_1134),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1251),
.B(n_1097),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1097),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1116),
.A2(n_1129),
.B(n_1213),
.C(n_1161),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1102),
.B(n_1171),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1147),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1147),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1134),
.A2(n_1138),
.B(n_1222),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1171),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1171),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1201),
.B(n_1219),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1166),
.B(n_1224),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1224),
.B(n_1204),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1138),
.A2(n_1222),
.B(n_1191),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1224),
.Y(n_1366)
);

O2A1O1Ixp5_ASAP7_75t_L g1367 ( 
.A1(n_1189),
.A2(n_1192),
.B(n_1252),
.C(n_1195),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1201),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1201),
.Y(n_1369)
);

OAI22x1_ASAP7_75t_L g1370 ( 
.A1(n_1228),
.A2(n_562),
.B1(n_981),
.B2(n_679),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1214),
.A2(n_1000),
.B(n_1160),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1214),
.A2(n_1000),
.B(n_1160),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1239),
.B(n_814),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1101),
.Y(n_1374)
);

AO31x2_ASAP7_75t_L g1375 ( 
.A1(n_1160),
.A2(n_966),
.A3(n_1092),
.B(n_1081),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1232),
.A2(n_1001),
.B1(n_952),
.B2(n_1008),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1121),
.A2(n_1214),
.B(n_1194),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1232),
.A2(n_1001),
.B1(n_952),
.B2(n_1008),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1239),
.B(n_814),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1160),
.A2(n_966),
.A3(n_1092),
.B(n_1081),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_SL g1381 ( 
.A1(n_1209),
.A2(n_812),
.B(n_1246),
.C(n_1188),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1167),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1121),
.A2(n_1214),
.B(n_1194),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1123),
.B(n_606),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1123),
.B(n_1059),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1123),
.B(n_606),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1202),
.B(n_625),
.Y(n_1387)
);

AO31x2_ASAP7_75t_L g1388 ( 
.A1(n_1160),
.A2(n_966),
.A3(n_1092),
.B(n_1081),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1101),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1214),
.A2(n_1000),
.B(n_1160),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1123),
.B(n_625),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1231),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1121),
.A2(n_1214),
.B(n_1194),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1121),
.A2(n_1214),
.B(n_1194),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1214),
.A2(n_1000),
.B(n_1160),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1121),
.A2(n_1214),
.B(n_1194),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1174),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1160),
.A2(n_1098),
.B(n_1119),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1239),
.B(n_814),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1245),
.A2(n_1023),
.B(n_1223),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1231),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1120),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1231),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1101),
.Y(n_1404)
);

AOI221xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1165),
.A2(n_1216),
.B1(n_1227),
.B2(n_1217),
.C(n_1118),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1214),
.A2(n_1000),
.B(n_1160),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1120),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1120),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1120),
.Y(n_1409)
);

AO21x1_ASAP7_75t_L g1410 ( 
.A1(n_1160),
.A2(n_1151),
.B(n_1010),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1214),
.A2(n_1000),
.B(n_1160),
.Y(n_1411)
);

OA21x2_ASAP7_75t_L g1412 ( 
.A1(n_1194),
.A2(n_1160),
.B(n_1214),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1245),
.A2(n_1023),
.B(n_1223),
.Y(n_1413)
);

CKINVDCx8_ASAP7_75t_R g1414 ( 
.A(n_1167),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1101),
.Y(n_1415)
);

NAND3x1_ASAP7_75t_L g1416 ( 
.A(n_1161),
.B(n_1084),
.C(n_826),
.Y(n_1416)
);

AOI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1160),
.A2(n_1214),
.B(n_1194),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_SL g1418 ( 
.A1(n_1209),
.A2(n_812),
.B(n_1246),
.C(n_1188),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1121),
.A2(n_1214),
.B(n_1194),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1245),
.A2(n_1023),
.B(n_1223),
.Y(n_1420)
);

AO31x2_ASAP7_75t_L g1421 ( 
.A1(n_1160),
.A2(n_966),
.A3(n_1092),
.B(n_1081),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1231),
.Y(n_1422)
);

NAND3xp33_ASAP7_75t_L g1423 ( 
.A(n_1232),
.B(n_825),
.C(n_1216),
.Y(n_1423)
);

OR2x6_ASAP7_75t_L g1424 ( 
.A(n_1120),
.B(n_943),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1423),
.A2(n_1370),
.B1(n_1376),
.B2(n_1378),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1355),
.A2(n_1333),
.B1(n_1423),
.B2(n_1281),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1316),
.A2(n_1348),
.B1(n_1376),
.B2(n_1378),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1316),
.A2(n_1391),
.B1(n_1336),
.B2(n_1399),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1269),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1326),
.A2(n_1329),
.B1(n_1373),
.B2(n_1379),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1289),
.B(n_1323),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1284),
.A2(n_1302),
.B1(n_1329),
.B2(n_1257),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1277),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1302),
.A2(n_1260),
.B1(n_1386),
.B2(n_1384),
.Y(n_1434)
);

CKINVDCx6p67_ASAP7_75t_R g1435 ( 
.A(n_1261),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1334),
.A2(n_1321),
.B1(n_1349),
.B2(n_1346),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1416),
.A2(n_1405),
.B1(n_1340),
.B2(n_1337),
.Y(n_1437)
);

INVx8_ASAP7_75t_L g1438 ( 
.A(n_1424),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1368),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1374),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1412),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1270),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1260),
.A2(n_1262),
.B1(n_1290),
.B2(n_1334),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1280),
.A2(n_1301),
.B1(n_1351),
.B2(n_1389),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1412),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1414),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1322),
.A2(n_1413),
.B1(n_1400),
.B2(n_1420),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1278),
.A2(n_1387),
.B1(n_1420),
.B2(n_1413),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1404),
.Y(n_1449)
);

BUFx4f_ASAP7_75t_SL g1450 ( 
.A(n_1255),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1382),
.Y(n_1451)
);

CKINVDCx11_ASAP7_75t_R g1452 ( 
.A(n_1267),
.Y(n_1452)
);

INVx4_ASAP7_75t_L g1453 ( 
.A(n_1327),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1322),
.A2(n_1400),
.B1(n_1422),
.B2(n_1401),
.Y(n_1454)
);

AOI22x1_ASAP7_75t_SL g1455 ( 
.A1(n_1264),
.A2(n_1291),
.B1(n_1408),
.B2(n_1402),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1392),
.A2(n_1403),
.B1(n_1259),
.B2(n_1415),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1328),
.A2(n_1339),
.B1(n_1341),
.B2(n_1337),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1287),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1293),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1298),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_SL g1461 ( 
.A1(n_1256),
.A2(n_1343),
.B1(n_1301),
.B2(n_1405),
.Y(n_1461)
);

OAI22xp33_ASAP7_75t_R g1462 ( 
.A1(n_1385),
.A2(n_1299),
.B1(n_1335),
.B2(n_1283),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1343),
.A2(n_1363),
.B1(n_1338),
.B2(n_1276),
.Y(n_1463)
);

OAI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1276),
.A2(n_1307),
.B1(n_1424),
.B2(n_1272),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1367),
.B(n_1274),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1342),
.Y(n_1466)
);

BUFx4f_ASAP7_75t_SL g1467 ( 
.A(n_1397),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1377),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1340),
.A2(n_1259),
.B1(n_1265),
.B2(n_1356),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1256),
.A2(n_1324),
.B1(n_1310),
.B2(n_1306),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1319),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1410),
.A2(n_1342),
.B1(n_1324),
.B2(n_1350),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1402),
.A2(n_1408),
.B1(n_1309),
.B2(n_1409),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1274),
.A2(n_1409),
.B1(n_1407),
.B2(n_1332),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1383),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1407),
.A2(n_1320),
.B1(n_1275),
.B2(n_1424),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1304),
.A2(n_1313),
.B1(n_1350),
.B2(n_1306),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1358),
.B(n_1360),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1368),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1362),
.B(n_1366),
.Y(n_1480)
);

CKINVDCx11_ASAP7_75t_R g1481 ( 
.A(n_1357),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1354),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1310),
.A2(n_1295),
.B1(n_1364),
.B2(n_1292),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1271),
.A2(n_1371),
.B1(n_1411),
.B2(n_1406),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1361),
.B(n_1369),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1372),
.A2(n_1390),
.B1(n_1395),
.B2(n_1359),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1331),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1295),
.A2(n_1292),
.B1(n_1365),
.B2(n_1285),
.Y(n_1488)
);

INVx6_ASAP7_75t_L g1489 ( 
.A(n_1347),
.Y(n_1489)
);

INVx3_ASAP7_75t_SL g1490 ( 
.A(n_1330),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1282),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_1279),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1311),
.A2(n_1308),
.B1(n_1303),
.B2(n_1300),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1312),
.A2(n_1279),
.B1(n_1344),
.B2(n_1258),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_1297),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1398),
.A2(n_1263),
.B1(n_1268),
.B2(n_1314),
.Y(n_1496)
);

BUFx8_ASAP7_75t_L g1497 ( 
.A(n_1381),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1288),
.A2(n_1417),
.B1(n_1418),
.B2(n_1266),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1352),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1352),
.B(n_1318),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1317),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1296),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1318),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1286),
.A2(n_1345),
.B1(n_1315),
.B2(n_1396),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1393),
.A2(n_1419),
.B1(n_1394),
.B2(n_1421),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1286),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1318),
.A2(n_1325),
.B1(n_1296),
.B2(n_1375),
.Y(n_1507)
);

INVx6_ASAP7_75t_L g1508 ( 
.A(n_1296),
.Y(n_1508)
);

AOI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1375),
.A2(n_1380),
.B1(n_1388),
.B2(n_1421),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1375),
.A2(n_1380),
.B1(n_1388),
.B2(n_1421),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1380),
.A2(n_1388),
.B1(n_1325),
.B2(n_1294),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1325),
.A2(n_915),
.B1(n_716),
.B2(n_410),
.Y(n_1512)
);

OAI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1423),
.A2(n_1281),
.B1(n_1378),
.B2(n_1376),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1355),
.A2(n_1333),
.B1(n_1001),
.B2(n_1423),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1255),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_SL g1517 ( 
.A1(n_1423),
.A2(n_915),
.B1(n_716),
.B2(n_410),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1305),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1305),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1348),
.A2(n_1370),
.B1(n_679),
.B2(n_729),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1348),
.A2(n_1084),
.B1(n_625),
.B2(n_850),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1384),
.B(n_1386),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1355),
.A2(n_1333),
.B1(n_1001),
.B2(n_1423),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1355),
.A2(n_1333),
.B1(n_1001),
.B2(n_1423),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1278),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_1255),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1255),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1423),
.A2(n_825),
.B(n_1302),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_SL g1531 ( 
.A1(n_1348),
.A2(n_1370),
.B1(n_679),
.B2(n_729),
.Y(n_1531)
);

CKINVDCx11_ASAP7_75t_R g1532 ( 
.A(n_1414),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1533)
);

CKINVDCx11_ASAP7_75t_R g1534 ( 
.A(n_1414),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1348),
.A2(n_1355),
.B(n_1084),
.Y(n_1535)
);

OAI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1423),
.A2(n_1281),
.B1(n_1378),
.B2(n_1376),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1537)
);

BUFx12f_ASAP7_75t_L g1538 ( 
.A(n_1261),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1539)
);

BUFx2_ASAP7_75t_SL g1540 ( 
.A(n_1255),
.Y(n_1540)
);

BUFx12f_ASAP7_75t_L g1541 ( 
.A(n_1261),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1542)
);

BUFx10_ASAP7_75t_L g1543 ( 
.A(n_1327),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1270),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1269),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1305),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_SL g1550 ( 
.A1(n_1423),
.A2(n_915),
.B1(n_716),
.B2(n_410),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_1255),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1373),
.B(n_1379),
.Y(n_1553)
);

INVx5_ASAP7_75t_L g1554 ( 
.A(n_1424),
.Y(n_1554)
);

CKINVDCx14_ASAP7_75t_R g1555 ( 
.A(n_1255),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1368),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1353),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1423),
.A2(n_1281),
.B1(n_1378),
.B2(n_1376),
.Y(n_1559)
);

CKINVDCx11_ASAP7_75t_R g1560 ( 
.A(n_1414),
.Y(n_1560)
);

INVx6_ASAP7_75t_L g1561 ( 
.A(n_1273),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1270),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_1255),
.Y(n_1564)
);

CKINVDCx11_ASAP7_75t_R g1565 ( 
.A(n_1414),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1423),
.A2(n_1281),
.B1(n_1378),
.B2(n_1376),
.Y(n_1566)
);

CKINVDCx11_ASAP7_75t_R g1567 ( 
.A(n_1414),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1353),
.B(n_1337),
.Y(n_1568)
);

INVx4_ASAP7_75t_L g1569 ( 
.A(n_1327),
.Y(n_1569)
);

INVx6_ASAP7_75t_L g1570 ( 
.A(n_1273),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1355),
.A2(n_1333),
.B1(n_1001),
.B2(n_1423),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1423),
.A2(n_915),
.B1(n_716),
.B2(n_410),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1423),
.A2(n_852),
.B1(n_1370),
.B2(n_981),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1442),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1466),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1446),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1532),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1427),
.A2(n_1535),
.B1(n_1447),
.B2(n_1522),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1491),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1429),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1554),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1544),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1492),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1530),
.A2(n_1524),
.B(n_1514),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1433),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1526),
.A2(n_1571),
.B(n_1426),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1440),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1562),
.Y(n_1588)
);

NOR2x1_ASAP7_75t_R g1589 ( 
.A(n_1534),
.B(n_1560),
.Y(n_1589)
);

OR2x6_ASAP7_75t_L g1590 ( 
.A(n_1438),
.B(n_1508),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1554),
.Y(n_1591)
);

OAI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1513),
.A2(n_1559),
.B1(n_1536),
.B2(n_1566),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1447),
.B(n_1506),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1431),
.B(n_1500),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1527),
.B(n_1450),
.Y(n_1595)
);

OA21x2_ASAP7_75t_L g1596 ( 
.A1(n_1496),
.A2(n_1511),
.B(n_1510),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1523),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1481),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1448),
.B(n_1443),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1449),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1458),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1443),
.B(n_1503),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1459),
.B(n_1460),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1428),
.A2(n_1436),
.B(n_1513),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1511),
.B(n_1425),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1554),
.B(n_1502),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1536),
.A2(n_1566),
.B(n_1559),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1484),
.A2(n_1496),
.B(n_1486),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1545),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1495),
.B(n_1568),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1441),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1441),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1438),
.Y(n_1613)
);

AO21x2_ASAP7_75t_L g1614 ( 
.A1(n_1509),
.A2(n_1507),
.B(n_1504),
.Y(n_1614)
);

NAND2x1p5_ASAP7_75t_L g1615 ( 
.A(n_1487),
.B(n_1437),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1438),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1498),
.A2(n_1505),
.B(n_1488),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1445),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1445),
.Y(n_1619)
);

AO31x2_ASAP7_75t_L g1620 ( 
.A1(n_1463),
.A2(n_1519),
.A3(n_1547),
.B(n_1518),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1485),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1499),
.B(n_1454),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1553),
.B(n_1430),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1490),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1468),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1490),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1468),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1497),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1425),
.B(n_1478),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1475),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1454),
.B(n_1434),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1510),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1456),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1489),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1456),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1489),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1489),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1434),
.B(n_1483),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1558),
.B(n_1444),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_SL g1640 ( 
.A(n_1538),
.B(n_1541),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1488),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1497),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1472),
.Y(n_1643)
);

INVx4_ASAP7_75t_L g1644 ( 
.A(n_1439),
.Y(n_1644)
);

BUFx2_ASAP7_75t_SL g1645 ( 
.A(n_1501),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1479),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_SL g1647 ( 
.A1(n_1476),
.A2(n_1474),
.B(n_1473),
.Y(n_1647)
);

NOR2x1_ASAP7_75t_R g1648 ( 
.A(n_1565),
.B(n_1567),
.Y(n_1648)
);

AO21x1_ASAP7_75t_L g1649 ( 
.A1(n_1464),
.A2(n_1465),
.B(n_1432),
.Y(n_1649)
);

NAND2x1_ASAP7_75t_L g1650 ( 
.A(n_1483),
.B(n_1482),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1461),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1494),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1464),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1556),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1450),
.B(n_1528),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1457),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1480),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1462),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1469),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1515),
.B(n_1537),
.Y(n_1660)
);

BUFx2_ASAP7_75t_L g1661 ( 
.A(n_1561),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1512),
.A2(n_1572),
.B1(n_1550),
.B2(n_1517),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1477),
.B(n_1569),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1470),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1493),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1515),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1520),
.B(n_1573),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1520),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1516),
.B(n_1529),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1525),
.B(n_1573),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1525),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1533),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1533),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1537),
.A2(n_1548),
.B(n_1546),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1570),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1539),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1539),
.B(n_1548),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1453),
.B(n_1569),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1471),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1594),
.B(n_1540),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1583),
.B(n_1555),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1583),
.B(n_1453),
.Y(n_1682)
);

AOI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1578),
.A2(n_1552),
.B1(n_1549),
.B2(n_1546),
.C(n_1557),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1646),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1611),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1608),
.A2(n_1542),
.B(n_1563),
.Y(n_1686)
);

O2A1O1Ixp33_ASAP7_75t_SL g1687 ( 
.A1(n_1592),
.A2(n_1564),
.B(n_1551),
.C(n_1455),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1597),
.B(n_1543),
.Y(n_1688)
);

A2O1A1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1604),
.A2(n_1557),
.B(n_1552),
.C(n_1549),
.Y(n_1689)
);

OA21x2_ASAP7_75t_L g1690 ( 
.A1(n_1608),
.A2(n_1563),
.B(n_1542),
.Y(n_1690)
);

OA21x2_ASAP7_75t_L g1691 ( 
.A1(n_1617),
.A2(n_1521),
.B(n_1531),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1590),
.B(n_1451),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1590),
.B(n_1467),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1590),
.B(n_1467),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1575),
.B(n_1435),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1580),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1646),
.B(n_1452),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1574),
.Y(n_1698)
);

AO32x2_ASAP7_75t_L g1699 ( 
.A1(n_1581),
.A2(n_1591),
.A3(n_1644),
.B1(n_1594),
.B2(n_1616),
.Y(n_1699)
);

AND2x6_ASAP7_75t_L g1700 ( 
.A(n_1638),
.B(n_1606),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1593),
.B(n_1641),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1607),
.A2(n_1584),
.B(n_1586),
.Y(n_1702)
);

OA21x2_ASAP7_75t_L g1703 ( 
.A1(n_1617),
.A2(n_1626),
.B(n_1665),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1611),
.Y(n_1704)
);

AOI221x1_ASAP7_75t_SL g1705 ( 
.A1(n_1658),
.A2(n_1667),
.B1(n_1623),
.B2(n_1652),
.C(n_1607),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1576),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1603),
.B(n_1657),
.Y(n_1707)
);

OA21x2_ASAP7_75t_L g1708 ( 
.A1(n_1626),
.A2(n_1665),
.B(n_1636),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_SL g1709 ( 
.A(n_1649),
.B(n_1599),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1661),
.Y(n_1710)
);

AOI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1638),
.A2(n_1649),
.B1(n_1599),
.B2(n_1660),
.C(n_1670),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1576),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1652),
.B(n_1593),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1610),
.B(n_1645),
.Y(n_1714)
);

AOI221xp5_ASAP7_75t_L g1715 ( 
.A1(n_1660),
.A2(n_1670),
.B1(n_1677),
.B2(n_1676),
.C(n_1673),
.Y(n_1715)
);

NAND2x1_ASAP7_75t_L g1716 ( 
.A(n_1647),
.B(n_1663),
.Y(n_1716)
);

AO21x2_ASAP7_75t_L g1717 ( 
.A1(n_1634),
.A2(n_1637),
.B(n_1636),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1677),
.A2(n_1674),
.B1(n_1631),
.B2(n_1662),
.Y(n_1718)
);

A2O1A1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1631),
.A2(n_1651),
.B(n_1653),
.C(n_1658),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1653),
.A2(n_1641),
.B(n_1674),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1577),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1621),
.B(n_1609),
.Y(n_1722)
);

NAND3xp33_ASAP7_75t_L g1723 ( 
.A(n_1666),
.B(n_1673),
.C(n_1671),
.Y(n_1723)
);

A2O1A1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1651),
.A2(n_1668),
.B(n_1666),
.C(n_1676),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1674),
.A2(n_1671),
.B1(n_1672),
.B2(n_1668),
.Y(n_1725)
);

O2A1O1Ixp33_ASAP7_75t_SL g1726 ( 
.A1(n_1650),
.A2(n_1628),
.B(n_1598),
.C(n_1595),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1585),
.B(n_1587),
.Y(n_1727)
);

CKINVDCx16_ASAP7_75t_R g1728 ( 
.A(n_1640),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1663),
.B(n_1650),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1582),
.B(n_1588),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1588),
.B(n_1654),
.Y(n_1731)
);

INVx5_ASAP7_75t_L g1732 ( 
.A(n_1624),
.Y(n_1732)
);

AO32x2_ASAP7_75t_L g1733 ( 
.A1(n_1581),
.A2(n_1591),
.A3(n_1644),
.B1(n_1616),
.B2(n_1613),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1600),
.B(n_1601),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1674),
.A2(n_1672),
.B(n_1605),
.Y(n_1735)
);

A2O1A1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1602),
.A2(n_1605),
.B(n_1664),
.C(n_1629),
.Y(n_1736)
);

AOI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1579),
.A2(n_1642),
.B(n_1678),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1642),
.A2(n_1628),
.B1(n_1664),
.B2(n_1643),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1643),
.A2(n_1679),
.B1(n_1615),
.B2(n_1602),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1620),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1659),
.A2(n_1656),
.B1(n_1633),
.B2(n_1635),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_SL g1742 ( 
.A1(n_1577),
.A2(n_1669),
.B1(n_1655),
.B2(n_1678),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1612),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1618),
.B(n_1619),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1675),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1659),
.A2(n_1639),
.B1(n_1622),
.B2(n_1615),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1701),
.B(n_1618),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1702),
.B(n_1678),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1685),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1685),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1743),
.B(n_1579),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1707),
.B(n_1614),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1699),
.B(n_1614),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1704),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1740),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1699),
.B(n_1614),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1699),
.B(n_1703),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1704),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1711),
.A2(n_1622),
.B1(n_1632),
.B2(n_1635),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1744),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1699),
.B(n_1703),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1729),
.B(n_1596),
.Y(n_1762)
);

INVx4_ASAP7_75t_L g1763 ( 
.A(n_1693),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1696),
.B(n_1720),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1729),
.B(n_1596),
.Y(n_1765)
);

NAND3xp33_ASAP7_75t_L g1766 ( 
.A(n_1711),
.B(n_1625),
.C(n_1627),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1709),
.A2(n_1632),
.B1(n_1633),
.B2(n_1656),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1732),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1727),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1684),
.B(n_1624),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1734),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1734),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1722),
.B(n_1630),
.Y(n_1773)
);

AOI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1683),
.A2(n_1705),
.B1(n_1689),
.B2(n_1715),
.C(n_1687),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1737),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1695),
.B(n_1680),
.Y(n_1776)
);

BUFx3_ASAP7_75t_L g1777 ( 
.A(n_1700),
.Y(n_1777)
);

BUFx8_ASAP7_75t_L g1778 ( 
.A(n_1733),
.Y(n_1778)
);

AOI211xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1774),
.A2(n_1687),
.B(n_1726),
.C(n_1683),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1753),
.B(n_1710),
.Y(n_1780)
);

OAI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1759),
.A2(n_1689),
.B1(n_1718),
.B2(n_1719),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1755),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_L g1783 ( 
.A(n_1774),
.B(n_1690),
.C(n_1715),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1750),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1749),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1747),
.B(n_1745),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1749),
.Y(n_1787)
);

INVxp67_ASAP7_75t_SL g1788 ( 
.A(n_1778),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1776),
.B(n_1706),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1760),
.B(n_1735),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1760),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1754),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1753),
.B(n_1756),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1753),
.B(n_1708),
.Y(n_1794)
);

AOI221xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1764),
.A2(n_1719),
.B1(n_1736),
.B2(n_1724),
.C(n_1725),
.Y(n_1795)
);

BUFx12f_ASAP7_75t_L g1796 ( 
.A(n_1763),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1771),
.B(n_1713),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1756),
.B(n_1708),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1756),
.B(n_1731),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1777),
.B(n_1700),
.Y(n_1800)
);

AOI211xp5_ASAP7_75t_L g1801 ( 
.A1(n_1766),
.A2(n_1726),
.B(n_1736),
.C(n_1724),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1777),
.B(n_1700),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1757),
.B(n_1733),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1771),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1757),
.B(n_1761),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1758),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1758),
.Y(n_1807)
);

BUFx2_ASAP7_75t_L g1808 ( 
.A(n_1778),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1757),
.B(n_1733),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1759),
.A2(n_1691),
.B1(n_1690),
.B2(n_1713),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1761),
.B(n_1733),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1761),
.B(n_1717),
.Y(n_1812)
);

AO21x2_ASAP7_75t_L g1813 ( 
.A1(n_1766),
.A2(n_1717),
.B(n_1746),
.Y(n_1813)
);

XNOR2xp5_ASAP7_75t_L g1814 ( 
.A(n_1752),
.B(n_1681),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1767),
.A2(n_1691),
.B1(n_1723),
.B2(n_1739),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1767),
.A2(n_1716),
.B1(n_1741),
.B2(n_1738),
.Y(n_1816)
);

INVx5_ASAP7_75t_L g1817 ( 
.A(n_1768),
.Y(n_1817)
);

NAND2xp33_ASAP7_75t_SL g1818 ( 
.A(n_1763),
.B(n_1697),
.Y(n_1818)
);

NAND3xp33_ASAP7_75t_L g1819 ( 
.A(n_1764),
.B(n_1695),
.C(n_1741),
.Y(n_1819)
);

AOI211xp5_ASAP7_75t_L g1820 ( 
.A1(n_1748),
.A2(n_1686),
.B(n_1742),
.C(n_1714),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1751),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1790),
.B(n_1747),
.Y(n_1822)
);

BUFx2_ASAP7_75t_L g1823 ( 
.A(n_1796),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1803),
.B(n_1775),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1796),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1790),
.B(n_1773),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1785),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1785),
.Y(n_1828)
);

NOR3xp33_ASAP7_75t_SL g1829 ( 
.A(n_1818),
.B(n_1721),
.C(n_1712),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1803),
.B(n_1775),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1803),
.B(n_1775),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1809),
.B(n_1775),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1782),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1786),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1821),
.B(n_1769),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1817),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1809),
.B(n_1775),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1811),
.B(n_1805),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1811),
.B(n_1805),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1787),
.Y(n_1840)
);

INVx3_ASAP7_75t_L g1841 ( 
.A(n_1817),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1817),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1787),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1821),
.B(n_1769),
.Y(n_1844)
);

BUFx2_ASAP7_75t_L g1845 ( 
.A(n_1796),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1792),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1805),
.B(n_1770),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1800),
.B(n_1777),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1792),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1791),
.B(n_1772),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1780),
.B(n_1762),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1800),
.B(n_1802),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1786),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1780),
.B(n_1765),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1780),
.B(n_1765),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1804),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1806),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1799),
.B(n_1765),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1843),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1833),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1838),
.B(n_1817),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1834),
.B(n_1819),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1843),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1833),
.Y(n_1864)
);

AOI21x1_ASAP7_75t_L g1865 ( 
.A1(n_1823),
.A2(n_1807),
.B(n_1784),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1843),
.Y(n_1866)
);

AOI21xp33_ASAP7_75t_L g1867 ( 
.A1(n_1826),
.A2(n_1801),
.B(n_1795),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1827),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1827),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1838),
.B(n_1817),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1838),
.B(n_1817),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1828),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1834),
.B(n_1819),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1828),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1839),
.B(n_1852),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1823),
.B(n_1589),
.Y(n_1876)
);

OR2x2_ASAP7_75t_SL g1877 ( 
.A(n_1822),
.B(n_1728),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1840),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1822),
.B(n_1797),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1853),
.A2(n_1779),
.B(n_1783),
.Y(n_1880)
);

NOR3xp33_ASAP7_75t_L g1881 ( 
.A(n_1823),
.B(n_1783),
.C(n_1845),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_1845),
.Y(n_1882)
);

INVxp67_ASAP7_75t_SL g1883 ( 
.A(n_1856),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1853),
.B(n_1797),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1840),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1822),
.B(n_1820),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1833),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1833),
.Y(n_1888)
);

INVx2_ASAP7_75t_SL g1889 ( 
.A(n_1852),
.Y(n_1889)
);

NAND4xp25_ASAP7_75t_L g1890 ( 
.A(n_1824),
.B(n_1779),
.C(n_1801),
.D(n_1795),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1852),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1826),
.B(n_1820),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1852),
.B(n_1800),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1846),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1826),
.B(n_1812),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1846),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1849),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1856),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1839),
.B(n_1817),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1824),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1835),
.B(n_1812),
.Y(n_1901)
);

OAI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1824),
.A2(n_1781),
.B(n_1816),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1849),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1847),
.Y(n_1904)
);

NAND2x1p5_ASAP7_75t_L g1905 ( 
.A(n_1836),
.B(n_1693),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1847),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1845),
.A2(n_1781),
.B(n_1816),
.Y(n_1907)
);

INVxp67_ASAP7_75t_L g1908 ( 
.A(n_1825),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1867),
.B(n_1830),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1880),
.B(n_1830),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1875),
.B(n_1852),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1875),
.B(n_1839),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1859),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1890),
.B(n_1830),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1859),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1893),
.B(n_1847),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1863),
.Y(n_1917)
);

BUFx2_ASAP7_75t_L g1918 ( 
.A(n_1890),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_1877),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1907),
.B(n_1831),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1863),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1893),
.B(n_1848),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1879),
.B(n_1835),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1866),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1866),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1868),
.Y(n_1926)
);

INVx2_ASAP7_75t_SL g1927 ( 
.A(n_1889),
.Y(n_1927)
);

OAI21xp33_ASAP7_75t_L g1928 ( 
.A1(n_1902),
.A2(n_1873),
.B(n_1862),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1879),
.B(n_1844),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1876),
.B(n_1648),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1868),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1869),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1900),
.Y(n_1933)
);

INVx2_ASAP7_75t_SL g1934 ( 
.A(n_1889),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1886),
.B(n_1831),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1892),
.B(n_1831),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1881),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1893),
.B(n_1848),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1882),
.B(n_1832),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1898),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1884),
.B(n_1844),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1895),
.B(n_1850),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1893),
.B(n_1848),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1891),
.B(n_1848),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1900),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_L g1946 ( 
.A1(n_1901),
.A2(n_1813),
.B1(n_1810),
.B2(n_1793),
.Y(n_1946)
);

NAND2x2_ASAP7_75t_L g1947 ( 
.A(n_1891),
.B(n_1825),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1883),
.B(n_1832),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1908),
.B(n_1832),
.Y(n_1949)
);

OAI21xp33_ASAP7_75t_SL g1950 ( 
.A1(n_1920),
.A2(n_1870),
.B(n_1861),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1926),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_L g1952 ( 
.A1(n_1946),
.A2(n_1813),
.B1(n_1793),
.B2(n_1837),
.Y(n_1952)
);

AOI31xp33_ASAP7_75t_L g1953 ( 
.A1(n_1937),
.A2(n_1905),
.A3(n_1871),
.B(n_1870),
.Y(n_1953)
);

INVxp67_ASAP7_75t_L g1954 ( 
.A(n_1918),
.Y(n_1954)
);

AOI32xp33_ASAP7_75t_L g1955 ( 
.A1(n_1918),
.A2(n_1837),
.A3(n_1900),
.B1(n_1793),
.B2(n_1855),
.Y(n_1955)
);

INVxp67_ASAP7_75t_L g1956 ( 
.A(n_1940),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1926),
.Y(n_1957)
);

AOI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1928),
.A2(n_1815),
.B1(n_1813),
.B2(n_1837),
.Y(n_1958)
);

O2A1O1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1914),
.A2(n_1872),
.B(n_1869),
.C(n_1874),
.Y(n_1959)
);

AOI211xp5_ASAP7_75t_SL g1960 ( 
.A1(n_1910),
.A2(n_1836),
.B(n_1841),
.C(n_1861),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1909),
.B(n_1904),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1931),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1931),
.Y(n_1963)
);

OAI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1919),
.A2(n_1815),
.B1(n_1788),
.B2(n_1808),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1932),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1912),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1935),
.A2(n_1813),
.B1(n_1812),
.B2(n_1798),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1936),
.B(n_1923),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1947),
.A2(n_1877),
.B1(n_1814),
.B2(n_1922),
.Y(n_1969)
);

A2O1A1Ixp33_ASAP7_75t_L g1970 ( 
.A1(n_1941),
.A2(n_1794),
.B(n_1798),
.C(n_1788),
.Y(n_1970)
);

NAND3x2_ASAP7_75t_L g1971 ( 
.A(n_1922),
.B(n_1943),
.C(n_1938),
.Y(n_1971)
);

AOI211xp5_ASAP7_75t_L g1972 ( 
.A1(n_1948),
.A2(n_1871),
.B(n_1899),
.C(n_1748),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1932),
.Y(n_1973)
);

INVxp67_ASAP7_75t_L g1974 ( 
.A(n_1930),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1912),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1923),
.B(n_1904),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1913),
.Y(n_1977)
);

O2A1O1Ixp33_ASAP7_75t_L g1978 ( 
.A1(n_1913),
.A2(n_1874),
.B(n_1872),
.C(n_1903),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1916),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1977),
.Y(n_1980)
);

AOI221xp5_ASAP7_75t_L g1981 ( 
.A1(n_1954),
.A2(n_1921),
.B1(n_1924),
.B2(n_1915),
.C(n_1925),
.Y(n_1981)
);

CKINVDCx20_ASAP7_75t_R g1982 ( 
.A(n_1974),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1954),
.A2(n_1917),
.B(n_1915),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1966),
.B(n_1929),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1953),
.B(n_1927),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1951),
.Y(n_1986)
);

OAI322xp33_ASAP7_75t_L g1987 ( 
.A1(n_1958),
.A2(n_1941),
.A3(n_1929),
.B1(n_1939),
.B2(n_1942),
.C1(n_1949),
.C2(n_1934),
.Y(n_1987)
);

NAND4xp25_ASAP7_75t_L g1988 ( 
.A(n_1959),
.B(n_1943),
.C(n_1938),
.D(n_1944),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1971),
.A2(n_1947),
.B1(n_1952),
.B2(n_1969),
.Y(n_1989)
);

AOI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1959),
.A2(n_1934),
.B(n_1927),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1968),
.B(n_1933),
.Y(n_1991)
);

OAI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1967),
.A2(n_1942),
.B1(n_1808),
.B2(n_1945),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1975),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1979),
.B(n_1911),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1956),
.B(n_1933),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1956),
.B(n_1945),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1978),
.A2(n_1921),
.B(n_1917),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1961),
.B(n_1976),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1957),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1962),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1963),
.B(n_1906),
.Y(n_2001)
);

NOR4xp25_ASAP7_75t_L g2002 ( 
.A(n_1978),
.B(n_1925),
.C(n_1924),
.D(n_1944),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1965),
.Y(n_2003)
);

BUFx2_ASAP7_75t_L g2004 ( 
.A(n_1982),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1994),
.B(n_1974),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1997),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_2002),
.B(n_1911),
.Y(n_2007)
);

INVxp67_ASAP7_75t_L g2008 ( 
.A(n_1985),
.Y(n_2008)
);

INVx3_ASAP7_75t_L g2009 ( 
.A(n_1998),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1984),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1995),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1997),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1996),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_2001),
.Y(n_2014)
);

INVx1_ASAP7_75t_SL g2015 ( 
.A(n_1991),
.Y(n_2015)
);

INVx2_ASAP7_75t_SL g2016 ( 
.A(n_1993),
.Y(n_2016)
);

INVxp67_ASAP7_75t_L g2017 ( 
.A(n_1990),
.Y(n_2017)
);

AOI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1987),
.A2(n_1964),
.B1(n_1887),
.B2(n_1864),
.Y(n_2018)
);

O2A1O1Ixp33_ASAP7_75t_L g2019 ( 
.A1(n_1983),
.A2(n_1970),
.B(n_1973),
.C(n_1960),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_2004),
.B(n_1916),
.Y(n_2020)
);

OAI211xp5_ASAP7_75t_L g2021 ( 
.A1(n_2007),
.A2(n_1981),
.B(n_1983),
.C(n_1988),
.Y(n_2021)
);

AOI21xp33_ASAP7_75t_L g2022 ( 
.A1(n_2006),
.A2(n_1986),
.B(n_1980),
.Y(n_2022)
);

INVx2_ASAP7_75t_SL g2023 ( 
.A(n_2004),
.Y(n_2023)
);

NAND3xp33_ASAP7_75t_L g2024 ( 
.A(n_2006),
.B(n_1981),
.C(n_1999),
.Y(n_2024)
);

NAND4xp25_ASAP7_75t_L g2025 ( 
.A(n_2007),
.B(n_1989),
.C(n_1955),
.D(n_2003),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_2009),
.B(n_1992),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_2012),
.B(n_2000),
.Y(n_2027)
);

OAI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_2008),
.A2(n_1972),
.B1(n_1905),
.B2(n_1906),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_2009),
.B(n_1950),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_2009),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2015),
.B(n_1851),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_2016),
.B(n_1851),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_2005),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_SL g2034 ( 
.A(n_2023),
.B(n_2010),
.Y(n_2034)
);

OAI311xp33_ASAP7_75t_L g2035 ( 
.A1(n_2025),
.A2(n_2012),
.A3(n_2019),
.B1(n_2017),
.C1(n_2018),
.Y(n_2035)
);

NOR2xp67_ASAP7_75t_L g2036 ( 
.A(n_2030),
.B(n_2016),
.Y(n_2036)
);

NAND5xp2_ASAP7_75t_L g2037 ( 
.A(n_2021),
.B(n_2014),
.C(n_2013),
.D(n_2011),
.E(n_1829),
.Y(n_2037)
);

AOI222xp33_ASAP7_75t_L g2038 ( 
.A1(n_2024),
.A2(n_1887),
.B1(n_1860),
.B2(n_1864),
.C1(n_1888),
.C2(n_1794),
.Y(n_2038)
);

AOI322xp5_ASAP7_75t_L g2039 ( 
.A1(n_2027),
.A2(n_1887),
.A3(n_1798),
.B1(n_1794),
.B2(n_1860),
.C1(n_1888),
.C2(n_1851),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2020),
.Y(n_2040)
);

OAI211xp5_ASAP7_75t_SL g2041 ( 
.A1(n_2026),
.A2(n_1836),
.B(n_1841),
.C(n_1829),
.Y(n_2041)
);

XNOR2x1_ASAP7_75t_L g2042 ( 
.A(n_2040),
.B(n_2033),
.Y(n_2042)
);

O2A1O1Ixp33_ASAP7_75t_L g2043 ( 
.A1(n_2035),
.A2(n_2027),
.B(n_2029),
.C(n_2022),
.Y(n_2043)
);

OAI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_2036),
.A2(n_2032),
.B1(n_2031),
.B2(n_2028),
.Y(n_2044)
);

AOI221xp5_ASAP7_75t_L g2045 ( 
.A1(n_2037),
.A2(n_1885),
.B1(n_1903),
.B2(n_1878),
.C(n_1897),
.Y(n_2045)
);

AOI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_2034),
.A2(n_1885),
.B(n_1878),
.Y(n_2046)
);

OAI211xp5_ASAP7_75t_L g2047 ( 
.A1(n_2041),
.A2(n_1865),
.B(n_1825),
.C(n_1841),
.Y(n_2047)
);

AOI221xp5_ASAP7_75t_L g2048 ( 
.A1(n_2038),
.A2(n_1897),
.B1(n_1896),
.B2(n_1894),
.C(n_1855),
.Y(n_2048)
);

OAI211xp5_ASAP7_75t_L g2049 ( 
.A1(n_2039),
.A2(n_1865),
.B(n_1825),
.C(n_1836),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_2042),
.B(n_1894),
.Y(n_2050)
);

OAI22xp5_ASAP7_75t_SL g2051 ( 
.A1(n_2044),
.A2(n_2043),
.B1(n_1905),
.B2(n_2047),
.Y(n_2051)
);

NOR2x1_ASAP7_75t_L g2052 ( 
.A(n_2049),
.B(n_1836),
.Y(n_2052)
);

NAND4xp75_ASAP7_75t_L g2053 ( 
.A(n_2046),
.B(n_1899),
.C(n_1842),
.D(n_1682),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2045),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2048),
.B(n_1789),
.Y(n_2055)
);

XNOR2xp5_ASAP7_75t_L g2056 ( 
.A(n_2051),
.B(n_1692),
.Y(n_2056)
);

INVx1_ASAP7_75t_SL g2057 ( 
.A(n_2050),
.Y(n_2057)
);

OAI221xp5_ASAP7_75t_SL g2058 ( 
.A1(n_2054),
.A2(n_1842),
.B1(n_1841),
.B2(n_1814),
.C(n_1896),
.Y(n_2058)
);

NAND4xp75_ASAP7_75t_L g2059 ( 
.A(n_2052),
.B(n_2055),
.C(n_2053),
.D(n_1842),
.Y(n_2059)
);

XNOR2x1_ASAP7_75t_L g2060 ( 
.A(n_2057),
.B(n_1692),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2059),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2060),
.Y(n_2062)
);

AND2x2_ASAP7_75t_SL g2063 ( 
.A(n_2062),
.B(n_2061),
.Y(n_2063)
);

INVx4_ASAP7_75t_L g2064 ( 
.A(n_2062),
.Y(n_2064)
);

AOI22x1_ASAP7_75t_L g2065 ( 
.A1(n_2064),
.A2(n_2056),
.B1(n_2063),
.B2(n_2058),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2063),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_2066),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_2067),
.B(n_2065),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2068),
.Y(n_2069)
);

AOI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_2069),
.A2(n_1858),
.B1(n_1855),
.B2(n_1854),
.Y(n_2070)
);

AOI221xp5_ASAP7_75t_L g2071 ( 
.A1(n_2070),
.A2(n_1688),
.B1(n_1776),
.B2(n_1698),
.C(n_1857),
.Y(n_2071)
);

AOI211xp5_ASAP7_75t_L g2072 ( 
.A1(n_2071),
.A2(n_1730),
.B(n_1694),
.C(n_1841),
.Y(n_2072)
);


endmodule