module fake_jpeg_16641_n_359 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_359);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_359;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_47),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_28),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_29),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_29),
.Y(n_64)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_37),
.B1(n_27),
.B2(n_31),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_37),
.B1(n_49),
.B2(n_27),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_80),
.Y(n_112)
);

NOR2x1_ASAP7_75t_R g105 ( 
.A(n_67),
.B(n_48),
.Y(n_105)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_74),
.Y(n_100)
);

CKINVDCx9p33_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_46),
.B(n_25),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_93),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_96),
.B1(n_102),
.B2(n_110),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_37),
.B1(n_31),
.B2(n_26),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_47),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_31),
.B1(n_49),
.B2(n_83),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_23),
.B(n_25),
.Y(n_136)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_79),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_30),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_69),
.A2(n_26),
.B1(n_49),
.B2(n_24),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_103),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_119),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_117),
.B(n_126),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_142),
.Y(n_147)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_54),
.B1(n_44),
.B2(n_42),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_45),
.Y(n_146)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_130),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_56),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_43),
.B(n_44),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_86),
.B(n_30),
.Y(n_126)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_84),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_139),
.Y(n_158)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_136),
.A2(n_24),
.B1(n_36),
.B2(n_35),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_69),
.B1(n_54),
.B2(n_74),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_137),
.A2(n_141),
.B(n_45),
.C(n_43),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_34),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_97),
.Y(n_140)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_94),
.A2(n_70),
.B1(n_45),
.B2(n_43),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_73),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_56),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_19),
.C(n_18),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_127),
.C(n_125),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_143),
.A2(n_92),
.B(n_107),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_145),
.A2(n_149),
.B(n_153),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_157),
.B1(n_133),
.B2(n_121),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_107),
.B(n_95),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_152),
.B(n_165),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_0),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_155),
.Y(n_176)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_131),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_63),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_166),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_SL g163 ( 
.A(n_122),
.B(n_19),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_141),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_117),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_65),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_71),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_169),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_124),
.A2(n_34),
.B(n_35),
.C(n_28),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_157),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_149),
.A2(n_142),
.B1(n_122),
.B2(n_137),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_171),
.A2(n_173),
.B1(n_184),
.B2(n_190),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_174),
.A2(n_187),
.B(n_194),
.Y(n_205)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_196),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_178),
.B(n_179),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_160),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_180),
.A2(n_193),
.B1(n_164),
.B2(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_121),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_183),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_132),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_100),
.B1(n_140),
.B2(n_127),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_125),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_165),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_129),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_186),
.B(n_188),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_144),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_123),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_146),
.A2(n_153),
.B1(n_147),
.B2(n_163),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_135),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_192),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_150),
.A2(n_120),
.B1(n_164),
.B2(n_114),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_19),
.Y(n_194)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_114),
.B1(n_100),
.B2(n_120),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_148),
.Y(n_201)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_206),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_205),
.A2(n_174),
.B(n_153),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_157),
.B(n_174),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_209),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_148),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_187),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_213),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_183),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_184),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_160),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_211),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_240),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_187),
.Y(n_226)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_177),
.C(n_196),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_244),
.C(n_249),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_195),
.B1(n_190),
.B2(n_189),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_233),
.A2(n_155),
.B1(n_88),
.B2(n_85),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_197),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_150),
.Y(n_236)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_239),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_167),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_214),
.B1(n_215),
.B2(n_223),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_219),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_171),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_205),
.A2(n_215),
.B(n_222),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_245),
.A2(n_223),
.B(n_198),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_203),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_240),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_198),
.B(n_191),
.C(n_167),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_246),
.B1(n_232),
.B2(n_241),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_SL g254 ( 
.A(n_226),
.B(n_212),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_256),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_203),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_236),
.C(n_248),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_263),
.C(n_265),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_264),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_259),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_191),
.C(n_224),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_206),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_146),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_169),
.Y(n_266)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_202),
.Y(n_268)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_242),
.A2(n_157),
.B1(n_200),
.B2(n_152),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_271),
.B1(n_235),
.B2(n_246),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_235),
.A2(n_157),
.B1(n_155),
.B2(n_160),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_44),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_95),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_229),
.C(n_228),
.Y(n_284)
);

INVx11_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_286),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_260),
.A2(n_262),
.B1(n_239),
.B2(n_269),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_278),
.A2(n_279),
.B1(n_285),
.B2(n_277),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_290),
.C(n_251),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_228),
.B1(n_231),
.B2(n_249),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_243),
.Y(n_287)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_17),
.Y(n_288)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_289),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_95),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_263),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_292),
.B(n_273),
.Y(n_301)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_295),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_283),
.A2(n_281),
.B(n_285),
.Y(n_296)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_296),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_257),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_302),
.Y(n_317)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_298),
.A2(n_304),
.B1(n_66),
.B2(n_65),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_305),
.C(n_289),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_276),
.B1(n_290),
.B2(n_282),
.Y(n_310)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_258),
.C(n_251),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_265),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_282),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_0),
.B(n_1),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_89),
.C(n_73),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_274),
.B(n_1),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_R g315 ( 
.A(n_306),
.B(n_1),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_291),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_313),
.C(n_316),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_22),
.C(n_71),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_17),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_320),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_315),
.A2(n_306),
.B1(n_308),
.B2(n_4),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_22),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_294),
.A2(n_36),
.B1(n_22),
.B2(n_50),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_318),
.B(n_320),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_33),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_66),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_317),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_334),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_295),
.C(n_309),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_325),
.B(n_329),
.C(n_321),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_326),
.B(n_331),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_299),
.C(n_296),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_307),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_L g344 ( 
.A1(n_332),
.A2(n_335),
.A3(n_50),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_8),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_304),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_327),
.A2(n_314),
.B(n_333),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_336),
.A2(n_2),
.B(n_8),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_337),
.B(n_2),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_33),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_339),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_328),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_33),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_340),
.B(n_18),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_330),
.A2(n_50),
.B1(n_3),
.B2(n_4),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_9),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_344),
.A2(n_2),
.B1(n_8),
.B2(n_9),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_345),
.B(n_346),
.Y(n_351)
);

NOR3xp33_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_341),
.C(n_11),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_349),
.A2(n_350),
.B(n_343),
.Y(n_352)
);

AOI322xp5_ASAP7_75t_L g354 ( 
.A1(n_352),
.A2(n_353),
.A3(n_348),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_10),
.Y(n_354)
);

AO21x1_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_351),
.B(n_348),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_339),
.B(n_14),
.Y(n_356)
);

AOI21x1_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_12),
.B(n_14),
.Y(n_357)
);

O2A1O1Ixp33_ASAP7_75t_SL g358 ( 
.A1(n_357),
.A2(n_15),
.B(n_18),
.C(n_315),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_15),
.B(n_18),
.Y(n_359)
);


endmodule