module fake_jpeg_8824_n_55 (n_3, n_2, n_1, n_0, n_4, n_5, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx10_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_9),
.Y(n_20)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_17),
.Y(n_19)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_12),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_21),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_24),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_17),
.B1(n_14),
.B2(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_19),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_12),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_31),
.B1(n_14),
.B2(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_32),
.Y(n_34)
);

MAJx2_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_26),
.C(n_17),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_32),
.C(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_34),
.B1(n_39),
.B2(n_33),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_47),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_8),
.B1(n_11),
.B2(n_2),
.Y(n_47)
);

OAI31xp33_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_42),
.A3(n_47),
.B(n_2),
.Y(n_50)
);

AOI322xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.A3(n_0),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_8),
.Y(n_52)
);

MAJx2_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_8),
.C(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_0),
.B(n_3),
.C(n_5),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_8),
.Y(n_55)
);


endmodule