module fake_jpeg_833_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

AOI21xp33_ASAP7_75t_L g27 ( 
.A1(n_1),
.A2(n_0),
.B(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_50),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_52),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_53),
.B(n_55),
.Y(n_130)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_13),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_56),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_57),
.B(n_63),
.Y(n_114)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_60),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_62),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_2),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_82),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_23),
.B(n_2),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_67),
.B(n_73),
.Y(n_142)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_72),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_32),
.B(n_4),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_23),
.B(n_5),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_74),
.B(n_6),
.Y(n_143)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_43),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_43),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_89),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_91),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_29),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_5),
.C(n_6),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_30),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_95),
.Y(n_138)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_93),
.B(n_94),
.Y(n_148)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_96),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_31),
.B1(n_42),
.B2(n_39),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_99),
.A2(n_100),
.B1(n_104),
.B2(n_139),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_27),
.B1(n_42),
.B2(n_39),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_31),
.B1(n_44),
.B2(n_26),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_115),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_60),
.Y(n_115)
);

OAI32xp33_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_44),
.A3(n_40),
.B1(n_36),
.B2(n_34),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_116),
.A2(n_56),
.B(n_62),
.C(n_85),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_54),
.B(n_40),
.C(n_36),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_137),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_51),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_140),
.Y(n_154)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_85),
.A2(n_34),
.B1(n_7),
.B2(n_8),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_48),
.B(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_130),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_76),
.A2(n_11),
.B1(n_66),
.B2(n_61),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_56),
.B(n_81),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_151),
.B(n_152),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_52),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_160),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_128),
.B1(n_113),
.B2(n_101),
.Y(n_197)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_156),
.A2(n_133),
.B(n_171),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_117),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_158),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_52),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_108),
.B(n_11),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_161),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_62),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_72),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_97),
.A2(n_58),
.B(n_147),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_165),
.B(n_188),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_105),
.B(n_114),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_167),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_147),
.A2(n_111),
.B(n_127),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_102),
.B(n_121),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_111),
.B(n_127),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_98),
.B(n_116),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_141),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_172),
.Y(n_195)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_118),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_107),
.B(n_103),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_175),
.Y(n_199)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_99),
.B(n_122),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_179),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_112),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_144),
.Y(n_180)
);

BUFx24_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_107),
.B(n_131),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_185),
.Y(n_211)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_182),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_122),
.B(n_136),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_126),
.B(n_109),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_187),
.Y(n_219)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_139),
.A2(n_137),
.B(n_129),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_134),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_169),
.A2(n_150),
.B1(n_178),
.B2(n_160),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_207),
.B1(n_175),
.B2(n_162),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_197),
.A2(n_198),
.B1(n_180),
.B2(n_166),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_150),
.A2(n_129),
.B1(n_134),
.B2(n_106),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_106),
.B1(n_113),
.B2(n_101),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_156),
.A2(n_128),
.B1(n_133),
.B2(n_155),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_210),
.A2(n_216),
.B1(n_175),
.B2(n_179),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_218),
.C(n_153),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_155),
.A2(n_185),
.B1(n_171),
.B2(n_168),
.Y(n_216)
);

NAND2xp67_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_182),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_193),
.B(n_206),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_221),
.B(n_238),
.Y(n_251)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

NOR3xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_232),
.C(n_236),
.Y(n_250)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_154),
.B(n_149),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_228),
.B(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_205),
.A2(n_163),
.B(n_172),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_152),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_233),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_230),
.A2(n_231),
.B1(n_243),
.B2(n_215),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_195),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_157),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_234),
.A2(n_239),
.B1(n_204),
.B2(n_219),
.Y(n_247)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_192),
.B(n_167),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_165),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_240),
.C(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_204),
.A2(n_200),
.B1(n_211),
.B2(n_199),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_190),
.B(n_196),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_201),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_241),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_205),
.A2(n_210),
.B(n_216),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_200),
.A2(n_189),
.B1(n_176),
.B2(n_177),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_242),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_252),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_222),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_219),
.C(n_215),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_226),
.C(n_228),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_232),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_194),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_240),
.B(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_258),
.B(n_259),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_230),
.B(n_208),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_231),
.B1(n_234),
.B2(n_243),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_263),
.C(n_265),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_273),
.B1(n_275),
.B2(n_249),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_220),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_255),
.A2(n_241),
.B(n_238),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_253),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_251),
.B(n_212),
.Y(n_268)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

A2O1A1O1Ixp25_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_225),
.B(n_223),
.C(n_227),
.D(n_214),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_271),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_261),
.A2(n_235),
.B1(n_187),
.B2(n_162),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_256),
.B1(n_254),
.B2(n_246),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_214),
.B(n_213),
.Y(n_273)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_162),
.B1(n_213),
.B2(n_209),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_282),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_281),
.A2(n_269),
.B1(n_248),
.B2(n_256),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_273),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_258),
.C(n_251),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_265),
.C(n_267),
.Y(n_291)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_252),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_286),
.B1(n_269),
.B2(n_283),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_262),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_291),
.C(n_293),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_280),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_294),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_245),
.C(n_250),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_276),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_295),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_293),
.C(n_280),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_284),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_288),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_289),
.A2(n_283),
.B(n_266),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_302),
.A2(n_247),
.B(n_292),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_292),
.C(n_290),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_307),
.C(n_298),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_310),
.C(n_303),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_281),
.C(n_272),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_312),
.B(n_313),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_248),
.B(n_254),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_260),
.C(n_194),
.Y(n_313)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_173),
.A3(n_184),
.B1(n_191),
.B2(n_209),
.C1(n_260),
.C2(n_303),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_315),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_314),
.Y(n_317)
);


endmodule