module fake_jpeg_15594_n_316 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_24),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_41),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_17),
.B1(n_21),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_32),
.B1(n_37),
.B2(n_36),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_60),
.B(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_18),
.B(n_30),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_32),
.B(n_20),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_51),
.B1(n_42),
.B2(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_21),
.B1(n_17),
.B2(n_15),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_21),
.B1(n_23),
.B2(n_15),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_53),
.Y(n_92)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_31),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_71),
.B(n_82),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_83),
.Y(n_88)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_39),
.B1(n_38),
.B2(n_33),
.Y(n_74)
);

AO22x1_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_50),
.B1(n_43),
.B2(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_28),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_17),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_24),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_89),
.B1(n_98),
.B2(n_80),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_86),
.B(n_92),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_32),
.B1(n_37),
.B2(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_103),
.B1(n_80),
.B2(n_59),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_24),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_34),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_104),
.C(n_107),
.Y(n_127)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_68),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_39),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_35),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_26),
.B(n_19),
.C(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_23),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_124),
.B1(n_125),
.B2(n_137),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_121),
.Y(n_167)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_59),
.B1(n_80),
.B2(n_79),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_74),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_101),
.C(n_105),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_9),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_85),
.A2(n_79),
.B1(n_73),
.B2(n_15),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_8),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_142),
.C(n_165),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_92),
.B(n_101),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_155),
.B(n_170),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_145),
.B(n_22),
.Y(n_172)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_92),
.B1(n_85),
.B2(n_89),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_110),
.B1(n_88),
.B2(n_108),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_87),
.B1(n_51),
.B2(n_74),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_108),
.B1(n_111),
.B2(n_100),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_157),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_23),
.B(n_22),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_100),
.C(n_91),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_109),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_168),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_58),
.B1(n_74),
.B2(n_39),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_120),
.B1(n_58),
.B2(n_132),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_118),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_39),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_169),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_0),
.B(n_1),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_172),
.B(n_189),
.Y(n_206)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_178),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_162),
.A2(n_122),
.B(n_25),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_174),
.A2(n_196),
.B(n_198),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

AOI22x1_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_147),
.B1(n_141),
.B2(n_163),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_201),
.B1(n_170),
.B2(n_168),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_186),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_193),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_195),
.B1(n_197),
.B2(n_193),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_143),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_169),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_190),
.B(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_164),
.Y(n_193)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_128),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_0),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_145),
.B(n_133),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_200),
.B(n_18),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_1),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_199),
.Y(n_202)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_184),
.Y(n_203)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_142),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_212),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_216),
.B1(n_221),
.B2(n_224),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_209),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_140),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_219),
.C(n_220),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_153),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_165),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_201),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_154),
.B1(n_152),
.B2(n_155),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_84),
.B(n_45),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_217),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_45),
.C(n_47),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_72),
.C(n_33),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_58),
.B1(n_84),
.B2(n_38),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_180),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_225),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_38),
.B1(n_33),
.B2(n_3),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_175),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_216),
.A2(n_196),
.B(n_174),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_227),
.A2(n_19),
.B(n_29),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_187),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_242),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_176),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_233),
.C(n_234),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_176),
.C(n_177),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_208),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_198),
.B(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_214),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_238),
.C(n_240),
.Y(n_261)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_175),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_181),
.C(n_178),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_195),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_185),
.Y(n_245)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_247),
.A2(n_16),
.B1(n_7),
.B2(n_8),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_215),
.B1(n_221),
.B2(n_220),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_254),
.B1(n_29),
.B2(n_16),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_207),
.B1(n_211),
.B2(n_204),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_252),
.B1(n_262),
.B2(n_234),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_217),
.B(n_224),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_246),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_260),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_19),
.B1(n_26),
.B2(n_173),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_230),
.B(n_30),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_30),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_238),
.B(n_20),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_239),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_263),
.A2(n_236),
.B1(n_22),
.B2(n_25),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_233),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_264),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_276),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_229),
.C(n_231),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_269),
.C(n_256),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_249),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_229),
.C(n_231),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_270),
.B(n_275),
.Y(n_279)
);

OAI22x1_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_30),
.B1(n_8),
.B2(n_7),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_252),
.B1(n_259),
.B2(n_249),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_282),
.C(n_287),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_255),
.Y(n_280)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_256),
.C(n_258),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_271),
.C(n_276),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_285),
.A2(n_12),
.B1(n_13),
.B2(n_4),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_20),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_277),
.A2(n_11),
.B(n_14),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_4),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_278),
.C(n_292),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_295),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_6),
.B1(n_13),
.B2(n_11),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_299),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_5),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_279),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_301),
.B(n_306),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_299),
.A2(n_282),
.B(n_285),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_305),
.B1(n_293),
.B2(n_291),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_298),
.A2(n_5),
.B(n_6),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_307),
.C(n_302),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_303),
.B(n_308),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_4),
.B(n_2),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_313),
.A2(n_1),
.B(n_2),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_2),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_3),
.B1(n_38),
.B2(n_20),
.Y(n_316)
);


endmodule