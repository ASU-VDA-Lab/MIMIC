module fake_jpeg_12196_n_200 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_200);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_8),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_90),
.Y(n_106)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_62),
.Y(n_97)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_93),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_73),
.B1(n_91),
.B2(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_109),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_53),
.B(n_76),
.C(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_98),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_65),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_55),
.B1(n_64),
.B2(n_83),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_108),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_57),
.B1(n_74),
.B2(n_59),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_65),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_74),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_115),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_86),
.B1(n_85),
.B2(n_56),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_71),
.B1(n_79),
.B2(n_82),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_80),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_127),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_69),
.Y(n_125)
);

OR2x2_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_126),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_63),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_66),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_63),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_130),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_98),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_80),
.Y(n_136)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_143),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_136),
.B(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_78),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_139),
.B(n_141),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_78),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_67),
.B1(n_61),
.B2(n_60),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_146),
.A2(n_147),
.B1(n_6),
.B2(n_7),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_129),
.B1(n_125),
.B2(n_118),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_125),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_9),
.B(n_10),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_157),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_145),
.B1(n_132),
.B2(n_147),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_156),
.B1(n_167),
.B2(n_14),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_151),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_3),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_166),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_162),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_29),
.Y(n_162)
);

AO221x1_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_148),
.B1(n_152),
.B2(n_137),
.C(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_8),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_156),
.B(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_12),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_171),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_136),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_155),
.B1(n_163),
.B2(n_170),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_180),
.B(n_21),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_178),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_162),
.A2(n_15),
.B(n_17),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_18),
.B(n_20),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_22),
.C(n_28),
.Y(n_186)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_186),
.A2(n_188),
.B1(n_178),
.B2(n_175),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_154),
.C(n_35),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_180),
.Y(n_189)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_190),
.B(n_173),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_193),
.A2(n_191),
.B1(n_177),
.B2(n_185),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_194),
.B(n_184),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_189),
.Y(n_196)
);

NOR4xp25_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_34),
.C(n_36),
.D(n_37),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_40),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_42),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_43),
.B(n_46),
.Y(n_200)
);


endmodule