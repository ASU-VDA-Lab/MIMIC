module real_aes_6191_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_756;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g520 ( .A1(n_0), .A2(n_167), .B(n_521), .C(n_524), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_1), .B(n_516), .Y(n_525) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g165 ( .A(n_3), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_4), .B(n_168), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_5), .A2(n_485), .B(n_560), .Y(n_559) );
OAI22xp5_ASAP7_75t_SL g767 ( .A1(n_6), .A2(n_768), .B1(n_771), .B2(n_772), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_6), .Y(n_772) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_7), .A2(n_175), .B(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_8), .A2(n_37), .B1(n_155), .B2(n_203), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_9), .B(n_175), .Y(n_183) );
AND2x6_ASAP7_75t_L g170 ( .A(n_10), .B(n_171), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_11), .A2(n_170), .B(n_490), .C(n_533), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_12), .A2(n_41), .B1(n_769), .B2(n_770), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_12), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_13), .B(n_115), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_13), .B(n_38), .Y(n_465) );
INVx1_ASAP7_75t_L g149 ( .A(n_14), .Y(n_149) );
INVx1_ASAP7_75t_L g146 ( .A(n_15), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_16), .B(n_151), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_17), .B(n_168), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_18), .B(n_142), .Y(n_249) );
AO32x2_ASAP7_75t_L g219 ( .A1(n_19), .A2(n_141), .A3(n_175), .B1(n_194), .B2(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_20), .B(n_155), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_21), .B(n_142), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_22), .A2(n_57), .B1(n_155), .B2(n_203), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g205 ( .A1(n_23), .A2(n_85), .B1(n_151), .B2(n_155), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_24), .B(n_155), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_25), .A2(n_194), .B(n_490), .C(n_508), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_26), .A2(n_194), .B(n_490), .C(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_27), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_28), .B(n_196), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_29), .A2(n_765), .B1(n_766), .B2(n_767), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_29), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_30), .A2(n_485), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_31), .B(n_196), .Y(n_237) );
INVx2_ASAP7_75t_L g153 ( .A(n_32), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_33), .A2(n_488), .B(n_492), .C(n_498), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_34), .B(n_155), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_35), .B(n_196), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_36), .B(n_214), .Y(n_543) );
INVx1_ASAP7_75t_L g115 ( .A(n_38), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_39), .B(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_40), .Y(n_537) );
INVx1_ASAP7_75t_L g770 ( .A(n_41), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_42), .B(n_168), .Y(n_554) );
OAI22xp5_ASAP7_75t_SL g452 ( .A1(n_43), .A2(n_453), .B1(n_456), .B2(n_457), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_43), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_44), .B(n_485), .Y(n_540) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_45), .A2(n_47), .B1(n_454), .B2(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_45), .Y(n_455) );
OAI22xp5_ASAP7_75t_SL g472 ( .A1(n_45), .A2(n_129), .B1(n_130), .B2(n_455), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_46), .A2(n_488), .B(n_498), .C(n_552), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_47), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_48), .B(n_155), .Y(n_178) );
INVx1_ASAP7_75t_L g522 ( .A(n_49), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_50), .A2(n_94), .B1(n_203), .B2(n_204), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_51), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_52), .B(n_155), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_53), .B(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g553 ( .A(n_54), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_55), .B(n_485), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_56), .B(n_163), .Y(n_182) );
AOI22xp33_ASAP7_75t_SL g247 ( .A1(n_58), .A2(n_62), .B1(n_151), .B2(n_155), .Y(n_247) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_59), .A2(n_69), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_59), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_60), .B(n_155), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_61), .B(n_155), .Y(n_211) );
INVx1_ASAP7_75t_L g171 ( .A(n_63), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_64), .B(n_485), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_65), .B(n_516), .Y(n_565) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_66), .A2(n_157), .B(n_163), .C(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_67), .B(n_155), .Y(n_166) );
INVx1_ASAP7_75t_L g145 ( .A(n_68), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_69), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_70), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_71), .B(n_168), .Y(n_496) );
AO32x2_ASAP7_75t_L g200 ( .A1(n_72), .A2(n_175), .A3(n_194), .B1(n_201), .B2(n_206), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_73), .B(n_169), .Y(n_534) );
INVx1_ASAP7_75t_L g190 ( .A(n_74), .Y(n_190) );
INVx1_ASAP7_75t_L g232 ( .A(n_75), .Y(n_232) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_76), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_77), .B(n_495), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_78), .A2(n_490), .B(n_498), .C(n_587), .Y(n_586) );
AOI222xp33_ASAP7_75t_L g470 ( .A1(n_79), .A2(n_471), .B1(n_763), .B2(n_764), .C1(n_773), .C2(n_777), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_80), .B(n_151), .Y(n_233) );
CKINVDCx16_ASAP7_75t_R g561 ( .A(n_81), .Y(n_561) );
INVx1_ASAP7_75t_L g113 ( .A(n_82), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_83), .A2(n_106), .B1(n_116), .B2(n_782), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_84), .B(n_494), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_86), .B(n_203), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_87), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_88), .B(n_151), .Y(n_236) );
INVx2_ASAP7_75t_L g143 ( .A(n_89), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_90), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_91), .B(n_193), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_92), .B(n_151), .Y(n_179) );
INVx2_ASAP7_75t_L g110 ( .A(n_93), .Y(n_110) );
OR2x2_ASAP7_75t_L g462 ( .A(n_93), .B(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g475 ( .A(n_93), .B(n_464), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_95), .A2(n_104), .B1(n_151), .B2(n_152), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_96), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g493 ( .A(n_97), .Y(n_493) );
INVxp67_ASAP7_75t_L g564 ( .A(n_98), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_99), .B(n_151), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_100), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g530 ( .A(n_101), .Y(n_530) );
INVx1_ASAP7_75t_L g588 ( .A(n_102), .Y(n_588) );
AND2x2_ASAP7_75t_L g555 ( .A(n_103), .B(n_196), .Y(n_555) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g783 ( .A(n_107), .Y(n_783) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_114), .Y(n_107) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_110), .C(n_111), .Y(n_108) );
AND2x2_ASAP7_75t_L g464 ( .A(n_109), .B(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g762 ( .A(n_110), .B(n_464), .Y(n_762) );
NOR2x2_ASAP7_75t_L g779 ( .A(n_110), .B(n_463), .Y(n_779) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_469), .Y(n_116) );
BUFx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g781 ( .A(n_120), .Y(n_781) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_459), .B(n_466), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_127), .B1(n_128), .B2(n_458), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_124), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_125), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_130), .B1(n_451), .B2(n_452), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_417), .Y(n_130) );
NOR3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_321), .C(n_405), .Y(n_131) );
NAND4xp25_ASAP7_75t_L g132 ( .A(n_133), .B(n_264), .C(n_286), .D(n_302), .Y(n_132) );
AOI221xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_197), .B1(n_223), .B2(n_242), .C(n_250), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_173), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_136), .B(n_242), .Y(n_276) );
NAND4xp25_ASAP7_75t_L g316 ( .A(n_136), .B(n_304), .C(n_317), .D(n_319), .Y(n_316) );
INVxp67_ASAP7_75t_L g433 ( .A(n_136), .Y(n_433) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g315 ( .A(n_137), .B(n_253), .Y(n_315) );
AND2x2_ASAP7_75t_L g339 ( .A(n_137), .B(n_173), .Y(n_339) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g306 ( .A(n_138), .B(n_241), .Y(n_306) );
AND2x2_ASAP7_75t_L g346 ( .A(n_138), .B(n_327), .Y(n_346) );
AND2x2_ASAP7_75t_L g363 ( .A(n_138), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_138), .B(n_174), .Y(n_387) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g240 ( .A(n_139), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g258 ( .A(n_139), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g270 ( .A(n_139), .B(n_174), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_139), .B(n_184), .Y(n_292) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_147), .B(n_172), .Y(n_139) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_140), .A2(n_185), .B(n_195), .Y(n_184) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_141), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_142), .Y(n_175) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x2_ASAP7_75t_SL g196 ( .A(n_143), .B(n_144), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_161), .B(n_170), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_154), .C(n_157), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_150), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_150), .A2(n_543), .B(n_544), .Y(n_542) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g156 ( .A(n_153), .Y(n_156) );
INVx1_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
INVx3_ASAP7_75t_L g231 ( .A(n_155), .Y(n_231) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_155), .Y(n_590) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g203 ( .A(n_156), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_156), .Y(n_204) );
AND2x6_ASAP7_75t_L g490 ( .A(n_156), .B(n_491), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g587 ( .A1(n_157), .A2(n_588), .B(n_589), .C(n_590), .Y(n_587) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_158), .A2(n_235), .B(n_236), .Y(n_234) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g495 ( .A(n_159), .Y(n_495) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g169 ( .A(n_160), .Y(n_169) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_160), .Y(n_193) );
INVx1_ASAP7_75t_L g214 ( .A(n_160), .Y(n_214) );
AND2x2_ASAP7_75t_L g486 ( .A(n_160), .B(n_164), .Y(n_486) );
INVx1_ASAP7_75t_L g491 ( .A(n_160), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_165), .B(n_166), .C(n_167), .Y(n_161) );
O2A1O1Ixp5_ASAP7_75t_L g189 ( .A1(n_162), .A2(n_190), .B(n_191), .C(n_192), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_162), .A2(n_509), .B(n_510), .Y(n_508) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_167), .A2(n_181), .B(n_182), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_167), .A2(n_193), .B1(n_221), .B2(n_222), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_167), .A2(n_193), .B1(n_246), .B2(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_168), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_168), .A2(n_187), .B(n_188), .Y(n_186) );
O2A1O1Ixp5_ASAP7_75t_SL g230 ( .A1(n_168), .A2(n_231), .B(n_232), .C(n_233), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_168), .B(n_564), .Y(n_563) );
INVx5_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g201 ( .A1(n_169), .A2(n_193), .B1(n_202), .B2(n_205), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g176 ( .A1(n_170), .A2(n_177), .B(n_180), .Y(n_176) );
BUFx3_ASAP7_75t_L g194 ( .A(n_170), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_170), .A2(n_210), .B(n_215), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_170), .A2(n_230), .B(n_234), .Y(n_229) );
AND2x4_ASAP7_75t_L g485 ( .A(n_170), .B(n_486), .Y(n_485) );
INVx4_ASAP7_75t_SL g499 ( .A(n_170), .Y(n_499) );
NAND2x1p5_ASAP7_75t_L g531 ( .A(n_170), .B(n_486), .Y(n_531) );
AND2x2_ASAP7_75t_L g273 ( .A(n_173), .B(n_274), .Y(n_273) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_173), .A2(n_323), .B1(n_326), .B2(n_328), .C(n_332), .Y(n_322) );
AND2x2_ASAP7_75t_L g381 ( .A(n_173), .B(n_346), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_173), .B(n_363), .Y(n_415) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_184), .Y(n_173) );
INVx3_ASAP7_75t_L g241 ( .A(n_174), .Y(n_241) );
AND2x2_ASAP7_75t_L g290 ( .A(n_174), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g344 ( .A(n_174), .B(n_259), .Y(n_344) );
AND2x2_ASAP7_75t_L g402 ( .A(n_174), .B(n_403), .Y(n_402) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_183), .Y(n_174) );
INVx4_ASAP7_75t_L g244 ( .A(n_175), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_175), .A2(n_540), .B(n_541), .Y(n_539) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_175), .Y(n_558) );
AND2x2_ASAP7_75t_L g242 ( .A(n_184), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g259 ( .A(n_184), .Y(n_259) );
INVx1_ASAP7_75t_L g314 ( .A(n_184), .Y(n_314) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_184), .Y(n_320) );
AND2x2_ASAP7_75t_L g365 ( .A(n_184), .B(n_241), .Y(n_365) );
OR2x2_ASAP7_75t_L g404 ( .A(n_184), .B(n_243), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_189), .B(n_194), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_192), .A2(n_216), .B(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx4_ASAP7_75t_L g523 ( .A(n_193), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g263 ( .A(n_194), .B(n_244), .C(n_245), .Y(n_263) );
INVx2_ASAP7_75t_L g206 ( .A(n_196), .Y(n_206) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_196), .A2(n_209), .B(n_218), .Y(n_208) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_196), .A2(n_229), .B(n_237), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_196), .A2(n_484), .B(n_487), .Y(n_483) );
INVx1_ASAP7_75t_L g513 ( .A(n_196), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_196), .A2(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_197), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_207), .Y(n_197) );
AND2x2_ASAP7_75t_L g400 ( .A(n_198), .B(n_397), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_198), .B(n_382), .Y(n_432) );
BUFx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g331 ( .A(n_199), .B(n_255), .Y(n_331) );
AND2x2_ASAP7_75t_L g380 ( .A(n_199), .B(n_226), .Y(n_380) );
INVx1_ASAP7_75t_L g426 ( .A(n_199), .Y(n_426) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_200), .Y(n_239) );
AND2x2_ASAP7_75t_L g281 ( .A(n_200), .B(n_255), .Y(n_281) );
INVx1_ASAP7_75t_L g298 ( .A(n_200), .Y(n_298) );
AND2x2_ASAP7_75t_L g304 ( .A(n_200), .B(n_219), .Y(n_304) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_204), .Y(n_497) );
INVx2_ASAP7_75t_L g524 ( .A(n_204), .Y(n_524) );
INVx1_ASAP7_75t_L g511 ( .A(n_206), .Y(n_511) );
AND2x2_ASAP7_75t_L g372 ( .A(n_207), .B(n_280), .Y(n_372) );
INVx2_ASAP7_75t_L g437 ( .A(n_207), .Y(n_437) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_219), .Y(n_207) );
AND2x2_ASAP7_75t_L g254 ( .A(n_208), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g267 ( .A(n_208), .B(n_227), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_208), .B(n_226), .Y(n_295) );
INVx1_ASAP7_75t_L g301 ( .A(n_208), .Y(n_301) );
INVx1_ASAP7_75t_L g318 ( .A(n_208), .Y(n_318) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_208), .Y(n_330) );
INVx2_ASAP7_75t_L g398 ( .A(n_208), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_210) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g255 ( .A(n_219), .Y(n_255) );
BUFx2_ASAP7_75t_L g352 ( .A(n_219), .Y(n_352) );
AND2x2_ASAP7_75t_L g397 ( .A(n_219), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_238), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_225), .B(n_334), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_225), .A2(n_396), .B(n_410), .Y(n_420) );
AND2x2_ASAP7_75t_L g445 ( .A(n_225), .B(n_331), .Y(n_445) );
BUFx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g367 ( .A(n_227), .Y(n_367) );
AND2x2_ASAP7_75t_L g396 ( .A(n_227), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_228), .Y(n_280) );
INVx2_ASAP7_75t_L g299 ( .A(n_228), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_228), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g253 ( .A(n_239), .Y(n_253) );
OR2x2_ASAP7_75t_L g266 ( .A(n_239), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g334 ( .A(n_239), .B(n_330), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_239), .B(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g435 ( .A(n_239), .B(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_239), .B(n_372), .Y(n_447) );
AND2x2_ASAP7_75t_L g326 ( .A(n_240), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g349 ( .A(n_240), .B(n_242), .Y(n_349) );
INVx2_ASAP7_75t_L g261 ( .A(n_241), .Y(n_261) );
AND2x2_ASAP7_75t_L g289 ( .A(n_241), .B(n_262), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_241), .B(n_314), .Y(n_370) );
AND2x2_ASAP7_75t_L g284 ( .A(n_242), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g431 ( .A(n_242), .Y(n_431) );
AND2x2_ASAP7_75t_L g443 ( .A(n_242), .B(n_306), .Y(n_443) );
AND2x2_ASAP7_75t_L g269 ( .A(n_243), .B(n_259), .Y(n_269) );
INVx1_ASAP7_75t_L g364 ( .A(n_243), .Y(n_364) );
AO21x1_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_248), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_244), .B(n_501), .Y(n_500) );
INVx3_ASAP7_75t_L g516 ( .A(n_244), .Y(n_516) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_244), .A2(n_529), .B(n_536), .Y(n_528) );
AO21x2_ASAP7_75t_L g584 ( .A1(n_244), .A2(n_585), .B(n_592), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_244), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x4_ASAP7_75t_L g262 ( .A(n_249), .B(n_263), .Y(n_262) );
INVxp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_256), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_253), .B(n_300), .Y(n_309) );
OR2x2_ASAP7_75t_L g441 ( .A(n_253), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g358 ( .A(n_254), .B(n_299), .Y(n_358) );
AND2x2_ASAP7_75t_L g366 ( .A(n_254), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g425 ( .A(n_254), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g449 ( .A(n_254), .B(n_296), .Y(n_449) );
NOR2xp67_ASAP7_75t_L g407 ( .A(n_255), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g436 ( .A(n_255), .B(n_299), .Y(n_436) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2x1p5_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
AND2x2_ASAP7_75t_L g288 ( .A(n_258), .B(n_289), .Y(n_288) );
INVxp67_ASAP7_75t_L g450 ( .A(n_258), .Y(n_450) );
NOR2x1_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g285 ( .A(n_261), .Y(n_285) );
AND2x2_ASAP7_75t_L g336 ( .A(n_261), .B(n_269), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_261), .B(n_404), .Y(n_430) );
INVx2_ASAP7_75t_L g275 ( .A(n_262), .Y(n_275) );
INVx3_ASAP7_75t_L g327 ( .A(n_262), .Y(n_327) );
OR2x2_ASAP7_75t_L g355 ( .A(n_262), .B(n_356), .Y(n_355) );
AOI311xp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_268), .A3(n_270), .B(n_271), .C(n_282), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g302 ( .A1(n_265), .A2(n_303), .B(n_305), .C(n_307), .Y(n_302) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_SL g287 ( .A(n_267), .Y(n_287) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g305 ( .A(n_269), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_269), .B(n_285), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_269), .B(n_270), .Y(n_438) );
AND2x2_ASAP7_75t_L g360 ( .A(n_270), .B(n_274), .Y(n_360) );
AOI21xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_276), .B(n_277), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g418 ( .A(n_274), .B(n_306), .Y(n_418) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_275), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g312 ( .A(n_275), .Y(n_312) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
AND2x2_ASAP7_75t_L g303 ( .A(n_279), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g348 ( .A(n_281), .Y(n_348) );
AND2x4_ASAP7_75t_L g410 ( .A(n_281), .B(n_379), .Y(n_410) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AOI222xp33_ASAP7_75t_L g361 ( .A1(n_284), .A2(n_350), .B1(n_362), .B2(n_366), .C1(n_368), .C2(n_372), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B(n_290), .C(n_293), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_287), .B(n_331), .Y(n_354) );
INVx1_ASAP7_75t_L g376 ( .A(n_289), .Y(n_376) );
INVx1_ASAP7_75t_L g310 ( .A(n_291), .Y(n_310) );
OR2x2_ASAP7_75t_L g375 ( .A(n_292), .B(n_376), .Y(n_375) );
OAI21xp33_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_296), .B(n_300), .Y(n_293) );
NAND3xp33_ASAP7_75t_L g311 ( .A(n_294), .B(n_312), .C(n_313), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g409 ( .A1(n_294), .A2(n_331), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_298), .Y(n_351) );
AND2x2_ASAP7_75t_SL g317 ( .A(n_299), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g408 ( .A(n_299), .Y(n_408) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_299), .Y(n_424) );
INVx2_ASAP7_75t_L g382 ( .A(n_300), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_304), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g356 ( .A(n_306), .Y(n_356) );
OAI221xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_310), .B1(n_311), .B2(n_315), .C(n_316), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_310), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g444 ( .A(n_310), .Y(n_444) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g325 ( .A(n_317), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_317), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g383 ( .A(n_317), .B(n_331), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_317), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g416 ( .A(n_317), .B(n_351), .Y(n_416) );
BUFx3_ASAP7_75t_L g379 ( .A(n_318), .Y(n_379) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND5xp2_ASAP7_75t_L g321 ( .A(n_322), .B(n_340), .C(n_361), .D(n_373), .E(n_388), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI32xp33_ASAP7_75t_L g413 ( .A1(n_325), .A2(n_352), .A3(n_368), .B1(n_414), .B2(n_416), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_327), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g337 ( .A(n_331), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B1(n_337), .B2(n_338), .Y(n_332) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_347), .B1(n_349), .B2(n_350), .C(n_353), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g412 ( .A(n_344), .B(n_363), .Y(n_412) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_349), .A2(n_410), .B1(n_428), .B2(n_433), .C(n_434), .Y(n_427) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx2_ASAP7_75t_L g393 ( .A(n_352), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_357), .B2(n_359), .Y(n_353) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx1_ASAP7_75t_L g371 ( .A(n_363), .Y(n_371) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .B1(n_381), .B2(n_382), .C1(n_383), .C2(n_384), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_382), .A2(n_429), .B1(n_431), .B2(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_394), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_399), .B(n_401), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g442 ( .A(n_397), .Y(n_442) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
A2O1A1Ixp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .B(n_411), .C(n_413), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI211xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B(n_421), .C(n_446), .Y(n_417) );
CKINVDCx16_ASAP7_75t_R g422 ( .A(n_418), .Y(n_422) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI211xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B(n_427), .C(n_439), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B(n_438), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_443), .B1(n_444), .B2(n_445), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI21xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B(n_450), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_453), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_462), .Y(n_468) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_466), .B(n_470), .C(n_780), .Y(n_469) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OAI22xp5_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_473), .B1(n_476), .B2(n_762), .Y(n_471) );
INVx1_ASAP7_75t_L g774 ( .A(n_472), .Y(n_774) );
OAI22x1_ASAP7_75t_SL g773 ( .A1(n_473), .A2(n_477), .B1(n_774), .B2(n_775), .Y(n_773) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OR3x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_676), .C(n_719), .Y(n_477) );
NAND5xp2_ASAP7_75t_L g478 ( .A(n_479), .B(n_603), .C(n_633), .D(n_650), .E(n_665), .Y(n_478) );
AOI221xp5_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_526), .B1(n_566), .B2(n_572), .C(n_576), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_502), .Y(n_480) );
OR2x2_ASAP7_75t_L g581 ( .A(n_481), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g620 ( .A(n_481), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g638 ( .A(n_481), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_481), .B(n_574), .Y(n_655) );
OR2x2_ASAP7_75t_L g667 ( .A(n_481), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_481), .B(n_626), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_481), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_481), .B(n_604), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_481), .B(n_612), .Y(n_718) );
AND2x2_ASAP7_75t_L g750 ( .A(n_481), .B(n_514), .Y(n_750) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_481), .Y(n_758) );
INVx5_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_482), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g578 ( .A(n_482), .B(n_556), .Y(n_578) );
BUFx2_ASAP7_75t_L g600 ( .A(n_482), .Y(n_600) );
AND2x2_ASAP7_75t_L g629 ( .A(n_482), .B(n_503), .Y(n_629) );
AND2x2_ASAP7_75t_L g684 ( .A(n_482), .B(n_582), .Y(n_684) );
OR2x6_ASAP7_75t_L g482 ( .A(n_483), .B(n_500), .Y(n_482) );
BUFx2_ASAP7_75t_L g506 ( .A(n_485), .Y(n_506) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_489), .A2(n_499), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g560 ( .A1(n_489), .A2(n_499), .B(n_561), .C(n_562), .Y(n_560) );
INVx5_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B(n_496), .C(n_497), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g552 ( .A1(n_494), .A2(n_497), .B(n_553), .C(n_554), .Y(n_552) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_502), .B(n_638), .Y(n_647) );
OAI32xp33_ASAP7_75t_L g661 ( .A1(n_502), .A2(n_597), .A3(n_662), .B1(n_663), .B2(n_664), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_502), .B(n_663), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_502), .B(n_581), .Y(n_704) );
INVx1_ASAP7_75t_SL g733 ( .A(n_502), .Y(n_733) );
NAND4xp25_ASAP7_75t_L g742 ( .A(n_502), .B(n_528), .C(n_684), .D(n_743), .Y(n_742) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_514), .Y(n_502) );
INVx5_ASAP7_75t_L g575 ( .A(n_503), .Y(n_575) );
AND2x2_ASAP7_75t_L g604 ( .A(n_503), .B(n_515), .Y(n_604) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_503), .Y(n_683) );
AND2x2_ASAP7_75t_L g753 ( .A(n_503), .B(n_700), .Y(n_753) );
OR2x6_ASAP7_75t_L g503 ( .A(n_504), .B(n_512), .Y(n_503) );
AOI21xp5_ASAP7_75t_SL g504 ( .A1(n_505), .A2(n_507), .B(n_511), .Y(n_504) );
AND2x4_ASAP7_75t_L g626 ( .A(n_514), .B(n_575), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_514), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g660 ( .A(n_514), .B(n_582), .Y(n_660) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g574 ( .A(n_515), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g612 ( .A(n_515), .B(n_584), .Y(n_612) );
AND2x2_ASAP7_75t_L g621 ( .A(n_515), .B(n_583), .Y(n_621) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_525), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
AOI222xp33_ASAP7_75t_L g689 ( .A1(n_526), .A2(n_690), .B1(n_692), .B2(n_694), .C1(n_697), .C2(n_698), .Y(n_689) );
AND2x4_ASAP7_75t_L g526 ( .A(n_527), .B(n_545), .Y(n_526) );
AND2x2_ASAP7_75t_L g622 ( .A(n_527), .B(n_623), .Y(n_622) );
NAND3xp33_ASAP7_75t_L g739 ( .A(n_527), .B(n_600), .C(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_538), .Y(n_527) );
INVx5_ASAP7_75t_SL g571 ( .A(n_528), .Y(n_571) );
OAI322xp33_ASAP7_75t_L g576 ( .A1(n_528), .A2(n_577), .A3(n_579), .B1(n_580), .B2(n_594), .C1(n_597), .C2(n_599), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_528), .B(n_569), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_528), .B(n_557), .Y(n_748) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_532), .Y(n_529) );
INVx2_ASAP7_75t_L g569 ( .A(n_538), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_538), .B(n_547), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_545), .B(n_607), .Y(n_662) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g641 ( .A(n_546), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_556), .Y(n_546) );
OR2x2_ASAP7_75t_L g570 ( .A(n_547), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_547), .B(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g609 ( .A(n_547), .B(n_557), .Y(n_609) );
AND2x2_ASAP7_75t_L g632 ( .A(n_547), .B(n_569), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_547), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g648 ( .A(n_547), .B(n_607), .Y(n_648) );
AND2x2_ASAP7_75t_L g656 ( .A(n_547), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_547), .B(n_616), .Y(n_706) );
INVx5_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g596 ( .A(n_548), .B(n_571), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_548), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g623 ( .A(n_548), .B(n_557), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_548), .B(n_670), .Y(n_711) );
OR2x2_ASAP7_75t_L g727 ( .A(n_548), .B(n_671), .Y(n_727) );
AND2x2_ASAP7_75t_SL g734 ( .A(n_548), .B(n_688), .Y(n_734) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_548), .Y(n_741) );
OR2x6_ASAP7_75t_L g548 ( .A(n_549), .B(n_555), .Y(n_548) );
AND2x2_ASAP7_75t_L g595 ( .A(n_556), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g645 ( .A(n_556), .B(n_569), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_556), .B(n_571), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_556), .B(n_607), .Y(n_729) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_557), .B(n_571), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_557), .B(n_569), .Y(n_617) );
OR2x2_ASAP7_75t_L g671 ( .A(n_557), .B(n_569), .Y(n_671) );
AND2x2_ASAP7_75t_L g688 ( .A(n_557), .B(n_568), .Y(n_688) );
INVxp67_ASAP7_75t_L g710 ( .A(n_557), .Y(n_710) );
AND2x2_ASAP7_75t_L g737 ( .A(n_557), .B(n_607), .Y(n_737) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_557), .Y(n_744) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B(n_565), .Y(n_557) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_568), .B(n_618), .Y(n_691) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g607 ( .A(n_569), .B(n_571), .Y(n_607) );
OR2x2_ASAP7_75t_L g674 ( .A(n_569), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g618 ( .A(n_570), .Y(n_618) );
OR2x2_ASAP7_75t_L g679 ( .A(n_570), .B(n_671), .Y(n_679) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g579 ( .A(n_574), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_574), .B(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g580 ( .A(n_575), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_575), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_575), .B(n_582), .Y(n_614) );
INVx2_ASAP7_75t_L g659 ( .A(n_575), .Y(n_659) );
AND2x2_ASAP7_75t_L g672 ( .A(n_575), .B(n_612), .Y(n_672) );
AND2x2_ASAP7_75t_L g697 ( .A(n_575), .B(n_621), .Y(n_697) );
INVx1_ASAP7_75t_L g649 ( .A(n_580), .Y(n_649) );
INVx2_ASAP7_75t_SL g636 ( .A(n_581), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_582), .Y(n_639) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_583), .Y(n_602) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx2_ASAP7_75t_L g700 ( .A(n_584), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_591), .Y(n_585) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g669 ( .A(n_596), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g675 ( .A(n_596), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_596), .A2(n_678), .B1(n_680), .B2(n_685), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_596), .B(n_688), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_597), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g631 ( .A(n_598), .Y(n_631) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
OR2x2_ASAP7_75t_L g613 ( .A(n_600), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_600), .B(n_604), .Y(n_664) );
AND2x2_ASAP7_75t_L g687 ( .A(n_600), .B(n_688), .Y(n_687) );
BUFx2_ASAP7_75t_L g663 ( .A(n_602), .Y(n_663) );
AOI211xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B(n_610), .C(n_624), .Y(n_603) );
INVx1_ASAP7_75t_L g627 ( .A(n_604), .Y(n_627) );
OAI221xp5_ASAP7_75t_SL g735 ( .A1(n_604), .A2(n_736), .B1(n_738), .B2(n_739), .C(n_742), .Y(n_735) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g754 ( .A(n_607), .Y(n_754) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g703 ( .A(n_609), .B(n_642), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .B(n_615), .C(n_619), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
OAI32xp33_ASAP7_75t_L g728 ( .A1(n_617), .A2(n_618), .A3(n_681), .B1(n_718), .B2(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
AND2x2_ASAP7_75t_L g760 ( .A(n_620), .B(n_659), .Y(n_760) );
AND2x2_ASAP7_75t_L g707 ( .A(n_621), .B(n_659), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_621), .B(n_629), .Y(n_725) );
AOI31xp33_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_627), .A3(n_628), .B(n_630), .Y(n_624) );
INVxp67_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_626), .B(n_638), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_626), .B(n_636), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g745 ( .A1(n_626), .A2(n_656), .B1(n_746), .B2(n_749), .C(n_751), .Y(n_745) );
CKINVDCx16_ASAP7_75t_R g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
AND2x2_ASAP7_75t_L g651 ( .A(n_631), .B(n_652), .Y(n_651) );
AOI222xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_640), .B1(n_643), .B2(n_646), .C1(n_648), .C2(n_649), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_635), .B(n_637), .Y(n_634) );
INVx1_ASAP7_75t_L g716 ( .A(n_635), .Y(n_716) );
INVx1_ASAP7_75t_L g738 ( .A(n_638), .Y(n_738) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_641), .A2(n_752), .B1(n_754), .B2(n_755), .Y(n_751) );
INVx1_ASAP7_75t_L g657 ( .A(n_642), .Y(n_657) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B1(n_656), .B2(n_658), .C(n_661), .Y(n_650) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g695 ( .A(n_653), .B(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g747 ( .A(n_653), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g722 ( .A(n_658), .Y(n_722) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx1_ASAP7_75t_L g686 ( .A(n_659), .Y(n_686) );
INVx1_ASAP7_75t_L g668 ( .A(n_660), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_663), .B(n_750), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_669), .B1(n_672), .B2(n_673), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g759 ( .A(n_672), .Y(n_759) );
INVxp33_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_674), .B(n_718), .Y(n_717) );
OAI32xp33_ASAP7_75t_L g708 ( .A1(n_675), .A2(n_709), .A3(n_710), .B1(n_711), .B2(n_712), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g676 ( .A(n_677), .B(n_689), .C(n_701), .D(n_713), .Y(n_676) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
NAND2xp33_ASAP7_75t_SL g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_684), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
CKINVDCx16_ASAP7_75t_R g694 ( .A(n_695), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_698), .A2(n_714), .B1(n_731), .B2(n_734), .C(n_735), .Y(n_730) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g749 ( .A(n_700), .B(n_750), .Y(n_749) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B1(n_705), .B2(n_707), .C(n_708), .Y(n_701) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_710), .B(n_741), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_716), .B(n_717), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND4xp25_ASAP7_75t_L g719 ( .A(n_720), .B(n_730), .C(n_745), .D(n_756), .Y(n_719) );
O2A1O1Ixp33_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_724), .B(n_726), .C(n_728), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVxp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g761 ( .A(n_748), .Y(n_761) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_760), .B(n_761), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g776 ( .A(n_762), .Y(n_776) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
CKINVDCx14_ASAP7_75t_R g771 ( .A(n_768), .Y(n_771) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
endmodule