module fake_jpeg_1450_n_225 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_225);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_4),
.B(n_16),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_63),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_45),
.B(n_44),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_83),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_51),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_94),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_80),
.B1(n_77),
.B2(n_72),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_60),
.B1(n_48),
.B2(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_110),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_74),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_101),
.B(n_104),
.Y(n_119)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_74),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_109),
.B1(n_116),
.B2(n_50),
.Y(n_130)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_47),
.B1(n_72),
.B2(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_58),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_108),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_60),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_56),
.B(n_49),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_52),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_48),
.B1(n_60),
.B2(n_47),
.Y(n_109)
);

OR2x2_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_49),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_88),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_113),
.B(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_61),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_50),
.B1(n_48),
.B2(n_69),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_83),
.B1(n_82),
.B2(n_89),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_122),
.B1(n_123),
.B2(n_135),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_89),
.B1(n_69),
.B2(n_57),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_104),
.A2(n_57),
.B1(n_62),
.B2(n_56),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_128),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_65),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_129),
.B(n_112),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_56),
.B1(n_59),
.B2(n_71),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_71),
.B1(n_64),
.B2(n_3),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_98),
.B1(n_105),
.B2(n_100),
.Y(n_149)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_127),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_110),
.Y(n_138)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_148),
.B1(n_140),
.B2(n_145),
.C(n_159),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_11),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_155),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_97),
.A3(n_98),
.B1(n_115),
.B2(n_105),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_147),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_149),
.A2(n_15),
.B1(n_17),
.B2(n_19),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_1),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_150),
.B(n_154),
.Y(n_179)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_2),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_4),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_6),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_37),
.Y(n_167)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_64),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_161),
.C(n_14),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_118),
.A2(n_43),
.B1(n_42),
.B2(n_41),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_160),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_6),
.B(n_7),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_39),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_135),
.B(n_38),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_162),
.A2(n_166),
.B(n_173),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_153),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_172),
.B1(n_174),
.B2(n_15),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_9),
.B(n_10),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_169),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_181),
.C(n_21),
.Y(n_197)
);

AO22x1_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_153),
.B1(n_141),
.B2(n_145),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_12),
.B(n_13),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_159),
.B1(n_143),
.B2(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_151),
.A2(n_25),
.B(n_33),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_183),
.A2(n_35),
.B(n_20),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_193),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_22),
.C(n_26),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_186),
.C(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_17),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_190),
.B(n_192),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_32),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_194),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_197),
.A2(n_172),
.B(n_177),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_175),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_200),
.C(n_203),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_177),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_205),
.A2(n_186),
.B(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_166),
.C(n_182),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_206),
.A2(n_173),
.B(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_198),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_210),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_212),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_191),
.B(n_196),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_202),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_189),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_174),
.B(n_184),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_202),
.B(n_185),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_219),
.B(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_216),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_221),
.B1(n_179),
.B2(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_222),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_223),
.B(n_163),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_178),
.Y(n_225)
);


endmodule