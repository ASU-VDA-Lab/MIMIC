module fake_ariane_538_n_2005 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2005);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2005;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_279;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_212;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_51),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_56),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_39),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_87),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_74),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_34),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_79),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_124),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_34),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_76),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_167),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_56),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_35),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_89),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_165),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_60),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_25),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_12),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_95),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_111),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_53),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_14),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_160),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_43),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_115),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_2),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_82),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_25),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_163),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_138),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_140),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_51),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_12),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_108),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_6),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_158),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_190),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_137),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_72),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_182),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_59),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_168),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_46),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_128),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_40),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_47),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_69),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_15),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_172),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_11),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_185),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_132),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_57),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_57),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_92),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_184),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_177),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_178),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_150),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_122),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_135),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_153),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_45),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_26),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_129),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_14),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_50),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_105),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_146),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_6),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_29),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_64),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_20),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_94),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_47),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_117),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_164),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_194),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_139),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_45),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_104),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_176),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_161),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_133),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_183),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_52),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_30),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_30),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_27),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_102),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_49),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_20),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_13),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_96),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_151),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_26),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_120),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_54),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_70),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_123),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_78),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_28),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_169),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_155),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_125),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_179),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_131),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_38),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_103),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_126),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_28),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_38),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_154),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_23),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_159),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_54),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_18),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_50),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_109),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_44),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_23),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_85),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_53),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_107),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_86),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_93),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_110),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_11),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_21),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_29),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_27),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_152),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_75),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_99),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_41),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_162),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_0),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_4),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_22),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_44),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_13),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_5),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_31),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_40),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_100),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_143),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_191),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_18),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_41),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_166),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_4),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_61),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_59),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_73),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_170),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_106),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_66),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_142),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_188),
.Y(n_359)
);

BUFx10_ASAP7_75t_L g360 ( 
.A(n_97),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_136),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_81),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_71),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_113),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_46),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_98),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_48),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_112),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_16),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_119),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_10),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_36),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_157),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_88),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_127),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_42),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_193),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_61),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_22),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_60),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_77),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_33),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_186),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_43),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_145),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_36),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_101),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_198),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_270),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_329),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_268),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_292),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_319),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_327),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_329),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_204),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_355),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_329),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_335),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_199),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_199),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_263),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_195),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_267),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_200),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_200),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_197),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_335),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_221),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_221),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_226),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_226),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_201),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_228),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_228),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_233),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_219),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_233),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_234),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_234),
.Y(n_420)
);

BUFx2_ASAP7_75t_SL g421 ( 
.A(n_360),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_220),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_253),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_222),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_267),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_288),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_239),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_239),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_225),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_242),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_311),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_296),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_227),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_296),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_253),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_323),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_349),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_242),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_349),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_244),
.Y(n_440)
);

INVxp33_ASAP7_75t_L g441 ( 
.A(n_232),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_244),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_235),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_241),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_328),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_243),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_247),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_247),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_217),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_249),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_249),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_253),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_256),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_248),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_256),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_261),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_229),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_250),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_229),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_253),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_344),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_261),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_254),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_276),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_196),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_276),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_303),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_253),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_277),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_277),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_282),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_282),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_264),
.Y(n_473)
);

INVxp33_ASAP7_75t_SL g474 ( 
.A(n_272),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_341),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_297),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_353),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_297),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_299),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_307),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_299),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_307),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_400),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_400),
.B(n_215),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_452),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_460),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_468),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_390),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_393),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_480),
.A2(n_330),
.B1(n_379),
.B2(n_245),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_402),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_390),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_423),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_394),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_401),
.B(n_215),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_395),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_423),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_395),
.B(n_306),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_426),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_435),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_396),
.B(n_449),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

AOI22x1_ASAP7_75t_SL g503 ( 
.A1(n_431),
.A2(n_312),
.B1(n_320),
.B2(n_321),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_475),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_421),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_398),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_404),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_475),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_397),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_467),
.B(n_360),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_437),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_388),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_398),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_401),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_405),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_405),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_482),
.A2(n_271),
.B1(n_386),
.B2(n_231),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_406),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_406),
.A2(n_309),
.B(n_306),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_465),
.B(n_399),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_409),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_409),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_410),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_410),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_437),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_411),
.B(n_313),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_411),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_391),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_R g529 ( 
.A(n_403),
.B(n_407),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_412),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_412),
.B(n_309),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_414),
.B(n_291),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_414),
.B(n_326),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_415),
.B(n_291),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_415),
.Y(n_535)
);

NOR2x1_ASAP7_75t_L g536 ( 
.A(n_421),
.B(n_265),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_436),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_416),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_416),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_418),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_418),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_419),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_419),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_420),
.B(n_326),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_408),
.B(n_216),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_420),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_427),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_427),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_428),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_428),
.B(n_347),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_430),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_430),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_438),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_438),
.B(n_298),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_440),
.B(n_313),
.Y(n_555)
);

AND3x2_ASAP7_75t_L g556 ( 
.A(n_439),
.B(n_224),
.C(n_298),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_440),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_442),
.B(n_347),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_442),
.B(n_341),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_447),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_445),
.B(n_275),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_447),
.B(n_354),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_493),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_514),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_514),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_511),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_514),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_514),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_493),
.Y(n_569)
);

BUFx10_ASAP7_75t_L g570 ( 
.A(n_489),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_514),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_514),
.Y(n_572)
);

AND2x2_ASAP7_75t_SL g573 ( 
.A(n_483),
.B(n_354),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_SL g574 ( 
.A(n_529),
.B(n_413),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_493),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_514),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_505),
.B(n_474),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_524),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_R g579 ( 
.A(n_494),
.B(n_389),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_505),
.B(n_485),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_524),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_547),
.B(n_448),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_524),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_524),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_547),
.B(n_448),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_520),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_524),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_524),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_517),
.A2(n_286),
.B1(n_289),
.B2(n_280),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_524),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_547),
.B(n_450),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_500),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_520),
.B(n_450),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_536),
.B(n_432),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_546),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_500),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_500),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_536),
.B(n_434),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_546),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_546),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_545),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_545),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_546),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_546),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_508),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_484),
.B(n_451),
.Y(n_606)
);

NOR2x1p5_ASAP7_75t_L g607 ( 
.A(n_509),
.B(n_392),
.Y(n_607)
);

CKINVDCx6p67_ASAP7_75t_R g608 ( 
.A(n_491),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_546),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_549),
.B(n_417),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_508),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_546),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_508),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_486),
.B(n_451),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_497),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_486),
.B(n_422),
.Y(n_616)
);

NAND2xp33_ASAP7_75t_L g617 ( 
.A(n_516),
.B(n_424),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_549),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_548),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_487),
.B(n_453),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_487),
.B(n_429),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_549),
.B(n_453),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_497),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_483),
.B(n_433),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_548),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_483),
.B(n_443),
.Y(n_626)
);

CKINVDCx6p67_ASAP7_75t_R g627 ( 
.A(n_499),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_497),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_483),
.B(n_444),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_548),
.B(n_455),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_497),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_497),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_497),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_497),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_517),
.A2(n_457),
.B1(n_459),
.B2(n_439),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_548),
.B(n_446),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_516),
.B(n_458),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_523),
.B(n_527),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_502),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_523),
.B(n_463),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_502),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_515),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_527),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_484),
.B(n_455),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_502),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_515),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_515),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_502),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_484),
.B(n_456),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_531),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_530),
.B(n_456),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_L g652 ( 
.A(n_530),
.B(n_473),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_502),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_535),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_502),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_502),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_518),
.Y(n_657)
);

OAI22xp33_ASAP7_75t_L g658 ( 
.A1(n_490),
.A2(n_425),
.B1(n_441),
.B2(n_454),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_518),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_518),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_534),
.A2(n_481),
.B1(n_479),
.B2(n_478),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_521),
.Y(n_662)
);

BUFx10_ASAP7_75t_L g663 ( 
.A(n_556),
.Y(n_663)
);

AO22x2_ASAP7_75t_L g664 ( 
.A1(n_490),
.A2(n_481),
.B1(n_479),
.B2(n_478),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_521),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_521),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_522),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_556),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_522),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_522),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_535),
.B(n_462),
.Y(n_671)
);

AND2x6_ASAP7_75t_L g672 ( 
.A(n_559),
.B(n_539),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_510),
.B(n_462),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_538),
.B(n_464),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_538),
.Y(n_675)
);

INVxp33_ASAP7_75t_L g676 ( 
.A(n_561),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_539),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_539),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_540),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_541),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_540),
.B(n_464),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_534),
.A2(n_338),
.B1(n_365),
.B2(n_367),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_541),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_542),
.B(n_466),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_541),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_542),
.B(n_466),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_551),
.B(n_469),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_543),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_543),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_543),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_511),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_R g692 ( 
.A(n_512),
.B(n_461),
.Y(n_692)
);

AND2x2_ASAP7_75t_SL g693 ( 
.A(n_559),
.B(n_356),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_534),
.B(n_554),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_552),
.Y(n_695)
);

INVxp67_ASAP7_75t_SL g696 ( 
.A(n_531),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_552),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_552),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_557),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_557),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_557),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_551),
.B(n_341),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_534),
.B(n_469),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_553),
.B(n_470),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_553),
.B(n_470),
.Y(n_705)
);

INVx5_ASAP7_75t_L g706 ( 
.A(n_526),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_560),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_504),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_504),
.Y(n_709)
);

BUFx4f_ASAP7_75t_L g710 ( 
.A(n_526),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_519),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_554),
.B(n_471),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_504),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_586),
.B(n_525),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_L g715 ( 
.A(n_577),
.B(n_501),
.Y(n_715)
);

BUFx6f_ASAP7_75t_SL g716 ( 
.A(n_570),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_643),
.Y(n_717)
);

INVxp67_ASAP7_75t_SL g718 ( 
.A(n_711),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_573),
.A2(n_560),
.B1(n_532),
.B2(n_495),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_650),
.B(n_495),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_573),
.B(n_519),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_696),
.B(n_495),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_638),
.A2(n_519),
.B(n_533),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_643),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_573),
.B(n_533),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_643),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_580),
.B(n_532),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_664),
.A2(n_476),
.B1(n_471),
.B2(n_472),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_586),
.B(n_532),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_654),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_593),
.B(n_544),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_566),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_654),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_654),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_SL g735 ( 
.A1(n_589),
.A2(n_477),
.B1(n_537),
.B2(n_528),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_675),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_563),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_693),
.B(n_544),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_703),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_711),
.B(n_550),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_L g741 ( 
.A1(n_589),
.A2(n_562),
.B1(n_558),
.B2(n_550),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_693),
.B(n_558),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_711),
.B(n_619),
.Y(n_743)
);

NOR2x2_ASAP7_75t_L g744 ( 
.A(n_703),
.B(n_712),
.Y(n_744)
);

O2A1O1Ixp5_ASAP7_75t_L g745 ( 
.A1(n_619),
.A2(n_496),
.B(n_513),
.C(n_488),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_619),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_711),
.B(n_619),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_675),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_691),
.B(n_525),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_563),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_703),
.B(n_554),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_675),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_693),
.B(n_562),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_624),
.B(n_554),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_579),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_711),
.B(n_559),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_618),
.B(n_625),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_618),
.B(n_559),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_703),
.B(n_488),
.Y(n_759)
);

OAI22xp33_ASAP7_75t_L g760 ( 
.A1(n_703),
.A2(n_472),
.B1(n_476),
.B2(n_498),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_629),
.B(n_492),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_625),
.B(n_492),
.Y(n_762)
);

INVxp67_ASAP7_75t_SL g763 ( 
.A(n_679),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_601),
.B(n_602),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_679),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_569),
.Y(n_766)
);

BUFx5_ASAP7_75t_L g767 ( 
.A(n_672),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_679),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_707),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_616),
.B(n_506),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_621),
.B(n_506),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_606),
.B(n_513),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_606),
.B(n_498),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_712),
.B(n_507),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_644),
.B(n_507),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_644),
.B(n_526),
.Y(n_776)
);

OAI22xp33_ASAP7_75t_L g777 ( 
.A1(n_712),
.A2(n_245),
.B1(n_317),
.B2(n_196),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_601),
.B(n_602),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_712),
.B(n_206),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_707),
.A2(n_308),
.B1(n_302),
.B2(n_337),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_649),
.B(n_526),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_649),
.B(n_526),
.Y(n_782)
);

OAI22x1_ASAP7_75t_SL g783 ( 
.A1(n_608),
.A2(n_293),
.B1(n_372),
.B2(n_342),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_673),
.B(n_526),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_569),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_686),
.A2(n_210),
.B(n_266),
.C(n_271),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_672),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_674),
.B(n_526),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_570),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_704),
.B(n_526),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_672),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_705),
.B(n_526),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_663),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_594),
.B(n_555),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_642),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_637),
.B(n_640),
.Y(n_796)
);

O2A1O1Ixp5_ASAP7_75t_L g797 ( 
.A1(n_687),
.A2(n_361),
.B(n_356),
.C(n_358),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_594),
.B(n_555),
.Y(n_798)
);

NAND2x1_ASAP7_75t_L g799 ( 
.A(n_672),
.B(n_555),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_712),
.A2(n_555),
.B1(n_375),
.B2(n_361),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_710),
.B(n_358),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_582),
.A2(n_314),
.B1(n_343),
.B2(n_331),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_569),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_570),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_710),
.B(n_375),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_672),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_575),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_594),
.B(n_598),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_594),
.B(n_555),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_575),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_598),
.B(n_555),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_608),
.B(n_627),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_692),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_617),
.A2(n_555),
.B1(n_364),
.B2(n_324),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_598),
.B(n_555),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_664),
.A2(n_635),
.B1(n_672),
.B2(n_694),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_598),
.B(n_555),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_646),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_585),
.B(n_504),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_636),
.B(n_348),
.Y(n_820)
);

INVxp67_ASAP7_75t_SL g821 ( 
.A(n_568),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_591),
.B(n_208),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_575),
.Y(n_823)
);

AND2x6_ASAP7_75t_L g824 ( 
.A(n_646),
.B(n_265),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_622),
.B(n_281),
.Y(n_825)
);

NOR3xp33_ASAP7_75t_L g826 ( 
.A(n_574),
.B(n_210),
.C(n_206),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_710),
.B(n_290),
.Y(n_827)
);

NOR3xp33_ASAP7_75t_L g828 ( 
.A(n_610),
.B(n_214),
.C(n_211),
.Y(n_828)
);

NOR3xp33_ASAP7_75t_L g829 ( 
.A(n_626),
.B(n_214),
.C(n_211),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_647),
.Y(n_830)
);

O2A1O1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_630),
.A2(n_246),
.B(n_386),
.C(n_231),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_690),
.B(n_290),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_647),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_682),
.A2(n_376),
.B1(n_352),
.B2(n_351),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_657),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_657),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_663),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_661),
.B(n_294),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_614),
.B(n_246),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_620),
.B(n_266),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_651),
.B(n_287),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_690),
.B(n_290),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_592),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_659),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_652),
.B(n_357),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_668),
.B(n_378),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_668),
.B(n_382),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_627),
.B(n_287),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_671),
.B(n_316),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_672),
.B(n_341),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_659),
.Y(n_851)
);

NAND2x1p5_ASAP7_75t_L g852 ( 
.A(n_706),
.B(n_274),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_694),
.A2(n_230),
.B1(n_387),
.B2(n_385),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_690),
.B(n_695),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_660),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_660),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_688),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_682),
.B(n_202),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_570),
.B(n_216),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_592),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_694),
.B(n_384),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_681),
.B(n_684),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_592),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_690),
.B(n_695),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_695),
.B(n_316),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_688),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_596),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_664),
.A2(n_318),
.B1(n_369),
.B2(n_340),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_664),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_694),
.A2(n_318),
.B1(n_369),
.B2(n_340),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_694),
.B(n_216),
.Y(n_871)
);

BUFx6f_ASAP7_75t_SL g872 ( 
.A(n_663),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_695),
.B(n_273),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_596),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_697),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_568),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_697),
.B(n_317),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_689),
.A2(n_339),
.B(n_380),
.C(n_371),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_597),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_697),
.B(n_290),
.Y(n_880)
);

OAI22xp33_ASAP7_75t_L g881 ( 
.A1(n_658),
.A2(n_371),
.B1(n_380),
.B2(n_339),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_727),
.B(n_697),
.Y(n_882)
);

NAND2x1p5_ASAP7_75t_L g883 ( 
.A(n_787),
.B(n_706),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_738),
.A2(n_590),
.B1(n_568),
.B2(n_708),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_731),
.B(n_689),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_769),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_795),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_770),
.B(n_698),
.Y(n_888)
);

OAI21xp33_ASAP7_75t_L g889 ( 
.A1(n_845),
.A2(n_700),
.B(n_708),
.Y(n_889)
);

BUFx6f_ASAP7_75t_SL g890 ( 
.A(n_774),
.Y(n_890)
);

OR2x6_ASAP7_75t_L g891 ( 
.A(n_812),
.B(n_607),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_737),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_818),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_771),
.B(n_700),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_SL g895 ( 
.A(n_813),
.B(n_676),
.Y(n_895)
);

NAND2x1p5_ASAP7_75t_L g896 ( 
.A(n_787),
.B(n_706),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_773),
.B(n_666),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_774),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_732),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_859),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_741),
.B(n_666),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_741),
.B(n_666),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_742),
.B(n_699),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_750),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_767),
.B(n_787),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_753),
.B(n_699),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_766),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_785),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_725),
.A2(n_568),
.B1(n_590),
.B2(n_708),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_716),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_716),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_868),
.A2(n_683),
.B1(n_667),
.B2(n_669),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_735),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_720),
.B(n_699),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_830),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_803),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_833),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_787),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_868),
.A2(n_683),
.B1(n_667),
.B2(n_669),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_SL g920 ( 
.A1(n_870),
.A2(n_503),
.B1(n_607),
.B2(n_663),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_SL g921 ( 
.A(n_872),
.B(n_360),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_808),
.B(n_708),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_722),
.B(n_862),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_SL g924 ( 
.A(n_775),
.B(n_503),
.C(n_205),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_791),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_791),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_755),
.B(n_590),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_791),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_791),
.Y(n_929)
);

NAND2x1p5_ASAP7_75t_L g930 ( 
.A(n_806),
.B(n_706),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_714),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_719),
.B(n_701),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_751),
.B(n_701),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_767),
.B(n_590),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_761),
.B(n_701),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_749),
.B(n_273),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_848),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_796),
.B(n_564),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_845),
.B(n_662),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_807),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_754),
.B(n_662),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_751),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_772),
.B(n_665),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_806),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_835),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_836),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_796),
.B(n_564),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_806),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_739),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_725),
.B(n_665),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_806),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_844),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_729),
.B(n_728),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_851),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_855),
.Y(n_955)
);

OR2x6_ASAP7_75t_L g956 ( 
.A(n_739),
.B(n_670),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_728),
.B(n_670),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_767),
.B(n_565),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_763),
.A2(n_612),
.B1(n_565),
.B2(n_567),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_759),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_816),
.A2(n_677),
.B1(n_685),
.B2(n_680),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_767),
.B(n_567),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_810),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_779),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_856),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_759),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_823),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_767),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_793),
.B(n_837),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_857),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_870),
.B(n_677),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_764),
.Y(n_972)
);

INVx5_ASAP7_75t_L g973 ( 
.A(n_746),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_764),
.Y(n_974)
);

INVx5_ASAP7_75t_L g975 ( 
.A(n_746),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_866),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_846),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_760),
.B(n_678),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_778),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_869),
.B(n_678),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_789),
.B(n_680),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_872),
.Y(n_982)
);

OAI22xp33_ASAP7_75t_L g983 ( 
.A1(n_777),
.A2(n_685),
.B1(n_341),
.B2(n_709),
.Y(n_983)
);

AND3x1_ASAP7_75t_L g984 ( 
.A(n_826),
.B(n_713),
.C(n_709),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_799),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_767),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_865),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_843),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_723),
.A2(n_713),
.B(n_609),
.C(n_578),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_760),
.B(n_721),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_778),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_875),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_877),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_R g994 ( 
.A(n_804),
.B(n_631),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_846),
.B(n_571),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_847),
.B(n_273),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_875),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_847),
.B(n_571),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_780),
.B(n_713),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_822),
.B(n_572),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_816),
.B(n_572),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_762),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_871),
.B(n_576),
.Y(n_1003)
);

BUFx12f_ASAP7_75t_L g1004 ( 
.A(n_824),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_860),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_861),
.B(n_605),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_871),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_762),
.Y(n_1008)
);

AO22x1_ASAP7_75t_L g1009 ( 
.A1(n_861),
.A2(n_706),
.B1(n_333),
.B2(n_274),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_776),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_834),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_783),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_721),
.B(n_576),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_873),
.B(n_578),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_781),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_717),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_881),
.A2(n_613),
.B1(n_611),
.B2(n_605),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_881),
.A2(n_613),
.B1(n_611),
.B2(n_333),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_777),
.A2(n_794),
.B1(n_809),
.B2(n_798),
.Y(n_1019)
);

INVx4_ASAP7_75t_L g1020 ( 
.A(n_824),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_873),
.B(n_581),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_715),
.B(n_706),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_724),
.A2(n_581),
.B1(n_584),
.B2(n_587),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_782),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_867),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_SL g1026 ( 
.A1(n_820),
.A2(n_702),
.B1(n_252),
.B2(n_255),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_820),
.B(n_583),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_811),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_R g1029 ( 
.A(n_850),
.B(n_631),
.Y(n_1029)
);

AOI211xp5_ASAP7_75t_L g1030 ( 
.A1(n_858),
.A2(n_583),
.B(n_584),
.C(n_612),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_815),
.B(n_587),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_817),
.B(n_588),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_744),
.Y(n_1033)
);

AND2x2_ASAP7_75t_SL g1034 ( 
.A(n_814),
.B(n_800),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_726),
.A2(n_588),
.B1(n_595),
.B2(n_609),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_874),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_879),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_825),
.B(n_595),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_730),
.B(n_599),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_733),
.B(n_599),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_839),
.B(n_600),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_734),
.B(n_600),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_736),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_748),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_752),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_840),
.B(n_603),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_863),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_864),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_718),
.A2(n_603),
.B(n_604),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_841),
.B(n_604),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_765),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_768),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_852),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_802),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_824),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_819),
.Y(n_1056)
);

NOR3xp33_ASAP7_75t_SL g1057 ( 
.A(n_878),
.B(n_218),
.C(n_383),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_849),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_829),
.A2(n_828),
.B1(n_801),
.B2(n_805),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_838),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_854),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_801),
.A2(n_633),
.B1(n_615),
.B2(n_653),
.Y(n_1062)
);

CKINVDCx8_ASAP7_75t_R g1063 ( 
.A(n_824),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_854),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_758),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_824),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_805),
.A2(n_756),
.B1(n_758),
.B2(n_784),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_821),
.B(n_631),
.Y(n_1068)
);

AND2x6_ASAP7_75t_SL g1069 ( 
.A(n_788),
.B(n_0),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_977),
.B(n_853),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_937),
.B(n_756),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_923),
.A2(n_740),
.B(n_743),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_885),
.A2(n_740),
.B(n_743),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_1007),
.A2(n_831),
.B(n_757),
.C(n_790),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_SL g1075 ( 
.A1(n_1011),
.A2(n_257),
.B1(n_203),
.B2(n_207),
.Y(n_1075)
);

INVxp67_ASAP7_75t_L g1076 ( 
.A(n_899),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_960),
.B(n_757),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_936),
.B(n_786),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_990),
.A2(n_792),
.B(n_745),
.C(n_747),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_925),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_935),
.A2(n_747),
.B(n_876),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_925),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_898),
.B(n_827),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_990),
.A2(n_852),
.B1(n_880),
.B2(n_842),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_888),
.A2(n_842),
.B(n_832),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_894),
.A2(n_1021),
.B(n_1014),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1058),
.B(n_631),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_931),
.A2(n_797),
.B(n_832),
.C(n_656),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_960),
.B(n_623),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_886),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_953),
.B(n_623),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_966),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_996),
.B(n_623),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_890),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_901),
.A2(n_902),
.B1(n_983),
.B2(n_1034),
.Y(n_1095)
);

INVx6_ASAP7_75t_L g1096 ( 
.A(n_933),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_887),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_995),
.A2(n_656),
.B(n_655),
.C(n_628),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_910),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_911),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_949),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_964),
.B(n_628),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_1054),
.B(n_655),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_L g1104 ( 
.A(n_920),
.B(n_656),
.C(n_655),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_893),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1060),
.B(n_615),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_938),
.B(n_632),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_942),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1013),
.A2(n_653),
.B(n_648),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_R g1110 ( 
.A(n_982),
.B(n_209),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1013),
.A2(n_648),
.B(n_645),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_895),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_925),
.B(n_632),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_933),
.B(n_633),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_913),
.B(n_1),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_925),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_938),
.B(n_634),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1011),
.B(n_634),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_995),
.A2(n_645),
.B(n_641),
.C(n_639),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1033),
.B(n_1),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_947),
.B(n_639),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_915),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1027),
.A2(n_641),
.B(n_381),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_947),
.B(n_2),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1056),
.B(n_3),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_983),
.A2(n_301),
.B1(n_374),
.B2(n_373),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1027),
.A2(n_377),
.B(n_370),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_890),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_928),
.B(n_212),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_998),
.B(n_3),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_928),
.B(n_1003),
.Y(n_1131)
);

CKINVDCx8_ASAP7_75t_R g1132 ( 
.A(n_982),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_998),
.B(n_5),
.Y(n_1133)
);

AO22x2_ASAP7_75t_L g1134 ( 
.A1(n_1001),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_933),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_969),
.B(n_7),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_969),
.B(n_8),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1034),
.A2(n_295),
.B1(n_366),
.B2(n_223),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_917),
.A2(n_368),
.B1(n_236),
.B2(n_362),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_R g1140 ( 
.A(n_921),
.B(n_213),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_R g1141 ( 
.A(n_900),
.B(n_1063),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_914),
.A2(n_237),
.B(n_359),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_945),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_946),
.A2(n_238),
.B1(n_350),
.B2(n_346),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_891),
.Y(n_1145)
);

AOI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_1003),
.A2(n_363),
.B(n_290),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_952),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_943),
.A2(n_285),
.B(n_345),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_972),
.B(n_240),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_974),
.B(n_251),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_897),
.A2(n_300),
.B(n_336),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_891),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_954),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_934),
.A2(n_284),
.B(n_334),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_934),
.A2(n_283),
.B(n_259),
.Y(n_1155)
);

OAI21xp33_ASAP7_75t_SL g1156 ( 
.A1(n_922),
.A2(n_9),
.B(n_10),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_979),
.B(n_991),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_955),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_882),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_965),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_969),
.B(n_258),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_928),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1006),
.B(n_17),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_928),
.B(n_305),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_891),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_956),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1059),
.A2(n_922),
.B(n_889),
.C(n_993),
.Y(n_1167)
);

AO22x1_ASAP7_75t_L g1168 ( 
.A1(n_1012),
.A2(n_1022),
.B1(n_981),
.B2(n_980),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_970),
.A2(n_304),
.B1(n_262),
.B2(n_325),
.Y(n_1169)
);

NOR2x1_ASAP7_75t_L g1170 ( 
.A(n_918),
.B(n_363),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_918),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_1057),
.B(n_310),
.C(n_269),
.Y(n_1172)
);

NOR2x1_ASAP7_75t_L g1173 ( 
.A(n_944),
.B(n_363),
.Y(n_1173)
);

OAI22x1_ASAP7_75t_L g1174 ( 
.A1(n_976),
.A2(n_260),
.B1(n_278),
.B2(n_279),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1002),
.A2(n_19),
.B(n_21),
.C(n_24),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1008),
.A2(n_19),
.B(n_24),
.C(n_31),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_978),
.A2(n_322),
.B1(n_315),
.B2(n_363),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_989),
.A2(n_1061),
.B(n_1064),
.C(n_1042),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_987),
.B(n_32),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_980),
.B(n_32),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_980),
.B(n_33),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_989),
.A2(n_35),
.B(n_37),
.C(n_42),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_932),
.A2(n_363),
.B1(n_332),
.B2(n_49),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_981),
.A2(n_332),
.B1(n_48),
.B2(n_52),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_984),
.B(n_332),
.C(n_55),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1018),
.A2(n_332),
.B1(n_55),
.B2(n_58),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_992),
.B(n_37),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1018),
.B(n_58),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1043),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1044),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_992),
.B(n_62),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1045),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_956),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1028),
.B(n_62),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_927),
.B(n_63),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_981),
.A2(n_332),
.B1(n_64),
.B2(n_65),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1042),
.A2(n_63),
.B(n_65),
.C(n_66),
.Y(n_1197)
);

INVx4_ASAP7_75t_L g1198 ( 
.A(n_944),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1051),
.A2(n_67),
.B(n_68),
.C(n_80),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1048),
.B(n_67),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_956),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_950),
.A2(n_1031),
.B(n_1032),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_948),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_892),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1048),
.B(n_68),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_904),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_994),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_903),
.B(n_83),
.Y(n_1208)
);

AOI21xp33_ASAP7_75t_L g1209 ( 
.A1(n_939),
.A2(n_999),
.B(n_957),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_1004),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_948),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_994),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_941),
.A2(n_84),
.B(n_90),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1019),
.A2(n_91),
.B1(n_114),
.B2(n_116),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1019),
.A2(n_118),
.B1(n_121),
.B2(n_130),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_927),
.B(n_134),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1052),
.A2(n_141),
.B(n_148),
.C(n_149),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_904),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_906),
.A2(n_156),
.B1(n_171),
.B2(n_173),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_929),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_884),
.A2(n_187),
.B(n_189),
.C(n_192),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1025),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1010),
.B(n_1015),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_SL g1224 ( 
.A1(n_1035),
.A2(n_1067),
.B(n_1065),
.Y(n_1224)
);

O2A1O1Ixp5_ASAP7_75t_L g1225 ( 
.A1(n_958),
.A2(n_962),
.B(n_959),
.C(n_1050),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_973),
.B(n_975),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_1036),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1022),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1067),
.A2(n_1046),
.B1(n_1041),
.B2(n_1035),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1086),
.A2(n_1068),
.B(n_958),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1095),
.A2(n_1183),
.A3(n_1229),
.B(n_1084),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1109),
.A2(n_1049),
.B(n_962),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1209),
.A2(n_1038),
.B(n_1000),
.Y(n_1233)
);

OR2x2_ASAP7_75t_L g1234 ( 
.A(n_1101),
.B(n_1037),
.Y(n_1234)
);

INVx4_ASAP7_75t_L g1235 ( 
.A(n_1099),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1095),
.B(n_1024),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1090),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1111),
.A2(n_968),
.B(n_905),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1202),
.A2(n_905),
.B(n_973),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1202),
.B(n_971),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1183),
.A2(n_1031),
.A3(n_1032),
.B(n_1023),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1223),
.B(n_1016),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1076),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1070),
.A2(n_1026),
.B(n_1069),
.Y(n_1244)
);

INVxp67_ASAP7_75t_SL g1245 ( 
.A(n_1103),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1118),
.B(n_924),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1107),
.A2(n_1121),
.B(n_1117),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1211),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1167),
.B(n_1016),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1075),
.A2(n_1022),
.B1(n_1030),
.B2(n_951),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1130),
.A2(n_909),
.B(n_1039),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1133),
.A2(n_1039),
.B(n_1040),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_SL g1253 ( 
.A1(n_1126),
.A2(n_1020),
.B(n_1055),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1092),
.Y(n_1254)
);

INVx5_ASAP7_75t_L g1255 ( 
.A(n_1096),
.Y(n_1255)
);

AOI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1084),
.A2(n_1009),
.B(n_1005),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1207),
.B(n_951),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1097),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1195),
.A2(n_1040),
.B(n_926),
.C(n_1055),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_SL g1260 ( 
.A1(n_1224),
.A2(n_1020),
.B(n_929),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1132),
.Y(n_1261)
);

NAND3xp33_ASAP7_75t_SL g1262 ( 
.A(n_1138),
.B(n_1140),
.C(n_1115),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1108),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1073),
.A2(n_968),
.B(n_1062),
.Y(n_1264)
);

AOI211x1_ASAP7_75t_L g1265 ( 
.A1(n_1124),
.A2(n_997),
.B(n_1017),
.C(n_926),
.Y(n_1265)
);

NAND2xp33_ASAP7_75t_L g1266 ( 
.A(n_1126),
.B(n_973),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1112),
.B(n_997),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1212),
.B(n_973),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1071),
.B(n_975),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1229),
.A2(n_1091),
.A3(n_1072),
.B(n_1208),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1211),
.Y(n_1271)
);

NAND3x1_ASAP7_75t_L g1272 ( 
.A(n_1104),
.B(n_1053),
.C(n_1004),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1209),
.B(n_961),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1210),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1178),
.A2(n_1062),
.B(n_967),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1168),
.B(n_961),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1105),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1216),
.A2(n_975),
.B(n_986),
.Y(n_1278)
);

INVxp67_ASAP7_75t_SL g1279 ( 
.A(n_1157),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1079),
.A2(n_940),
.B(n_1005),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_SL g1281 ( 
.A1(n_1125),
.A2(n_1182),
.B(n_1098),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1122),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1081),
.A2(n_963),
.B(n_988),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1211),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1078),
.B(n_1017),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1100),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1131),
.A2(n_975),
.B(n_986),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1188),
.A2(n_1066),
.B(n_1053),
.C(n_919),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1214),
.A2(n_988),
.A3(n_1047),
.B(n_907),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_SL g1290 ( 
.A1(n_1226),
.A2(n_908),
.B(n_916),
.C(n_963),
.Y(n_1290)
);

NAND2x1_ASAP7_75t_L g1291 ( 
.A(n_1220),
.B(n_985),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1214),
.A2(n_908),
.A3(n_916),
.B(n_940),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1143),
.B(n_912),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1225),
.A2(n_919),
.B(n_912),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1210),
.B(n_985),
.Y(n_1295)
);

OA21x2_ASAP7_75t_L g1296 ( 
.A1(n_1146),
.A2(n_1029),
.B(n_1066),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1147),
.B(n_985),
.Y(n_1297)
);

NAND2x1_ASAP7_75t_L g1298 ( 
.A(n_1220),
.B(n_985),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_1193),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1210),
.B(n_883),
.Y(n_1300)
);

CKINVDCx11_ASAP7_75t_R g1301 ( 
.A(n_1128),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1180),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1165),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1186),
.A2(n_1029),
.B1(n_896),
.B2(n_930),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1085),
.A2(n_883),
.B(n_896),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1114),
.B(n_930),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1153),
.B(n_1158),
.Y(n_1307)
);

BUFx2_ASAP7_75t_R g1308 ( 
.A(n_1145),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1160),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1161),
.B(n_1149),
.Y(n_1310)
);

INVx8_ASAP7_75t_L g1311 ( 
.A(n_1210),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1119),
.A2(n_1213),
.B(n_1170),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1110),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1189),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1190),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1192),
.Y(n_1316)
);

AO21x2_ASAP7_75t_L g1317 ( 
.A1(n_1146),
.A2(n_1123),
.B(n_1200),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1228),
.B(n_1093),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1186),
.A2(n_1150),
.B1(n_1215),
.B2(n_1169),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1173),
.A2(n_1221),
.B(n_1113),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_SL g1321 ( 
.A1(n_1125),
.A2(n_1215),
.B(n_1179),
.C(n_1129),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1177),
.A2(n_1206),
.A3(n_1204),
.B(n_1218),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1077),
.A2(n_1088),
.B(n_1162),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1136),
.B(n_1137),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1083),
.B(n_1163),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1222),
.Y(n_1326)
);

BUFx4_ASAP7_75t_SL g1327 ( 
.A(n_1152),
.Y(n_1327)
);

INVxp33_ASAP7_75t_SL g1328 ( 
.A(n_1141),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1074),
.A2(n_1185),
.B(n_1205),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1227),
.B(n_1135),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1219),
.A2(n_1177),
.B(n_1087),
.Y(n_1331)
);

AOI211x1_ASAP7_75t_L g1332 ( 
.A1(n_1194),
.A2(n_1181),
.B(n_1144),
.C(n_1169),
.Y(n_1332)
);

AO31x2_ASAP7_75t_L g1333 ( 
.A1(n_1219),
.A2(n_1174),
.A3(n_1106),
.B(n_1142),
.Y(n_1333)
);

INVx4_ASAP7_75t_L g1334 ( 
.A(n_1198),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1166),
.B(n_1201),
.Y(n_1335)
);

OAI22x1_ASAP7_75t_L g1336 ( 
.A1(n_1184),
.A2(n_1196),
.B1(n_1128),
.B2(n_1120),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1089),
.B(n_1077),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_SL g1338 ( 
.A1(n_1175),
.A2(n_1176),
.B(n_1197),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1096),
.B(n_1171),
.Y(n_1339)
);

AO31x2_ASAP7_75t_L g1340 ( 
.A1(n_1151),
.A2(n_1148),
.A3(n_1191),
.B(n_1187),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1198),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1134),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1096),
.B(n_1144),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1080),
.Y(n_1344)
);

AO32x2_ASAP7_75t_L g1345 ( 
.A1(n_1134),
.A2(n_1139),
.A3(n_1156),
.B1(n_1159),
.B2(n_1199),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1139),
.B(n_1094),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_SL g1347 ( 
.A1(n_1217),
.A2(n_1102),
.B(n_1154),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1127),
.A2(n_1164),
.B(n_1162),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1116),
.A2(n_1134),
.B(n_1114),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1116),
.A2(n_1203),
.B(n_1155),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1089),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1080),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1080),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1082),
.B(n_1172),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1082),
.A2(n_1086),
.B(n_718),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1082),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1090),
.Y(n_1357)
);

INVxp67_ASAP7_75t_SL g1358 ( 
.A(n_1103),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1209),
.A2(n_989),
.B(n_1086),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1100),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1109),
.A2(n_1111),
.B(n_1073),
.Y(n_1361)
);

AO31x2_ASAP7_75t_L g1362 ( 
.A1(n_1086),
.A2(n_1095),
.A3(n_1183),
.B(n_1229),
.Y(n_1362)
);

AOI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1109),
.A2(n_1111),
.B(n_1086),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1109),
.A2(n_1111),
.B(n_1073),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1095),
.B(n_923),
.Y(n_1365)
);

OAI22x1_ASAP7_75t_L g1366 ( 
.A1(n_1070),
.A2(n_589),
.B1(n_913),
.B2(n_1138),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1086),
.A2(n_718),
.B(n_923),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1070),
.B(n_489),
.Y(n_1368)
);

O2A1O1Ixp33_ASAP7_75t_SL g1369 ( 
.A1(n_1130),
.A2(n_1133),
.B(n_1124),
.C(n_923),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1070),
.A2(n_1011),
.B1(n_1054),
.B2(n_494),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1095),
.B(n_923),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1109),
.A2(n_1111),
.B(n_1073),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1086),
.A2(n_718),
.B(n_923),
.Y(n_1373)
);

O2A1O1Ixp5_ASAP7_75t_L g1374 ( 
.A1(n_1130),
.A2(n_990),
.B(n_1133),
.C(n_1195),
.Y(n_1374)
);

NOR2xp67_ASAP7_75t_L g1375 ( 
.A(n_1128),
.B(n_755),
.Y(n_1375)
);

AOI21xp33_ASAP7_75t_L g1376 ( 
.A1(n_1095),
.A2(n_1133),
.B(n_1130),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1095),
.A2(n_1167),
.B(n_990),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1086),
.A2(n_1095),
.A3(n_1183),
.B(n_1229),
.Y(n_1378)
);

O2A1O1Ixp5_ASAP7_75t_L g1379 ( 
.A1(n_1130),
.A2(n_990),
.B(n_1133),
.C(n_1195),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1118),
.B(n_936),
.Y(n_1380)
);

AOI211x1_ASAP7_75t_L g1381 ( 
.A1(n_1124),
.A2(n_741),
.B(n_1133),
.C(n_1130),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1211),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1090),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1118),
.B(n_936),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1103),
.B(n_1007),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1118),
.B(n_936),
.Y(n_1386)
);

OA22x2_ASAP7_75t_L g1387 ( 
.A1(n_1138),
.A2(n_589),
.B1(n_735),
.B2(n_920),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1209),
.A2(n_1146),
.B(n_1086),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1095),
.A2(n_1130),
.B1(n_1133),
.B2(n_1124),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1070),
.B(n_520),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1090),
.Y(n_1391)
);

AOI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1389),
.A2(n_1363),
.B(n_1331),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1263),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1377),
.A2(n_1364),
.B(n_1361),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1319),
.A2(n_1377),
.B(n_1374),
.C(n_1379),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1372),
.A2(n_1232),
.B(n_1312),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1368),
.A2(n_1244),
.B1(n_1370),
.B2(n_1366),
.Y(n_1397)
);

AO31x2_ASAP7_75t_L g1398 ( 
.A1(n_1389),
.A2(n_1247),
.A3(n_1342),
.B(n_1236),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1230),
.A2(n_1283),
.B(n_1264),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_1327),
.Y(n_1400)
);

OR2x6_ASAP7_75t_L g1401 ( 
.A(n_1311),
.B(n_1253),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1238),
.A2(n_1280),
.B(n_1355),
.Y(n_1402)
);

OR2x6_ASAP7_75t_L g1403 ( 
.A(n_1311),
.B(n_1349),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1255),
.B(n_1337),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1313),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1275),
.A2(n_1323),
.B(n_1367),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1373),
.A2(n_1305),
.B(n_1320),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1311),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1387),
.A2(n_1262),
.B1(n_1310),
.B2(n_1285),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1307),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1307),
.Y(n_1411)
);

AOI222xp33_ASAP7_75t_L g1412 ( 
.A1(n_1244),
.A2(n_1390),
.B1(n_1380),
.B2(n_1386),
.C1(n_1384),
.C2(n_1245),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1387),
.A2(n_1376),
.B1(n_1371),
.B2(n_1365),
.Y(n_1413)
);

BUFx12f_ASAP7_75t_L g1414 ( 
.A(n_1286),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1239),
.A2(n_1256),
.B(n_1359),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1376),
.A2(n_1371),
.B1(n_1365),
.B2(n_1358),
.Y(n_1416)
);

AO21x2_ASAP7_75t_L g1417 ( 
.A1(n_1294),
.A2(n_1388),
.B(n_1281),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1359),
.A2(n_1249),
.B(n_1260),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1294),
.A2(n_1388),
.B(n_1329),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1301),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1249),
.A2(n_1278),
.B(n_1350),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1295),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1326),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1254),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1347),
.A2(n_1236),
.B(n_1287),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1252),
.A2(n_1251),
.B(n_1385),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1329),
.A2(n_1348),
.B(n_1240),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1237),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1343),
.B(n_1279),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_SL g1430 ( 
.A1(n_1252),
.A2(n_1251),
.B(n_1354),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1258),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1317),
.A2(n_1273),
.B(n_1276),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_SL g1433 ( 
.A(n_1308),
.B(n_1328),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1325),
.A2(n_1338),
.B1(n_1336),
.B2(n_1242),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1277),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_SL g1436 ( 
.A1(n_1354),
.A2(n_1338),
.B(n_1242),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1240),
.A2(n_1304),
.B(n_1233),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1246),
.B(n_1234),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1325),
.B(n_1243),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1282),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1304),
.A2(n_1233),
.B(n_1297),
.Y(n_1441)
);

CKINVDCx11_ASAP7_75t_R g1442 ( 
.A(n_1261),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1266),
.A2(n_1324),
.B(n_1346),
.C(n_1259),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1337),
.B(n_1269),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1235),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1303),
.B(n_1267),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1297),
.A2(n_1273),
.B(n_1296),
.Y(n_1447)
);

AND2x4_ASAP7_75t_SL g1448 ( 
.A(n_1248),
.B(n_1300),
.Y(n_1448)
);

OA21x2_ASAP7_75t_L g1449 ( 
.A1(n_1288),
.A2(n_1293),
.B(n_1276),
.Y(n_1449)
);

NAND2x1p5_ASAP7_75t_L g1450 ( 
.A(n_1255),
.B(n_1300),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1271),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1296),
.A2(n_1291),
.B(n_1298),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1293),
.A2(n_1272),
.B(n_1318),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1318),
.A2(n_1353),
.B(n_1352),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_SL g1455 ( 
.A1(n_1334),
.A2(n_1341),
.B(n_1274),
.Y(n_1455)
);

AO21x2_ASAP7_75t_L g1456 ( 
.A1(n_1317),
.A2(n_1321),
.B(n_1290),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1271),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1339),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1284),
.Y(n_1459)
);

OAI221xp5_ASAP7_75t_L g1460 ( 
.A1(n_1369),
.A2(n_1302),
.B1(n_1250),
.B2(n_1375),
.C(n_1330),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1381),
.A2(n_1332),
.B1(n_1265),
.B2(n_1334),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1257),
.A2(n_1268),
.B(n_1356),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1309),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1344),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1299),
.A2(n_1351),
.B1(n_1360),
.B2(n_1357),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1314),
.A2(n_1316),
.B(n_1383),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1315),
.B(n_1391),
.Y(n_1467)
);

NAND2x1_ASAP7_75t_L g1468 ( 
.A(n_1274),
.B(n_1344),
.Y(n_1468)
);

BUFx2_ASAP7_75t_R g1469 ( 
.A(n_1335),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1284),
.A2(n_1382),
.B(n_1306),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1289),
.A2(n_1292),
.B(n_1378),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1362),
.A2(n_1378),
.B(n_1255),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1270),
.A2(n_1292),
.B(n_1289),
.Y(n_1473)
);

AO31x2_ASAP7_75t_L g1474 ( 
.A1(n_1231),
.A2(n_1378),
.A3(n_1362),
.B(n_1270),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1299),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1362),
.A2(n_1231),
.B(n_1241),
.Y(n_1476)
);

INVx3_ASAP7_75t_SL g1477 ( 
.A(n_1341),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1322),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1231),
.A2(n_1241),
.B(n_1345),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1241),
.A2(n_1333),
.B(n_1340),
.Y(n_1480)
);

A2O1A1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1345),
.A2(n_1333),
.B(n_1340),
.C(n_1322),
.Y(n_1481)
);

AND2x6_ASAP7_75t_L g1482 ( 
.A(n_1345),
.B(n_1319),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_SL g1483 ( 
.A1(n_1368),
.A2(n_1244),
.B(n_1319),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1377),
.A2(n_1364),
.B(n_1361),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1363),
.A2(n_1364),
.B(n_1361),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1363),
.A2(n_1364),
.B(n_1361),
.Y(n_1486)
);

INVx6_ASAP7_75t_L g1487 ( 
.A(n_1255),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1307),
.Y(n_1488)
);

A2O1A1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1319),
.A2(n_1377),
.B(n_1374),
.C(n_1379),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1313),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1307),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1245),
.B(n_1358),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1319),
.A2(n_1368),
.B1(n_1070),
.B2(n_1358),
.Y(n_1493)
);

INVx5_ASAP7_75t_L g1494 ( 
.A(n_1311),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1380),
.B(n_1384),
.Y(n_1495)
);

CKINVDCx6p67_ASAP7_75t_R g1496 ( 
.A(n_1286),
.Y(n_1496)
);

AO21x1_ASAP7_75t_L g1497 ( 
.A1(n_1389),
.A2(n_1376),
.B(n_1319),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1307),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1319),
.A2(n_1368),
.B1(n_1070),
.B2(n_1358),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1307),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1328),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1342),
.Y(n_1502)
);

O2A1O1Ixp33_ASAP7_75t_SL g1503 ( 
.A1(n_1376),
.A2(n_1389),
.B(n_1371),
.C(n_1365),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1328),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1307),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1307),
.Y(n_1506)
);

INVx8_ASAP7_75t_L g1507 ( 
.A(n_1311),
.Y(n_1507)
);

AO31x2_ASAP7_75t_L g1508 ( 
.A1(n_1389),
.A2(n_1247),
.A3(n_1342),
.B(n_1236),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1307),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1368),
.B(n_1389),
.C(n_1310),
.Y(n_1510)
);

AO32x2_ASAP7_75t_L g1511 ( 
.A1(n_1389),
.A2(n_1183),
.A3(n_1095),
.B1(n_1186),
.B2(n_1229),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1307),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1307),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1368),
.B(n_1389),
.C(n_1310),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1307),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1263),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1376),
.A2(n_1377),
.B(n_1256),
.Y(n_1517)
);

AO21x2_ASAP7_75t_L g1518 ( 
.A1(n_1376),
.A2(n_1377),
.B(n_1256),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1255),
.B(n_1337),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1307),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1245),
.B(n_1358),
.Y(n_1521)
);

BUFx12f_ASAP7_75t_L g1522 ( 
.A(n_1313),
.Y(n_1522)
);

BUFx12f_ASAP7_75t_L g1523 ( 
.A(n_1313),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1255),
.B(n_1337),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1313),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1245),
.B(n_1358),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1380),
.B(n_1384),
.Y(n_1527)
);

OA21x2_ASAP7_75t_L g1528 ( 
.A1(n_1377),
.A2(n_1364),
.B(n_1361),
.Y(n_1528)
);

CKINVDCx14_ASAP7_75t_R g1529 ( 
.A(n_1313),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1328),
.Y(n_1530)
);

NAND2xp33_ASAP7_75t_L g1531 ( 
.A(n_1365),
.B(n_1371),
.Y(n_1531)
);

AOI22x1_ASAP7_75t_L g1532 ( 
.A1(n_1366),
.A2(n_1054),
.B1(n_1134),
.B2(n_789),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1245),
.B(n_1358),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1307),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1342),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1307),
.Y(n_1536)
);

AOI222xp33_ASAP7_75t_L g1537 ( 
.A1(n_1366),
.A2(n_517),
.B1(n_490),
.B2(n_881),
.C1(n_735),
.C2(n_920),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1307),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1439),
.B(n_1429),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1510),
.A2(n_1514),
.B1(n_1483),
.B2(n_1499),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1493),
.A2(n_1397),
.B1(n_1413),
.B2(n_1443),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1479),
.B(n_1482),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1398),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1429),
.B(n_1492),
.Y(n_1544)
);

O2A1O1Ixp5_ASAP7_75t_L g1545 ( 
.A1(n_1497),
.A2(n_1434),
.B(n_1489),
.C(n_1395),
.Y(n_1545)
);

O2A1O1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1443),
.A2(n_1503),
.B(n_1489),
.C(n_1395),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1533),
.B(n_1521),
.Y(n_1547)
);

O2A1O1Ixp5_ASAP7_75t_L g1548 ( 
.A1(n_1434),
.A2(n_1461),
.B(n_1426),
.C(n_1472),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1420),
.Y(n_1549)
);

O2A1O1Ixp33_ASAP7_75t_L g1550 ( 
.A1(n_1503),
.A2(n_1531),
.B(n_1537),
.C(n_1413),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1428),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_SL g1552 ( 
.A1(n_1401),
.A2(n_1460),
.B(n_1403),
.Y(n_1552)
);

INVx4_ASAP7_75t_L g1553 ( 
.A(n_1401),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1424),
.B(n_1495),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1431),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1410),
.B(n_1411),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1438),
.B(n_1527),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1446),
.B(n_1475),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1393),
.B(n_1516),
.Y(n_1559)
);

BUFx12f_ASAP7_75t_L g1560 ( 
.A(n_1442),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1444),
.B(n_1412),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1416),
.A2(n_1409),
.B1(n_1532),
.B2(n_1465),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1444),
.B(n_1451),
.Y(n_1563)
);

OA21x2_ASAP7_75t_L g1564 ( 
.A1(n_1473),
.A2(n_1480),
.B(n_1481),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_R g1565 ( 
.A(n_1529),
.B(n_1433),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1467),
.B(n_1488),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1403),
.B(n_1401),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1491),
.B(n_1498),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1500),
.B(n_1505),
.Y(n_1569)
);

AOI21x1_ASAP7_75t_SL g1570 ( 
.A1(n_1445),
.A2(n_1477),
.B(n_1442),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1435),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1479),
.B(n_1482),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1416),
.A2(n_1409),
.B1(n_1477),
.B2(n_1501),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1506),
.B(n_1509),
.Y(n_1574)
);

O2A1O1Ixp5_ASAP7_75t_L g1575 ( 
.A1(n_1392),
.A2(n_1462),
.B(n_1481),
.C(n_1468),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1479),
.B(n_1482),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1512),
.B(n_1513),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1531),
.A2(n_1425),
.B(n_1417),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1515),
.B(n_1520),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1459),
.B(n_1458),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1440),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1501),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1504),
.A2(n_1530),
.B1(n_1469),
.B2(n_1400),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1463),
.B(n_1534),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1536),
.B(n_1538),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1504),
.A2(n_1530),
.B1(n_1420),
.B2(n_1408),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1466),
.Y(n_1587)
);

OA22x2_ASAP7_75t_L g1588 ( 
.A1(n_1436),
.A2(n_1430),
.B1(n_1453),
.B2(n_1519),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1457),
.B(n_1482),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1482),
.B(n_1423),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1502),
.B(n_1535),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1457),
.B(n_1422),
.Y(n_1592)
);

NAND2xp33_ASAP7_75t_SL g1593 ( 
.A(n_1408),
.B(n_1405),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1496),
.A2(n_1490),
.B1(n_1525),
.B2(n_1405),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1473),
.A2(n_1480),
.B(n_1415),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_SL g1596 ( 
.A1(n_1403),
.A2(n_1450),
.B(n_1524),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1490),
.A2(n_1525),
.B1(n_1494),
.B2(n_1464),
.Y(n_1597)
);

O2A1O1Ixp5_ASAP7_75t_L g1598 ( 
.A1(n_1464),
.A2(n_1519),
.B(n_1524),
.C(n_1404),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1404),
.B(n_1524),
.Y(n_1599)
);

O2A1O1Ixp5_ASAP7_75t_L g1600 ( 
.A1(n_1511),
.A2(n_1535),
.B(n_1502),
.C(n_1398),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1508),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1419),
.A2(n_1517),
.B(n_1518),
.C(n_1455),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1494),
.B(n_1454),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1508),
.B(n_1419),
.Y(n_1604)
);

NOR2xp67_ASAP7_75t_L g1605 ( 
.A(n_1522),
.B(n_1523),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1508),
.B(n_1432),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1453),
.B(n_1432),
.Y(n_1607)
);

AOI21x1_ASAP7_75t_SL g1608 ( 
.A1(n_1414),
.A2(n_1523),
.B(n_1522),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1474),
.B(n_1449),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1454),
.B(n_1452),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1470),
.B(n_1511),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1474),
.B(n_1449),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1474),
.B(n_1448),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1407),
.A2(n_1456),
.B(n_1421),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1507),
.A2(n_1511),
.B1(n_1487),
.B2(n_1414),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1415),
.A2(n_1476),
.B(n_1399),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1470),
.B(n_1511),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1474),
.B(n_1448),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1449),
.B(n_1427),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1507),
.A2(n_1487),
.B1(n_1450),
.B2(n_1528),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1427),
.B(n_1476),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1437),
.B(n_1441),
.Y(n_1622)
);

A2O1A1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1437),
.A2(n_1441),
.B(n_1418),
.C(n_1447),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_SL g1624 ( 
.A1(n_1394),
.A2(n_1528),
.B(n_1484),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1507),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1447),
.B(n_1418),
.Y(n_1626)
);

NOR2xp67_ASAP7_75t_L g1627 ( 
.A(n_1456),
.B(n_1421),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1478),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1471),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1394),
.A2(n_1484),
.B1(n_1528),
.B2(n_1471),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_SL g1631 ( 
.A1(n_1406),
.A2(n_1407),
.B(n_1402),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1399),
.B(n_1402),
.Y(n_1632)
);

NOR2x1_ASAP7_75t_SL g1633 ( 
.A(n_1396),
.B(n_1485),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1485),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1486),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1495),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1479),
.B(n_1482),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1398),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1526),
.B(n_1533),
.Y(n_1639)
);

NOR2xp67_ASAP7_75t_L g1640 ( 
.A(n_1510),
.B(n_1514),
.Y(n_1640)
);

AOI21x1_ASAP7_75t_SL g1641 ( 
.A1(n_1439),
.A2(n_1124),
.B(n_1130),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1473),
.A2(n_1480),
.B(n_1481),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1510),
.A2(n_1514),
.B1(n_1483),
.B2(n_1319),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1510),
.A2(n_1514),
.B1(n_1483),
.B2(n_1319),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1479),
.B(n_1482),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1439),
.B(n_1429),
.Y(n_1646)
);

INVx5_ASAP7_75t_L g1647 ( 
.A(n_1401),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1398),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1428),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_SL g1650 ( 
.A1(n_1443),
.A2(n_1095),
.B(n_1365),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1551),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1639),
.B(n_1547),
.Y(n_1652)
);

AO21x2_ASAP7_75t_L g1653 ( 
.A1(n_1607),
.A2(n_1630),
.B(n_1624),
.Y(n_1653)
);

OA21x2_ASAP7_75t_L g1654 ( 
.A1(n_1614),
.A2(n_1623),
.B(n_1578),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1629),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1582),
.B(n_1549),
.Y(n_1656)
);

OR2x6_ASAP7_75t_L g1657 ( 
.A(n_1596),
.B(n_1552),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1555),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1591),
.B(n_1544),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1571),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1581),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1539),
.B(n_1646),
.Y(n_1662)
);

AO21x2_ASAP7_75t_L g1663 ( 
.A1(n_1624),
.A2(n_1627),
.B(n_1623),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1587),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1610),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1649),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1542),
.B(n_1572),
.Y(n_1667)
);

OA21x2_ASAP7_75t_L g1668 ( 
.A1(n_1548),
.A2(n_1619),
.B(n_1600),
.Y(n_1668)
);

OR2x6_ASAP7_75t_L g1669 ( 
.A(n_1596),
.B(n_1552),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1542),
.B(n_1572),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1602),
.A2(n_1631),
.B(n_1621),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1563),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1576),
.B(n_1637),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1556),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1610),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1546),
.A2(n_1550),
.B(n_1541),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1585),
.B(n_1584),
.Y(n_1677)
);

OR2x6_ASAP7_75t_L g1678 ( 
.A(n_1567),
.B(n_1650),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1576),
.B(n_1637),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1545),
.A2(n_1640),
.B(n_1540),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1645),
.B(n_1611),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1568),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1569),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1579),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1580),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1645),
.B(n_1617),
.Y(n_1686)
);

CKINVDCx16_ASAP7_75t_R g1687 ( 
.A(n_1565),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1574),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1610),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1626),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1577),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1643),
.A2(n_1644),
.B1(n_1650),
.B2(n_1561),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1554),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1543),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1626),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1557),
.B(n_1589),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1616),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1562),
.A2(n_1573),
.B(n_1575),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1543),
.Y(n_1699)
);

AO21x2_ASAP7_75t_L g1700 ( 
.A1(n_1601),
.A2(n_1648),
.B(n_1638),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1566),
.B(n_1638),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1601),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1615),
.A2(n_1553),
.B(n_1620),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1648),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1590),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1606),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1603),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1604),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1636),
.B(n_1609),
.Y(n_1709)
);

INVxp67_ASAP7_75t_SL g1710 ( 
.A(n_1612),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1588),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1588),
.Y(n_1712)
);

OA21x2_ASAP7_75t_L g1713 ( 
.A1(n_1622),
.A2(n_1634),
.B(n_1635),
.Y(n_1713)
);

CKINVDCx16_ASAP7_75t_R g1714 ( 
.A(n_1565),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1559),
.B(n_1558),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1655),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1695),
.B(n_1690),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1692),
.A2(n_1633),
.B(n_1632),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1659),
.B(n_1595),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1713),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1707),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1701),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1659),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1695),
.B(n_1616),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1695),
.B(n_1690),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1692),
.A2(n_1680),
.B1(n_1676),
.B2(n_1698),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1690),
.B(n_1595),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1674),
.B(n_1603),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1709),
.B(n_1595),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1655),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1681),
.B(n_1642),
.Y(n_1731)
);

BUFx2_ASAP7_75t_L g1732 ( 
.A(n_1713),
.Y(n_1732)
);

BUFx2_ASAP7_75t_L g1733 ( 
.A(n_1713),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1681),
.B(n_1642),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1651),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1651),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1709),
.B(n_1564),
.Y(n_1737)
);

OAI221xp5_ASAP7_75t_SL g1738 ( 
.A1(n_1676),
.A2(n_1641),
.B1(n_1592),
.B2(n_1618),
.C(n_1613),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1680),
.A2(n_1583),
.B1(n_1560),
.B2(n_1647),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1658),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1665),
.B(n_1564),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1665),
.B(n_1564),
.Y(n_1742)
);

INVx4_ASAP7_75t_L g1743 ( 
.A(n_1657),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1675),
.B(n_1642),
.Y(n_1744)
);

AOI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1698),
.A2(n_1586),
.B1(n_1598),
.B2(n_1594),
.C(n_1549),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1675),
.B(n_1599),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1652),
.B(n_1628),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1687),
.A2(n_1553),
.B1(n_1647),
.B2(n_1560),
.Y(n_1748)
);

INVxp67_ASAP7_75t_SL g1749 ( 
.A(n_1697),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1689),
.B(n_1599),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1664),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1735),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1726),
.A2(n_1712),
.B(n_1711),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1735),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1726),
.A2(n_1712),
.B1(n_1705),
.B2(n_1684),
.C(n_1674),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_SL g1756 ( 
.A1(n_1720),
.A2(n_1714),
.B1(n_1687),
.B2(n_1653),
.Y(n_1756)
);

OR2x6_ASAP7_75t_L g1757 ( 
.A(n_1748),
.B(n_1657),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1746),
.B(n_1672),
.Y(n_1758)
);

AOI33xp33_ASAP7_75t_L g1759 ( 
.A1(n_1745),
.A2(n_1666),
.A3(n_1661),
.B1(n_1660),
.B2(n_1702),
.B3(n_1704),
.Y(n_1759)
);

AOI211xp5_ASAP7_75t_L g1760 ( 
.A1(n_1745),
.A2(n_1738),
.B(n_1718),
.C(n_1720),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_SL g1761 ( 
.A1(n_1720),
.A2(n_1714),
.B1(n_1653),
.B2(n_1668),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1723),
.B(n_1652),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1738),
.A2(n_1739),
.B1(n_1678),
.B2(n_1718),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1747),
.B(n_1686),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1736),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1728),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1746),
.B(n_1693),
.Y(n_1767)
);

OAI33xp33_ASAP7_75t_L g1768 ( 
.A1(n_1722),
.A2(n_1662),
.A3(n_1682),
.B1(n_1683),
.B2(n_1684),
.B3(n_1688),
.Y(n_1768)
);

AOI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1732),
.A2(n_1705),
.B1(n_1682),
.B2(n_1683),
.C(n_1662),
.Y(n_1769)
);

AOI222xp33_ASAP7_75t_L g1770 ( 
.A1(n_1732),
.A2(n_1710),
.B1(n_1708),
.B2(n_1706),
.C1(n_1670),
.C2(n_1667),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1732),
.A2(n_1708),
.B1(n_1688),
.B2(n_1691),
.C(n_1653),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1733),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1746),
.B(n_1696),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1747),
.B(n_1686),
.Y(n_1774)
);

AOI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1733),
.A2(n_1691),
.B1(n_1653),
.B2(n_1706),
.C(n_1661),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1728),
.B(n_1677),
.Y(n_1776)
);

OAI211xp5_ASAP7_75t_L g1777 ( 
.A1(n_1749),
.A2(n_1668),
.B(n_1654),
.C(n_1703),
.Y(n_1777)
);

INVxp67_ASAP7_75t_L g1778 ( 
.A(n_1719),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1750),
.B(n_1678),
.Y(n_1779)
);

AOI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1731),
.A2(n_1660),
.B1(n_1666),
.B2(n_1685),
.C(n_1677),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1747),
.B(n_1673),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1750),
.B(n_1707),
.Y(n_1782)
);

OAI221xp5_ASAP7_75t_L g1783 ( 
.A1(n_1737),
.A2(n_1703),
.B1(n_1679),
.B2(n_1673),
.C(n_1668),
.Y(n_1783)
);

BUFx3_ASAP7_75t_L g1784 ( 
.A(n_1721),
.Y(n_1784)
);

AO21x2_ASAP7_75t_L g1785 ( 
.A1(n_1716),
.A2(n_1730),
.B(n_1751),
.Y(n_1785)
);

OAI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1741),
.A2(n_1671),
.B(n_1668),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1736),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1740),
.Y(n_1788)
);

AOI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1731),
.A2(n_1699),
.B1(n_1694),
.B2(n_1704),
.C(n_1702),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1731),
.A2(n_1669),
.B1(n_1668),
.B2(n_1700),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1734),
.B(n_1715),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1748),
.A2(n_1663),
.B(n_1593),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1740),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1752),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1754),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1765),
.Y(n_1796)
);

INVxp67_ASAP7_75t_L g1797 ( 
.A(n_1783),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1791),
.B(n_1719),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1779),
.B(n_1750),
.Y(n_1799)
);

INVx3_ASAP7_75t_L g1800 ( 
.A(n_1782),
.Y(n_1800)
);

NOR3xp33_ASAP7_75t_SL g1801 ( 
.A(n_1777),
.B(n_1597),
.C(n_1625),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1787),
.Y(n_1802)
);

INVx4_ASAP7_75t_SL g1803 ( 
.A(n_1757),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1756),
.B(n_1750),
.Y(n_1804)
);

INVx4_ASAP7_75t_L g1805 ( 
.A(n_1757),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1769),
.B(n_1719),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1788),
.Y(n_1807)
);

NOR2x1p5_ASAP7_75t_L g1808 ( 
.A(n_1784),
.B(n_1743),
.Y(n_1808)
);

BUFx3_ASAP7_75t_L g1809 ( 
.A(n_1784),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1766),
.B(n_1734),
.Y(n_1810)
);

INVxp67_ASAP7_75t_SL g1811 ( 
.A(n_1760),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1793),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1766),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1756),
.B(n_1750),
.Y(n_1814)
);

OA21x2_ASAP7_75t_L g1815 ( 
.A1(n_1786),
.A2(n_1749),
.B(n_1724),
.Y(n_1815)
);

OA21x2_ASAP7_75t_L g1816 ( 
.A1(n_1775),
.A2(n_1724),
.B(n_1671),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1785),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1762),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1764),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1772),
.Y(n_1820)
);

OA21x2_ASAP7_75t_L g1821 ( 
.A1(n_1790),
.A2(n_1724),
.B(n_1671),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1774),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1759),
.B(n_1734),
.Y(n_1823)
);

OA21x2_ASAP7_75t_L g1824 ( 
.A1(n_1790),
.A2(n_1744),
.B(n_1727),
.Y(n_1824)
);

NAND3xp33_ASAP7_75t_SL g1825 ( 
.A(n_1761),
.B(n_1742),
.C(n_1656),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1813),
.Y(n_1826)
);

AND2x4_ASAP7_75t_SL g1827 ( 
.A(n_1805),
.B(n_1782),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1800),
.B(n_1773),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1794),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1800),
.B(n_1758),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1800),
.B(n_1767),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1794),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1823),
.B(n_1776),
.Y(n_1833)
);

NAND2x1_ASAP7_75t_L g1834 ( 
.A(n_1815),
.B(n_1717),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1795),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1795),
.Y(n_1836)
);

NOR2xp67_ASAP7_75t_L g1837 ( 
.A(n_1825),
.B(n_1792),
.Y(n_1837)
);

INVx3_ASAP7_75t_SL g1838 ( 
.A(n_1809),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1811),
.B(n_1809),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1824),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1818),
.B(n_1759),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1809),
.B(n_1761),
.Y(n_1842)
);

INVx1_ASAP7_75t_SL g1843 ( 
.A(n_1822),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1796),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1796),
.Y(n_1845)
);

NOR2x1_ASAP7_75t_L g1846 ( 
.A(n_1825),
.B(n_1605),
.Y(n_1846)
);

INVx3_ASAP7_75t_L g1847 ( 
.A(n_1815),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1823),
.B(n_1729),
.Y(n_1848)
);

AND2x4_ASAP7_75t_L g1849 ( 
.A(n_1808),
.B(n_1803),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1802),
.Y(n_1850)
);

INVxp67_ASAP7_75t_L g1851 ( 
.A(n_1797),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1803),
.B(n_1778),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1819),
.B(n_1781),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1806),
.B(n_1778),
.Y(n_1854)
);

INVxp67_ASAP7_75t_SL g1855 ( 
.A(n_1797),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1806),
.B(n_1737),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1815),
.B(n_1725),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1802),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1824),
.Y(n_1859)
);

INVx1_ASAP7_75t_SL g1860 ( 
.A(n_1803),
.Y(n_1860)
);

BUFx2_ASAP7_75t_L g1861 ( 
.A(n_1815),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1807),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1849),
.B(n_1803),
.Y(n_1863)
);

NOR2x2_ASAP7_75t_L g1864 ( 
.A(n_1840),
.B(n_1820),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1833),
.B(n_1810),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1828),
.B(n_1799),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1835),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1861),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1828),
.B(n_1799),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1845),
.Y(n_1870)
);

OR4x1_ASAP7_75t_L g1871 ( 
.A(n_1834),
.B(n_1812),
.C(n_1807),
.D(n_1817),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1861),
.Y(n_1872)
);

AND2x2_ASAP7_75t_SL g1873 ( 
.A(n_1839),
.B(n_1824),
.Y(n_1873)
);

INVx3_ASAP7_75t_L g1874 ( 
.A(n_1847),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1829),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1833),
.B(n_1810),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1829),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1855),
.B(n_1812),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_1838),
.Y(n_1879)
);

NOR2x1_ASAP7_75t_R g1880 ( 
.A(n_1849),
.B(n_1625),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1853),
.B(n_1798),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1832),
.Y(n_1882)
);

NOR2x1_ASAP7_75t_L g1883 ( 
.A(n_1846),
.B(n_1804),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1838),
.B(n_1768),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1851),
.B(n_1789),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1827),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1832),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1840),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1826),
.B(n_1780),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1843),
.B(n_1770),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1841),
.B(n_1755),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1837),
.B(n_1771),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1838),
.B(n_1799),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1836),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1846),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1853),
.B(n_1798),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1837),
.B(n_1824),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1854),
.B(n_1820),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1840),
.A2(n_1816),
.B1(n_1821),
.B2(n_1753),
.Y(n_1899)
);

CKINVDCx16_ASAP7_75t_R g1900 ( 
.A(n_1863),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1875),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1866),
.B(n_1831),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1875),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1873),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1885),
.B(n_1842),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1881),
.B(n_1854),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1864),
.Y(n_1907)
);

AND3x1_ASAP7_75t_L g1908 ( 
.A(n_1883),
.B(n_1842),
.C(n_1801),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1868),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_1863),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1888),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1864),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1871),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1866),
.B(n_1831),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1881),
.B(n_1856),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1869),
.B(n_1830),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1896),
.B(n_1856),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1888),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1877),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1882),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1887),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1894),
.Y(n_1922)
);

CKINVDCx16_ASAP7_75t_R g1923 ( 
.A(n_1863),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1879),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1868),
.Y(n_1925)
);

OAI21xp33_ASAP7_75t_L g1926 ( 
.A1(n_1873),
.A2(n_1847),
.B(n_1859),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1900),
.B(n_1886),
.Y(n_1927)
);

OAI22xp5_ASAP7_75t_SL g1928 ( 
.A1(n_1908),
.A2(n_1871),
.B1(n_1895),
.B2(n_1890),
.Y(n_1928)
);

AOI21xp33_ASAP7_75t_L g1929 ( 
.A1(n_1913),
.A2(n_1892),
.B(n_1891),
.Y(n_1929)
);

NOR4xp25_ASAP7_75t_SL g1930 ( 
.A(n_1926),
.B(n_1867),
.C(n_1870),
.D(n_1814),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1900),
.A2(n_1897),
.B1(n_1889),
.B2(n_1899),
.Y(n_1931)
);

INVx2_ASAP7_75t_SL g1932 ( 
.A(n_1923),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1905),
.A2(n_1859),
.B1(n_1884),
.B2(n_1816),
.Y(n_1933)
);

OAI322xp33_ASAP7_75t_L g1934 ( 
.A1(n_1913),
.A2(n_1872),
.A3(n_1878),
.B1(n_1847),
.B2(n_1898),
.C1(n_1834),
.C2(n_1865),
.Y(n_1934)
);

OAI22xp33_ASAP7_75t_L g1935 ( 
.A1(n_1907),
.A2(n_1847),
.B1(n_1816),
.B2(n_1848),
.Y(n_1935)
);

OAI21xp5_ASAP7_75t_SL g1936 ( 
.A1(n_1904),
.A2(n_1893),
.B(n_1886),
.Y(n_1936)
);

OAI211xp5_ASAP7_75t_L g1937 ( 
.A1(n_1904),
.A2(n_1872),
.B(n_1874),
.C(n_1893),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1904),
.A2(n_1874),
.B(n_1898),
.Y(n_1938)
);

OAI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1923),
.A2(n_1896),
.B1(n_1827),
.B2(n_1849),
.Y(n_1939)
);

OAI221xp5_ASAP7_75t_L g1940 ( 
.A1(n_1926),
.A2(n_1816),
.B1(n_1860),
.B2(n_1848),
.C(n_1821),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1909),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1906),
.B(n_1869),
.Y(n_1942)
);

AOI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1907),
.A2(n_1912),
.B1(n_1918),
.B2(n_1911),
.Y(n_1943)
);

NAND3xp33_ASAP7_75t_L g1944 ( 
.A(n_1912),
.B(n_1874),
.C(n_1821),
.Y(n_1944)
);

NAND2xp33_ASAP7_75t_SL g1945 ( 
.A(n_1906),
.B(n_1865),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1902),
.B(n_1830),
.Y(n_1946)
);

OAI221xp5_ASAP7_75t_L g1947 ( 
.A1(n_1915),
.A2(n_1821),
.B1(n_1876),
.B2(n_1805),
.C(n_1763),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1946),
.B(n_1924),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1941),
.Y(n_1949)
);

INVx1_ASAP7_75t_SL g1950 ( 
.A(n_1945),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1942),
.B(n_1910),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1932),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1929),
.B(n_1902),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1927),
.B(n_1914),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1930),
.B(n_1914),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1928),
.Y(n_1956)
);

NOR2x1_ASAP7_75t_L g1957 ( 
.A(n_1936),
.B(n_1925),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1931),
.B(n_1916),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1939),
.B(n_1916),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1943),
.B(n_1915),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1950),
.B(n_1925),
.Y(n_1961)
);

AOI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1960),
.A2(n_1934),
.B(n_1938),
.Y(n_1962)
);

OAI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1955),
.A2(n_1957),
.B(n_1956),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1952),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1948),
.Y(n_1965)
);

AOI21xp33_ASAP7_75t_L g1966 ( 
.A1(n_1953),
.A2(n_1938),
.B(n_1937),
.Y(n_1966)
);

AOI221xp5_ASAP7_75t_L g1967 ( 
.A1(n_1955),
.A2(n_1935),
.B1(n_1940),
.B2(n_1944),
.C(n_1933),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_SL g1968 ( 
.A1(n_1958),
.A2(n_1880),
.B(n_1849),
.Y(n_1968)
);

INVxp67_ASAP7_75t_L g1969 ( 
.A(n_1954),
.Y(n_1969)
);

NAND4xp25_ASAP7_75t_SL g1970 ( 
.A(n_1951),
.B(n_1947),
.C(n_1917),
.D(n_1922),
.Y(n_1970)
);

AOI221xp5_ASAP7_75t_L g1971 ( 
.A1(n_1949),
.A2(n_1911),
.B1(n_1918),
.B2(n_1922),
.C(n_1921),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1969),
.Y(n_1972)
);

NAND5xp2_ASAP7_75t_L g1973 ( 
.A(n_1967),
.B(n_1954),
.C(n_1959),
.D(n_1903),
.E(n_1901),
.Y(n_1973)
);

AOI21xp5_ASAP7_75t_L g1974 ( 
.A1(n_1962),
.A2(n_1901),
.B(n_1903),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1961),
.Y(n_1975)
);

INVx2_ASAP7_75t_SL g1976 ( 
.A(n_1964),
.Y(n_1976)
);

O2A1O1Ixp33_ASAP7_75t_L g1977 ( 
.A1(n_1963),
.A2(n_1921),
.B(n_1920),
.C(n_1919),
.Y(n_1977)
);

INVx3_ASAP7_75t_L g1978 ( 
.A(n_1976),
.Y(n_1978)
);

INVxp67_ASAP7_75t_SL g1979 ( 
.A(n_1977),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1975),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1972),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1974),
.Y(n_1982)
);

INVx1_ASAP7_75t_SL g1983 ( 
.A(n_1973),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_R g1984 ( 
.A(n_1978),
.B(n_1965),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_R g1985 ( 
.A(n_1978),
.B(n_1970),
.Y(n_1985)
);

OAI211xp5_ASAP7_75t_L g1986 ( 
.A1(n_1982),
.A2(n_1966),
.B(n_1968),
.C(n_1971),
.Y(n_1986)
);

AOI311xp33_ASAP7_75t_L g1987 ( 
.A1(n_1979),
.A2(n_1920),
.A3(n_1919),
.B(n_1836),
.C(n_1844),
.Y(n_1987)
);

INVx2_ASAP7_75t_SL g1988 ( 
.A(n_1978),
.Y(n_1988)
);

OAI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1986),
.A2(n_1982),
.B(n_1983),
.Y(n_1989)
);

NAND4xp75_ASAP7_75t_L g1990 ( 
.A(n_1988),
.B(n_1980),
.C(n_1981),
.D(n_1857),
.Y(n_1990)
);

NOR2x1_ASAP7_75t_L g1991 ( 
.A(n_1984),
.B(n_1981),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1991),
.B(n_1985),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1992),
.B(n_1917),
.Y(n_1993)
);

OR3x2_ASAP7_75t_L g1994 ( 
.A(n_1993),
.B(n_1980),
.C(n_1989),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1993),
.Y(n_1995)
);

AOI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1995),
.A2(n_1994),
.B1(n_1990),
.B2(n_1987),
.Y(n_1996)
);

INVx2_ASAP7_75t_SL g1997 ( 
.A(n_1995),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1997),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1996),
.A2(n_1876),
.B(n_1844),
.Y(n_1999)
);

OAI22x1_ASAP7_75t_L g2000 ( 
.A1(n_1998),
.A2(n_1852),
.B1(n_1805),
.B2(n_1608),
.Y(n_2000)
);

NAND3xp33_ASAP7_75t_L g2001 ( 
.A(n_2000),
.B(n_1999),
.C(n_1852),
.Y(n_2001)
);

OAI21xp5_ASAP7_75t_SL g2002 ( 
.A1(n_2001),
.A2(n_1852),
.B(n_1827),
.Y(n_2002)
);

CKINVDCx20_ASAP7_75t_R g2003 ( 
.A(n_2002),
.Y(n_2003)
);

OAI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_2003),
.A2(n_1850),
.B1(n_1858),
.B2(n_1862),
.Y(n_2004)
);

AOI211xp5_ASAP7_75t_L g2005 ( 
.A1(n_2004),
.A2(n_1852),
.B(n_1570),
.C(n_1817),
.Y(n_2005)
);


endmodule