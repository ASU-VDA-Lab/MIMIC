module fake_jpeg_20419_n_261 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_20),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_31),
.C(n_24),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_47),
.C(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_49),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_19),
.B1(n_28),
.B2(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_19),
.B1(n_28),
.B2(n_24),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_53),
.A2(n_65),
.B1(n_67),
.B2(n_44),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_61),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_28),
.B1(n_21),
.B2(n_25),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_63),
.B1(n_64),
.B2(n_18),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_20),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_59),
.B(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_29),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_25),
.B1(n_17),
.B2(n_23),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_25),
.B1(n_17),
.B2(n_23),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_29),
.B1(n_26),
.B2(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_34),
.B1(n_26),
.B2(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_31),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_96),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_68),
.C(n_50),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_74),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_38),
.C(n_37),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_81),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_78),
.A2(n_86),
.B1(n_103),
.B2(n_3),
.Y(n_125)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_82),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_33),
.B(n_27),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_51),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_84),
.Y(n_119)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_89),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_33),
.B1(n_46),
.B2(n_62),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_91),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_59),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_37),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_15),
.Y(n_117)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_97),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_61),
.A2(n_27),
.B1(n_30),
.B2(n_18),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_99),
.B1(n_56),
.B2(n_30),
.Y(n_107)
);

AND2x4_ASAP7_75t_SL g96 ( 
.A(n_53),
.B(n_38),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_67),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_48),
.A2(n_64),
.B1(n_27),
.B2(n_18),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_16),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_104),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g102 ( 
.A1(n_49),
.A2(n_44),
.B1(n_38),
.B2(n_37),
.Y(n_102)
);

AO22x1_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_57),
.A2(n_30),
.B1(n_34),
.B2(n_2),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_69),
.A2(n_44),
.B1(n_38),
.B2(n_34),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_111),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_38),
.B1(n_1),
.B2(n_2),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_69),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_130),
.Y(n_147)
);

AO22x1_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_96),
.B1(n_99),
.B2(n_102),
.Y(n_137)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_92),
.CI(n_102),
.CON(n_144),
.SN(n_144)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_73),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_6),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_7),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_74),
.C(n_70),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_126),
.C(n_106),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_87),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_124),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_152),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_138),
.B(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_93),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_143),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_96),
.B(n_95),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_146),
.B(n_154),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_110),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_124),
.C(n_105),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_145),
.B(n_151),
.Y(n_175)
);

OR2x6_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_92),
.Y(n_146)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_149),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_114),
.B(n_79),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_85),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_117),
.B(n_8),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_8),
.Y(n_179)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_152),
.B(n_144),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_124),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_180),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_129),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_169),
.B(n_178),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_176),
.C(n_181),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_108),
.B(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_116),
.B1(n_109),
.B2(n_107),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_172),
.A2(n_84),
.B1(n_80),
.B2(n_83),
.Y(n_200)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_154),
.A2(n_116),
.B1(n_122),
.B2(n_128),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_141),
.B1(n_133),
.B2(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_146),
.A2(n_126),
.B(n_115),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_179),
.B(n_182),
.Y(n_192)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_113),
.C(n_112),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_113),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_183),
.B(n_185),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_173),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_146),
.B(n_142),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_188),
.B(n_199),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_134),
.B(n_133),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_196),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_134),
.B1(n_137),
.B2(n_140),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_190),
.A2(n_170),
.B1(n_172),
.B2(n_159),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_170),
.A2(n_137),
.B1(n_144),
.B2(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_194),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_136),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_167),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_169),
.A2(n_150),
.B(n_112),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_200),
.A2(n_166),
.B1(n_171),
.B2(n_180),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_163),
.B(n_150),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_217),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_181),
.C(n_168),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_206),
.C(n_208),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_176),
.C(n_198),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_211),
.B1(n_200),
.B2(n_199),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_164),
.C(n_162),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_213),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_190),
.B1(n_195),
.B2(n_184),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_161),
.B(n_166),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_212),
.B(n_184),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_161),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_220),
.A2(n_213),
.B1(n_175),
.B2(n_94),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_187),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_221),
.A2(n_209),
.B1(n_211),
.B2(n_214),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_228),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_186),
.C(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

FAx1_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_183),
.CI(n_187),
.CON(n_227),
.SN(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_193),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_205),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_231),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_193),
.C(n_191),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_230),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_232),
.A2(n_233),
.B1(n_239),
.B2(n_227),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_207),
.B1(n_203),
.B2(n_204),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_233),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_89),
.B1(n_79),
.B2(n_11),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_241),
.A2(n_243),
.B1(n_244),
.B2(n_247),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_219),
.C(n_229),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_225),
.C(n_231),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_225),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_244),
.A2(n_232),
.B1(n_237),
.B2(n_245),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_13),
.B(n_14),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_242),
.A2(n_9),
.B(n_10),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_10),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_253),
.A2(n_256),
.B(n_248),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_251),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_255),
.C(n_13),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_12),
.C(n_13),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_258),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_14),
.B(n_15),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_15),
.Y(n_261)
);


endmodule