module fake_jpeg_24115_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_9),
.A2(n_0),
.B(n_2),
.C(n_4),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_17),
.A2(n_22),
.B1(n_13),
.B2(n_11),
.Y(n_35)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_21),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_13),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

OR2x4_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_0),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_32),
.B(n_10),
.Y(n_39)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_10),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_24),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_30),
.B1(n_32),
.B2(n_20),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_29),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_39),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_15),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_40),
.C(n_26),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_45),
.B(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_49),
.C(n_46),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_33),
.B(n_25),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

AOI322xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_40),
.A3(n_37),
.B1(n_31),
.B2(n_51),
.C1(n_41),
.C2(n_28),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_16),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_33),
.B(n_27),
.Y(n_55)
);


endmodule