module real_jpeg_27623_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx5_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_0),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_53),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_1),
.A2(n_53),
.B1(n_63),
.B2(n_64),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_1),
.A2(n_32),
.B1(n_34),
.B2(n_53),
.Y(n_158)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_3),
.A2(n_63),
.B1(n_64),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_3),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_143),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_143),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_3),
.A2(n_32),
.B1(n_34),
.B2(n_143),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_4),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_173),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_173),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_4),
.A2(n_32),
.B1(n_34),
.B2(n_173),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_7),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_56),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_7),
.A2(n_32),
.B1(n_34),
.B2(n_56),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_8),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_167),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_167),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_8),
.A2(n_32),
.B1(n_34),
.B2(n_167),
.Y(n_250)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_9),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_9),
.B(n_59),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_9),
.B(n_46),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_9),
.A2(n_46),
.B(n_210),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_171),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_9),
.A2(n_32),
.B(n_35),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_9),
.B(n_139),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_9),
.A2(n_87),
.B1(n_93),
.B2(n_258),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_10),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_66),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_10),
.A2(n_32),
.B1(n_34),
.B2(n_66),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_12),
.A2(n_32),
.B1(n_34),
.B2(n_38),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_12),
.A2(n_38),
.B1(n_63),
.B2(n_64),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_12),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_114)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_120),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_20),
.B(n_103),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_84),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_21),
.A2(n_22),
.B1(n_74),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_22)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_24),
.A2(n_25),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_24),
.B(n_40),
.C(n_57),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_36),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_26),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_26),
.A2(n_31),
.B1(n_98),
.B2(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_26),
.A2(n_36),
.B(n_99),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_26),
.A2(n_31),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_26),
.A2(n_79),
.B(n_218),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_26),
.A2(n_31),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_26),
.A2(n_31),
.B1(n_217),
.B2(n_235),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g208 ( 
.A1(n_28),
.A2(n_47),
.A3(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g211 ( 
.A(n_29),
.B(n_44),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_29),
.A2(n_30),
.B(n_171),
.C(n_237),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_31)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_31),
.A2(n_81),
.B(n_137),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_31),
.B(n_171),
.Y(n_256)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_34),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_34),
.B(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_37),
.B(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_51),
.B(n_54),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_41),
.A2(n_113),
.B(n_182),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_41),
.A2(n_54),
.B(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_50),
.B1(n_52),
.B2(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_42),
.B(n_55),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_42),
.A2(n_50),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_42),
.A2(n_50),
.B1(n_166),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_42),
.A2(n_50),
.B1(n_196),
.B2(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_43)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_44),
.Y(n_209)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_47),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_46),
.B(n_60),
.Y(n_185)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_47),
.A2(n_69),
.B1(n_170),
.B2(n_185),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_50),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_50),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_73),
.B1(n_105),
.B2(n_117),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_67),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_71),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_58),
.A2(n_62),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_58),
.A2(n_107),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_58),
.A2(n_107),
.B1(n_142),
.B2(n_179),
.Y(n_294)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_60),
.B(n_64),
.C(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_59),
.B(n_101),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_59),
.A2(n_68),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_64),
.Y(n_69)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g170 ( 
.A(n_64),
.B(n_171),
.CON(n_170),
.SN(n_170)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_74),
.A2(n_75),
.B(n_78),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_74),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_77),
.A2(n_115),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_84),
.A2(n_85),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_96),
.B(n_100),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_86),
.A2(n_100),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_86),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_86),
.A2(n_97),
.B1(n_126),
.B2(n_311),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_91),
.B(n_94),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_87),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_87),
.A2(n_91),
.B1(n_158),
.B2(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_87),
.A2(n_135),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_87),
.A2(n_250),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_88),
.A2(n_95),
.B(n_160),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_88),
.A2(n_92),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_95),
.Y(n_135)
);

INVx11_ASAP7_75t_L g259 ( 
.A(n_92),
.Y(n_259)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_93),
.B(n_134),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_93),
.A2(n_132),
.B(n_187),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_93),
.B(n_171),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_97),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_118),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_116),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_107),
.A2(n_142),
.B(n_144),
.Y(n_141)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_114),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_149),
.B(n_320),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_145),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_122),
.B(n_145),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.C(n_128),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_123),
.B(n_127),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_128),
.A2(n_129),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_138),
.C(n_140),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_130),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_131),
.B(n_136),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_138),
.A2(n_140),
.B1(n_141),
.B2(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_138),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_314),
.B(n_319),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_301),
.B(n_313),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_200),
.B(n_282),
.C(n_300),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_188),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_153),
.B(n_188),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_174),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_155),
.B(n_161),
.C(n_174),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_156),
.B(n_157),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_169),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_183),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_176),
.B(n_181),
.C(n_183),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_186),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_189),
.A2(n_190),
.B1(n_277),
.B2(n_279),
.Y(n_276)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_194),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.C(n_199),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_199),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_281),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_274),
.B(n_280),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_228),
.B(n_273),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_219),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_204),
.B(n_219),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_212),
.C(n_215),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_205),
.A2(n_206),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_208),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_220),
.B(n_226),
.C(n_227),
.Y(n_275)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_267),
.B(n_272),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_246),
.B(n_266),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_238),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_231),
.B(n_238),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_253),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_236),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_244),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_243),
.C(n_244),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_245),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_254),
.B(n_265),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_248),
.B(n_252),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_260),
.B(n_264),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_256),
.B(n_257),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_275),
.B(n_276),
.Y(n_280)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_277),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_284),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_298),
.B2(n_299),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_290),
.C(n_299),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_293),
.C(n_296),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_298),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_302),
.B(n_303),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_312),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_309),
.B2(n_310),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_310),
.C(n_312),
.Y(n_315)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);


endmodule