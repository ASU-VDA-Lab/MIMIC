module fake_netlist_5_2013_n_2227 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2227);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2227;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_2031;
wire n_556;
wire n_2076;
wire n_1728;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_314;
wire n_433;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_1138;
wire n_364;
wire n_927;
wire n_1089;
wire n_2044;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_3),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_109),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_41),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_59),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_81),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_56),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_111),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_50),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_157),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_33),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_84),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_120),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_219),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_150),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_162),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_137),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_19),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_20),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_170),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_208),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_179),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_17),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_163),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_141),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_46),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_41),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_2),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_27),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_72),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_160),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_15),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_45),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_113),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_184),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_16),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_121),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_175),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_168),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_53),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_92),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_94),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_61),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_4),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_6),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_183),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_216),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_176),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_127),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_116),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_115),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_145),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_172),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_129),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_146),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_169),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_98),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_60),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_90),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_164),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_87),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_73),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_85),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_152),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_173),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_104),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_155),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_87),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_197),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_147),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_124),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_74),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_213),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_199),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_83),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_165),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_6),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_51),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_48),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_81),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_46),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_23),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_61),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_15),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_29),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_32),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_18),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_132),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_158),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_58),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_82),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_159),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_212),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_17),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_80),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_50),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_142),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_18),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_161),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_112),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_68),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_84),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_118),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_123),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_95),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_66),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_186),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_51),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_189),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_37),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_106),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_153),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_68),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_102),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_220),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_214),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_70),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_31),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_48),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_3),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_117),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_72),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_215),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_177),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_43),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_134),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_91),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_211),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_149),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_37),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_217),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_26),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_108),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_143),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_206),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_56),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_22),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_130),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_22),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_79),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_54),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_107),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_24),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_154),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_144),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_78),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_171),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_20),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_205),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_86),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_19),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_125),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_93),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_210),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_11),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_122),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_21),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_221),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_148),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_83),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_35),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_209),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_192),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_4),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_140),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_194),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_26),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_30),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_79),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_181),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_77),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_14),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_110),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_80),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_33),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_55),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_201),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_198),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_12),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_126),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_13),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_166),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_45),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_174),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_34),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_180),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_85),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_139),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_103),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_182),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_38),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_75),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_43),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_101),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_7),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_58),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_0),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_10),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_14),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_82),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_78),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_30),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_59),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_44),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_187),
.Y(n_429)
);

BUFx5_ASAP7_75t_L g430 ( 
.A(n_10),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_185),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_96),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_40),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_2),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_11),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_55),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_255),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_231),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_430),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_430),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_256),
.B(n_0),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_430),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_430),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_430),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_359),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_430),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_430),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_430),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_236),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_430),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_228),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_375),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_248),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_375),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_237),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_359),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_375),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_238),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_242),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_368),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_297),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_243),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_228),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_267),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_267),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_375),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_380),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_375),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_405),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_368),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_247),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_405),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_285),
.B(n_1),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_259),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_262),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_417),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_263),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_265),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_405),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_266),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_271),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_275),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_276),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_405),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_224),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_417),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_L g487 ( 
.A(n_292),
.B(n_1),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_405),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_228),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_235),
.B(n_5),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_235),
.B(n_5),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_264),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_277),
.Y(n_493)
);

BUFx6f_ASAP7_75t_SL g494 ( 
.A(n_293),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_278),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_279),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_382),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_280),
.Y(n_498)
);

INVxp33_ASAP7_75t_SL g499 ( 
.A(n_226),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_429),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_264),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_284),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_225),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_302),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_273),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_302),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_341),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_308),
.B(n_7),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_289),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_341),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_225),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_273),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_381),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_362),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_381),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_362),
.Y(n_516)
);

INVxp33_ASAP7_75t_SL g517 ( 
.A(n_372),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_308),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_346),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_228),
.Y(n_520)
);

BUFx6f_ASAP7_75t_SL g521 ( 
.A(n_293),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_228),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_224),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_223),
.B(n_229),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_223),
.B(n_8),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_295),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_229),
.B(n_8),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_227),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_383),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_346),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_227),
.Y(n_531)
);

INVxp33_ASAP7_75t_L g532 ( 
.A(n_232),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_261),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_298),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_232),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_233),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_300),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_233),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_251),
.Y(n_539)
);

NOR2xp67_ASAP7_75t_L g540 ( 
.A(n_292),
.B(n_9),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_230),
.Y(n_541)
);

INVxp67_ASAP7_75t_SL g542 ( 
.A(n_240),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_313),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_234),
.B(n_9),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_316),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_317),
.Y(n_546)
);

CKINVDCx14_ASAP7_75t_R g547 ( 
.A(n_293),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_323),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_251),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_234),
.B(n_12),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_222),
.B(n_13),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_244),
.B(n_16),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_361),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_463),
.B(n_290),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_524),
.B(n_324),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_452),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_445),
.B(n_329),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_452),
.Y(n_558)
);

INVx6_ASAP7_75t_L g559 ( 
.A(n_460),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_456),
.B(n_331),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_454),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_450),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_508),
.B(n_272),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_508),
.B(n_290),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_463),
.B(n_312),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_553),
.B(n_361),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_533),
.B(n_293),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_454),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_463),
.B(n_312),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_438),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_470),
.B(n_428),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_451),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_460),
.B(n_428),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_490),
.B(n_333),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_450),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_457),
.B(n_335),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_457),
.B(n_336),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_466),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_463),
.Y(n_579)
);

BUFx8_ASAP7_75t_L g580 ( 
.A(n_494),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_451),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_466),
.B(n_355),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_533),
.B(n_386),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_468),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_460),
.Y(n_585)
);

BUFx8_ASAP7_75t_L g586 ( 
.A(n_494),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_468),
.B(n_340),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_469),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_451),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_449),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_450),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_469),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_472),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_489),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_489),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_489),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_520),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_472),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_479),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_479),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_484),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_520),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_484),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_488),
.B(n_350),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_485),
.B(n_244),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_520),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_522),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_522),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_522),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_519),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_488),
.B(n_352),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_439),
.B(n_272),
.Y(n_612)
);

OA21x2_ASAP7_75t_L g613 ( 
.A1(n_439),
.A2(n_249),
.B(n_245),
.Y(n_613)
);

OA21x2_ASAP7_75t_L g614 ( 
.A1(n_440),
.A2(n_249),
.B(n_245),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_503),
.B(n_386),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_440),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_523),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_485),
.B(n_258),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_442),
.B(n_355),
.Y(n_619)
);

AND2x2_ASAP7_75t_SL g620 ( 
.A(n_491),
.B(n_371),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_530),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_R g622 ( 
.A(n_499),
.B(n_239),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_523),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_442),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_SL g625 ( 
.A(n_486),
.B(n_379),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_517),
.A2(n_426),
.B1(n_422),
.B2(n_253),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_443),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_443),
.B(n_444),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_505),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_444),
.B(n_446),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_518),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_518),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_446),
.B(n_371),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_447),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_447),
.B(n_353),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_448),
.B(n_357),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_448),
.A2(n_378),
.B(n_270),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_487),
.B(n_378),
.Y(n_638)
);

CKINVDCx6p67_ASAP7_75t_R g639 ( 
.A(n_494),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_492),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_SL g641 ( 
.A(n_491),
.B(n_254),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_528),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_528),
.B(n_258),
.Y(n_643)
);

CKINVDCx8_ASAP7_75t_R g644 ( 
.A(n_503),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_L g645 ( 
.A(n_563),
.B(n_455),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_575),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_630),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_575),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_630),
.Y(n_649)
);

AO21x2_ASAP7_75t_L g650 ( 
.A1(n_635),
.A2(n_283),
.B(n_270),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_575),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_555),
.B(n_458),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_620),
.A2(n_441),
.B1(n_473),
.B2(n_547),
.Y(n_653)
);

INVxp33_ASAP7_75t_L g654 ( 
.A(n_610),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_573),
.B(n_437),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_630),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_573),
.B(n_486),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_555),
.B(n_459),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_570),
.B(n_462),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_635),
.B(n_471),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_559),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_559),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_630),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_630),
.Y(n_664)
);

AND2x2_ASAP7_75t_SL g665 ( 
.A(n_620),
.B(n_272),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_575),
.Y(n_666)
);

INVx5_ASAP7_75t_L g667 ( 
.A(n_563),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_616),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_616),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_557),
.B(n_474),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_559),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_629),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_636),
.B(n_475),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_591),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_616),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_562),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_624),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_591),
.Y(n_678)
);

INVxp67_ASAP7_75t_SL g679 ( 
.A(n_585),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_624),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_591),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_624),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_562),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_573),
.B(n_542),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_627),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_627),
.Y(n_686)
);

NAND3xp33_ASAP7_75t_SL g687 ( 
.A(n_625),
.B(n_514),
.C(n_512),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_625),
.B(n_541),
.C(n_478),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_562),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_641),
.A2(n_620),
.B1(n_622),
.B2(n_583),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_597),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_627),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_591),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_636),
.B(n_477),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_559),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_562),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_634),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_590),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_L g699 ( 
.A(n_571),
.B(n_481),
.C(n_480),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_634),
.Y(n_700)
);

BUFx4f_ASAP7_75t_L g701 ( 
.A(n_613),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_562),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_634),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_567),
.B(n_482),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_637),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_637),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_557),
.B(n_483),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_637),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_631),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_562),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_560),
.B(n_493),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_556),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_605),
.B(n_283),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_560),
.B(n_495),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_562),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_605),
.B(n_492),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_612),
.Y(n_717)
);

INVx5_ASAP7_75t_L g718 ( 
.A(n_563),
.Y(n_718)
);

INVx4_ASAP7_75t_L g719 ( 
.A(n_612),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_580),
.B(n_496),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_559),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_615),
.A2(n_534),
.B1(n_545),
.B2(n_543),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_556),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_558),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_572),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_597),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_644),
.Y(n_727)
);

BUFx10_ASAP7_75t_L g728 ( 
.A(n_564),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_572),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_558),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_572),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_644),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_561),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_597),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_564),
.A2(n_527),
.B1(n_544),
.B2(n_525),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_597),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_574),
.B(n_498),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_644),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_597),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_581),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_581),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_561),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_568),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_568),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_580),
.B(n_502),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_574),
.B(n_509),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_578),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_631),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_632),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_581),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_597),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_578),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_619),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_619),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_605),
.B(n_501),
.Y(n_755)
);

BUFx4f_ASAP7_75t_L g756 ( 
.A(n_613),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_619),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_589),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_L g759 ( 
.A(n_563),
.B(n_526),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_612),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_584),
.Y(n_761)
);

BUFx4f_ASAP7_75t_L g762 ( 
.A(n_613),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_584),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_621),
.A2(n_529),
.B1(n_546),
.B2(n_537),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_629),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_632),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_588),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_580),
.B(n_548),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_588),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_592),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_564),
.B(n_281),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_612),
.Y(n_772)
);

INVxp67_ASAP7_75t_SL g773 ( 
.A(n_628),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_589),
.Y(n_774)
);

AND2x6_ASAP7_75t_L g775 ( 
.A(n_564),
.B(n_272),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_592),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_589),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_618),
.B(n_501),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_580),
.B(n_511),
.Y(n_779)
);

NOR2x1p5_ASAP7_75t_L g780 ( 
.A(n_639),
.B(n_257),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_621),
.B(n_511),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_576),
.B(n_294),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_639),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_593),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_610),
.B(n_465),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_576),
.B(n_394),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_586),
.B(n_516),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_593),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_586),
.B(n_465),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_597),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_577),
.B(n_404),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_596),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_586),
.B(n_487),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_598),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_596),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_579),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_596),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_602),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_773),
.B(n_638),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_647),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_657),
.B(n_571),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_665),
.B(n_628),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_647),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_746),
.B(n_453),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_670),
.B(n_638),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_649),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_690),
.A2(n_618),
.B1(n_571),
.B2(n_566),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_649),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_656),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_656),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_665),
.B(n_619),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_707),
.B(n_638),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_663),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_663),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_664),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_664),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_712),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_652),
.B(n_461),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_665),
.A2(n_658),
.B1(n_737),
.B2(n_735),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_712),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_660),
.B(n_638),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_728),
.B(n_633),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_653),
.A2(n_694),
.B1(n_673),
.B2(n_711),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_723),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_714),
.A2(n_618),
.B1(n_566),
.B2(n_467),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_L g826 ( 
.A(n_796),
.B(n_563),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_753),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_L g828 ( 
.A(n_796),
.B(n_563),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_796),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_657),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_728),
.B(n_633),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_781),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_782),
.B(n_577),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_786),
.B(n_587),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_713),
.A2(n_639),
.B1(n_500),
.B2(n_497),
.Y(n_835)
);

NAND3x1_ASAP7_75t_L g836 ( 
.A(n_722),
.B(n_626),
.C(n_552),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_791),
.B(n_587),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_728),
.B(n_633),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_699),
.B(n_566),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_728),
.B(n_701),
.Y(n_840)
);

BUFx6f_ASAP7_75t_SL g841 ( 
.A(n_748),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_684),
.A2(n_655),
.B1(n_771),
.B2(n_713),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_684),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_701),
.A2(n_762),
.B(n_756),
.C(n_550),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_796),
.B(n_604),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_753),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_716),
.B(n_604),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_713),
.A2(n_563),
.B1(n_633),
.B2(n_614),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_723),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_701),
.B(n_272),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_L g851 ( 
.A(n_687),
.B(n_626),
.C(n_476),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_701),
.B(n_274),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_716),
.B(n_611),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_755),
.B(n_611),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_753),
.Y(n_855)
);

BUFx5_ASAP7_75t_L g856 ( 
.A(n_705),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_754),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_755),
.B(n_563),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_724),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_778),
.B(n_563),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_754),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_724),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_756),
.B(n_274),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_756),
.B(n_274),
.Y(n_864)
);

NAND2xp33_ASAP7_75t_L g865 ( 
.A(n_705),
.B(n_274),
.Y(n_865)
);

NOR3xp33_ASAP7_75t_L g866 ( 
.A(n_688),
.B(n_464),
.C(n_419),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_754),
.Y(n_867)
);

OAI22xp33_ASAP7_75t_L g868 ( 
.A1(n_713),
.A2(n_540),
.B1(n_291),
.B2(n_321),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_756),
.B(n_274),
.Y(n_869)
);

NAND2x1p5_ASAP7_75t_L g870 ( 
.A(n_757),
.B(n_667),
.Y(n_870)
);

INVxp67_ASAP7_75t_L g871 ( 
.A(n_709),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_709),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_757),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_757),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_778),
.B(n_679),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_730),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_654),
.B(n_494),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_730),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_733),
.B(n_579),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_733),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_713),
.A2(n_614),
.B1(n_613),
.B2(n_643),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_742),
.B(n_643),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_742),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_743),
.B(n_643),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_661),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_743),
.B(n_643),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_744),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_744),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_747),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_L g890 ( 
.A(n_706),
.B(n_339),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_747),
.B(n_643),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_752),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_752),
.B(n_613),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_655),
.A2(n_418),
.B1(n_366),
.B2(n_369),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_761),
.B(n_614),
.Y(n_895)
);

NAND2x1_ASAP7_75t_L g896 ( 
.A(n_717),
.B(n_612),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_764),
.B(n_521),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_766),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_659),
.B(n_521),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_761),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_762),
.B(n_339),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_763),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_704),
.B(n_521),
.Y(n_903)
);

NAND2x1_ASAP7_75t_L g904 ( 
.A(n_717),
.B(n_612),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_748),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_763),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_767),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_762),
.B(n_339),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_767),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_769),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_762),
.B(n_339),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_749),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_769),
.B(n_770),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_661),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_667),
.B(n_339),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_770),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_776),
.B(n_614),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_698),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_776),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_784),
.B(n_788),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_749),
.B(n_521),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_784),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_788),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_661),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_794),
.B(n_614),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_645),
.A2(n_623),
.B(n_642),
.C(n_617),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_667),
.B(n_406),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_785),
.B(n_532),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_794),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_785),
.B(n_551),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_650),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_672),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_668),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_669),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_727),
.B(n_551),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_650),
.B(n_569),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_650),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_706),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_793),
.B(n_241),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_669),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_675),
.Y(n_941)
);

BUFx8_ASAP7_75t_L g942 ( 
.A(n_775),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_759),
.A2(n_623),
.B(n_642),
.C(n_617),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_696),
.B(n_569),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_765),
.B(n_531),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_708),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_708),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_783),
.B(n_531),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_696),
.B(n_569),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_720),
.B(n_246),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_662),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_696),
.B(n_569),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_702),
.B(n_554),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_675),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_745),
.B(n_250),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_667),
.B(n_406),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_702),
.B(n_721),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_768),
.B(n_252),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_721),
.A2(n_565),
.B(n_554),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_702),
.B(n_676),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_789),
.B(n_268),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_677),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_667),
.B(n_406),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_780),
.A2(n_373),
.B1(n_387),
.B2(n_358),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_677),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_680),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_662),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_680),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_662),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_800),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_829),
.A2(n_695),
.B(n_671),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_800),
.Y(n_972)
);

NOR2x1p5_ASAP7_75t_L g973 ( 
.A(n_918),
.B(n_779),
.Y(n_973)
);

NOR2xp67_ASAP7_75t_L g974 ( 
.A(n_932),
.B(n_787),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_832),
.B(n_732),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_829),
.B(n_667),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_833),
.B(n_676),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_829),
.A2(n_695),
.B(n_671),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_834),
.B(n_837),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_819),
.A2(n_685),
.B(n_686),
.C(n_682),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_822),
.A2(n_695),
.B(n_671),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_805),
.B(n_676),
.Y(n_982)
);

INVxp67_ASAP7_75t_SL g983 ( 
.A(n_827),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_823),
.A2(n_775),
.B1(n_780),
.B2(n_738),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_822),
.A2(n_715),
.B(n_718),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_930),
.B(n_945),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_812),
.B(n_676),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_L g988 ( 
.A1(n_830),
.A2(n_282),
.B(n_269),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_L g989 ( 
.A(n_804),
.B(n_540),
.C(n_291),
.Y(n_989)
);

AOI21x1_ASAP7_75t_L g990 ( 
.A1(n_850),
.A2(n_685),
.B(n_682),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_806),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_801),
.B(n_535),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_831),
.A2(n_715),
.B(n_718),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_799),
.B(n_683),
.Y(n_994)
);

NAND2x1_ASAP7_75t_L g995 ( 
.A(n_885),
.B(n_715),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_843),
.B(n_535),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_839),
.A2(n_775),
.B1(n_689),
.B2(n_710),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_842),
.A2(n_288),
.B(n_327),
.C(n_321),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_847),
.B(n_853),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_843),
.B(n_718),
.Y(n_1000)
);

AOI21x1_ASAP7_75t_L g1001 ( 
.A1(n_850),
.A2(n_692),
.B(n_686),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_854),
.B(n_683),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_861),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_821),
.B(n_683),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_861),
.B(n_718),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_831),
.A2(n_715),
.B(n_718),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_871),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_852),
.A2(n_697),
.B(n_692),
.Y(n_1008)
);

NOR2x1_ASAP7_75t_R g1009 ( 
.A(n_918),
.B(n_286),
.Y(n_1009)
);

NOR3xp33_ASAP7_75t_L g1010 ( 
.A(n_818),
.B(n_327),
.C(n_288),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_872),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_838),
.A2(n_718),
.B(n_717),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_838),
.A2(n_719),
.B(n_717),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_845),
.A2(n_760),
.B(n_719),
.Y(n_1014)
);

BUFx4_ASAP7_75t_SL g1015 ( 
.A(n_878),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_826),
.A2(n_760),
.B(n_719),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_875),
.B(n_683),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_807),
.A2(n_775),
.B1(n_710),
.B2(n_689),
.Y(n_1018)
);

NOR2x1_ASAP7_75t_L g1019 ( 
.A(n_835),
.B(n_719),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_883),
.B(n_689),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_887),
.B(n_689),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_861),
.B(n_760),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_888),
.B(n_710),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_928),
.B(n_536),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_802),
.A2(n_700),
.B(n_703),
.C(n_697),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_802),
.A2(n_296),
.B1(n_299),
.B2(n_257),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_948),
.B(n_536),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_809),
.Y(n_1028)
);

NAND2x1_ASAP7_75t_L g1029 ( 
.A(n_885),
.B(n_710),
.Y(n_1029)
);

AOI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_961),
.A2(n_586),
.B(n_338),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_825),
.B(n_260),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_889),
.B(n_700),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_898),
.B(n_538),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_902),
.B(n_703),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_826),
.A2(n_772),
.B(n_760),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_861),
.B(n_772),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_828),
.A2(n_772),
.B(n_734),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_905),
.B(n_332),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_907),
.B(n_646),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_828),
.A2(n_772),
.B(n_734),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_905),
.B(n_344),
.Y(n_1041)
);

AND2x6_ASAP7_75t_L g1042 ( 
.A(n_938),
.B(n_328),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_885),
.A2(n_734),
.B(n_691),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_924),
.A2(n_863),
.B(n_852),
.Y(n_1044)
);

AO21x1_ASAP7_75t_L g1045 ( 
.A1(n_863),
.A2(n_338),
.B(n_328),
.Y(n_1045)
);

OAI21xp33_ASAP7_75t_SL g1046 ( 
.A1(n_811),
.A2(n_347),
.B(n_345),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_931),
.A2(n_296),
.B1(n_306),
.B2(n_299),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_873),
.B(n_815),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_924),
.A2(n_734),
.B(n_691),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_909),
.B(n_646),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_844),
.A2(n_347),
.B1(n_348),
.B2(n_345),
.Y(n_1051)
);

AOI33xp33_ASAP7_75t_L g1052 ( 
.A1(n_912),
.A2(n_374),
.A3(n_349),
.B1(n_318),
.B2(n_310),
.B3(n_307),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_816),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_816),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_924),
.A2(n_734),
.B(n_691),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_864),
.A2(n_901),
.B(n_869),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_864),
.A2(n_648),
.B(n_646),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_841),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_931),
.A2(n_307),
.B1(n_310),
.B2(n_306),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_939),
.A2(n_348),
.B(n_376),
.C(n_351),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_916),
.B(n_648),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_922),
.B(n_648),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_869),
.A2(n_734),
.B(n_691),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_929),
.B(n_651),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_803),
.B(n_651),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_935),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_808),
.B(n_651),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_873),
.Y(n_1068)
);

AOI21x1_ASAP7_75t_L g1069 ( 
.A1(n_908),
.A2(n_674),
.B(n_666),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_950),
.A2(n_351),
.B(n_376),
.C(n_377),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_L g1071 ( 
.A(n_955),
.B(n_397),
.C(n_377),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_911),
.A2(n_736),
.B(n_726),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_810),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_813),
.B(n_814),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_873),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_817),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_913),
.B(n_367),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_811),
.A2(n_412),
.B(n_408),
.C(n_397),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_920),
.B(n_666),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_894),
.B(n_391),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_817),
.B(n_666),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_820),
.B(n_674),
.Y(n_1082)
);

AO21x1_ASAP7_75t_L g1083 ( 
.A1(n_865),
.A2(n_412),
.B(n_408),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_836),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_820),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_873),
.B(n_736),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_824),
.B(n_674),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_824),
.B(n_678),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_840),
.A2(n_739),
.B(n_736),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_849),
.B(n_678),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_958),
.A2(n_432),
.B(n_681),
.C(n_678),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_827),
.B(n_538),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_841),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_844),
.A2(n_432),
.B1(n_415),
.B2(n_693),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_967),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_849),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_840),
.A2(n_751),
.B(n_739),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_859),
.B(n_681),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_846),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_862),
.B(n_693),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_862),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_876),
.B(n_693),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_937),
.A2(n_349),
.B(n_435),
.C(n_318),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_876),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_855),
.A2(n_857),
.B1(n_874),
.B2(n_867),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_880),
.B(n_892),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_881),
.A2(n_895),
.B(n_893),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_880),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_892),
.B(n_775),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_858),
.A2(n_790),
.B(n_751),
.C(n_582),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_827),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_836),
.A2(n_775),
.B1(n_790),
.B2(n_554),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_856),
.B(n_790),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_914),
.Y(n_1114)
);

NOR3xp33_ASAP7_75t_L g1115 ( 
.A(n_897),
.B(n_301),
.C(n_287),
.Y(n_1115)
);

AND2x6_ASAP7_75t_L g1116 ( 
.A(n_946),
.B(n_790),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_944),
.A2(n_565),
.B(n_554),
.Y(n_1117)
);

O2A1O1Ixp5_ASAP7_75t_L g1118 ( 
.A1(n_900),
.A2(n_582),
.B(n_565),
.C(n_554),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_900),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_914),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_856),
.B(n_406),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_906),
.B(n_775),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_949),
.A2(n_565),
.B(n_725),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_906),
.B(n_775),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_910),
.B(n_303),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_866),
.B(n_539),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_919),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_919),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_923),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_952),
.A2(n_565),
.B(n_725),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_917),
.A2(n_729),
.B(n_725),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_957),
.A2(n_731),
.B(n_729),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_923),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_877),
.B(n_539),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_841),
.B(n_304),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_925),
.A2(n_731),
.B(n_729),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_953),
.A2(n_740),
.B(n_731),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_860),
.A2(n_937),
.B(n_936),
.Y(n_1138)
);

NOR2xp67_ASAP7_75t_L g1139 ( 
.A(n_899),
.B(n_549),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_868),
.A2(n_598),
.B(n_599),
.C(n_600),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_851),
.B(n_305),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_865),
.A2(n_741),
.B(n_740),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_856),
.B(n_406),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_914),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_882),
.B(n_740),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_856),
.B(n_798),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_884),
.B(n_741),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_964),
.Y(n_1148)
);

AOI33xp33_ASAP7_75t_L g1149 ( 
.A1(n_848),
.A2(n_360),
.A3(n_407),
.B1(n_409),
.B2(n_399),
.B3(n_416),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_886),
.B(n_741),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_891),
.A2(n_758),
.B(n_750),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_979),
.B(n_921),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_999),
.B(n_903),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_972),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1007),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1053),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1129),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1054),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1056),
.A2(n_890),
.B(n_926),
.C(n_943),
.Y(n_1159)
);

OAI21xp33_ASAP7_75t_SL g1160 ( 
.A1(n_1107),
.A2(n_947),
.B(n_879),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1138),
.B(n_1068),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1010),
.A2(n_890),
.B(n_968),
.C(n_962),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1077),
.B(n_549),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1015),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1044),
.A2(n_947),
.B(n_870),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_992),
.B(n_933),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1026),
.A2(n_954),
.B(n_934),
.C(n_966),
.Y(n_1167)
);

NOR2xp67_ASAP7_75t_L g1168 ( 
.A(n_986),
.B(n_933),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1016),
.A2(n_870),
.B(n_896),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1096),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1027),
.B(n_1129),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1026),
.A2(n_1077),
.B(n_1031),
.C(n_1080),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1035),
.A2(n_904),
.B(n_959),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1104),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1119),
.Y(n_1175)
);

AOI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1048),
.A2(n_960),
.B(n_940),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1084),
.A2(n_934),
.B1(n_940),
.B2(n_966),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1134),
.B(n_941),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1011),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1141),
.A2(n_941),
.B(n_965),
.C(n_364),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1004),
.A2(n_951),
.B(n_914),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1127),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1024),
.B(n_965),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_970),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1141),
.A2(n_360),
.B(n_364),
.C(n_435),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_991),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1111),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_996),
.B(n_967),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1070),
.A2(n_374),
.B(n_434),
.C(n_427),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1133),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1068),
.B(n_856),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1071),
.A2(n_384),
.B(n_434),
.C(n_427),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1014),
.A2(n_976),
.B(n_982),
.Y(n_1193)
);

AOI221xp5_ASAP7_75t_L g1194 ( 
.A1(n_1031),
.A2(n_334),
.B1(n_311),
.B2(n_314),
.C(n_315),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1068),
.B(n_856),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1128),
.B(n_856),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1068),
.B(n_951),
.Y(n_1197)
);

AO21x1_ASAP7_75t_L g1198 ( 
.A1(n_1051),
.A2(n_927),
.B(n_915),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_996),
.B(n_969),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1148),
.A2(n_969),
.B1(n_951),
.B2(n_390),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1089),
.A2(n_927),
.B(n_915),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1015),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1073),
.B(n_951),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1028),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1066),
.B(n_504),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_1003),
.B(n_956),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_976),
.A2(n_963),
.B(n_956),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_987),
.A2(n_963),
.B(n_758),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1110),
.A2(n_758),
.B(n_750),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_SL g1211 ( 
.A(n_1115),
.B(n_319),
.C(n_309),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1092),
.B(n_942),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1022),
.A2(n_774),
.B(n_750),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1076),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1092),
.B(n_942),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_977),
.B(n_942),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_973),
.B(n_504),
.Y(n_1217)
);

OAI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_1080),
.A2(n_322),
.B(n_320),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1038),
.B(n_506),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1085),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1101),
.Y(n_1221)
);

OR2x6_ASAP7_75t_L g1222 ( 
.A(n_974),
.B(n_384),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1125),
.B(n_640),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_975),
.B(n_325),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1022),
.A2(n_777),
.B(n_774),
.Y(n_1225)
);

BUFx12f_ASAP7_75t_L g1226 ( 
.A(n_1058),
.Y(n_1226)
);

BUFx12f_ASAP7_75t_L g1227 ( 
.A(n_1093),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1149),
.A2(n_393),
.B(n_395),
.C(n_396),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1125),
.B(n_640),
.Y(n_1229)
);

AOI221xp5_ASAP7_75t_L g1230 ( 
.A1(n_1041),
.A2(n_411),
.B1(n_330),
.B2(n_337),
.C(n_342),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_998),
.A2(n_421),
.B(n_393),
.C(n_395),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1036),
.A2(n_994),
.B(n_1013),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1108),
.B(n_640),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1097),
.A2(n_798),
.B(n_797),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1099),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1106),
.Y(n_1236)
);

OAI21xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1074),
.A2(n_416),
.B(n_396),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1114),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_975),
.B(n_1099),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1126),
.B(n_506),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1139),
.B(n_774),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1060),
.A2(n_421),
.B(n_409),
.C(n_407),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1032),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1034),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1039),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1050),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1061),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1047),
.A2(n_399),
.B(n_326),
.C(n_424),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1036),
.A2(n_798),
.B(n_797),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_971),
.A2(n_797),
.B(n_795),
.Y(n_1250)
);

BUFx8_ASAP7_75t_L g1251 ( 
.A(n_1033),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_984),
.B(n_343),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1030),
.A2(n_603),
.B(n_601),
.C(n_600),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_978),
.A2(n_795),
.B(n_792),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1062),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1002),
.B(n_640),
.Y(n_1256)
);

OR2x6_ASAP7_75t_SL g1257 ( 
.A(n_1094),
.B(n_354),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1047),
.B(n_582),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1064),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1111),
.Y(n_1260)
);

NOR2xp67_ASAP7_75t_L g1261 ( 
.A(n_1135),
.B(n_389),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1037),
.A2(n_795),
.B(n_792),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1114),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1059),
.A2(n_356),
.B(n_363),
.C(n_365),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1040),
.A2(n_792),
.B(n_777),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_995),
.A2(n_1147),
.B(n_1145),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1059),
.B(n_582),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1150),
.A2(n_777),
.B(n_582),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1135),
.B(n_507),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_SL g1270 ( 
.A(n_989),
.B(n_392),
.C(n_388),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_988),
.Y(n_1271)
);

OAI22x1_ASAP7_75t_L g1272 ( 
.A1(n_1105),
.A2(n_400),
.B1(n_398),
.B2(n_385),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1095),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1052),
.A2(n_425),
.B(n_370),
.C(n_436),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1009),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1095),
.B(n_599),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1043),
.A2(n_594),
.B(n_595),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1019),
.A2(n_413),
.B1(n_401),
.B2(n_402),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1017),
.B(n_601),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1048),
.B(n_403),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1003),
.B(n_1075),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1103),
.A2(n_433),
.B(n_423),
.C(n_420),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1103),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1078),
.A2(n_513),
.B(n_515),
.C(n_510),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1112),
.A2(n_410),
.B1(n_414),
.B2(n_431),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1081),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1075),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1114),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1046),
.A2(n_1091),
.B(n_1140),
.C(n_1023),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_983),
.B(n_603),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1114),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1120),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1079),
.B(n_602),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1049),
.A2(n_595),
.B(n_594),
.Y(n_1294)
);

NOR3xp33_ASAP7_75t_L g1295 ( 
.A(n_1118),
.B(n_507),
.C(n_510),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1055),
.A2(n_594),
.B(n_595),
.Y(n_1296)
);

O2A1O1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1020),
.A2(n_513),
.B(n_515),
.C(n_607),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1082),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1021),
.B(n_21),
.Y(n_1299)
);

OAI221xp5_ASAP7_75t_L g1300 ( 
.A1(n_1018),
.A2(n_997),
.B1(n_1117),
.B2(n_1067),
.C(n_1065),
.Y(n_1300)
);

NAND3xp33_ASAP7_75t_SL g1301 ( 
.A(n_1083),
.B(n_386),
.C(n_608),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_980),
.A2(n_609),
.B(n_608),
.C(n_607),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1008),
.A2(n_606),
.B1(n_609),
.B2(n_608),
.Y(n_1303)
);

NOR2x1_ASAP7_75t_L g1304 ( 
.A(n_1144),
.B(n_594),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_981),
.A2(n_595),
.B(n_609),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1087),
.B(n_23),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1100),
.B(n_602),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1088),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1100),
.B(n_386),
.Y(n_1309)
);

NAND2x1p5_ASAP7_75t_L g1310 ( 
.A(n_1144),
.B(n_606),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1120),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1120),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1157),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1172),
.B(n_1086),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1155),
.Y(n_1315)
);

INVx3_ASAP7_75t_SL g1316 ( 
.A(n_1164),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1157),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1152),
.B(n_1042),
.Y(n_1318)
);

OR2x6_ASAP7_75t_L g1319 ( 
.A(n_1212),
.B(n_1120),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1172),
.A2(n_1025),
.B(n_1130),
.C(n_1123),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_SL g1321 ( 
.A1(n_1153),
.A2(n_1143),
.B(n_1121),
.C(n_1000),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1152),
.B(n_1042),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1234),
.A2(n_1069),
.B(n_1001),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1160),
.A2(n_1137),
.B(n_1132),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1179),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1171),
.B(n_1090),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1238),
.Y(n_1327)
);

AO31x2_ASAP7_75t_L g1328 ( 
.A1(n_1198),
.A2(n_1045),
.A3(n_1063),
.B(n_1142),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_1251),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1238),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1235),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1243),
.B(n_1042),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1165),
.A2(n_990),
.B(n_1072),
.Y(n_1333)
);

AOI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1161),
.A2(n_1121),
.B(n_1143),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1185),
.A2(n_1000),
.B(n_1086),
.C(n_1122),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1239),
.B(n_1042),
.Y(n_1336)
);

AO21x2_ASAP7_75t_L g1337 ( 
.A1(n_1161),
.A2(n_1151),
.B(n_1136),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1207),
.B(n_1042),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1244),
.B(n_1098),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1251),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1263),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1292),
.Y(n_1342)
);

AOI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1232),
.A2(n_1266),
.B(n_1176),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1236),
.B(n_1102),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1239),
.B(n_1109),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1201),
.A2(n_1057),
.B(n_1131),
.Y(n_1346)
);

OR2x6_ASAP7_75t_L g1347 ( 
.A(n_1215),
.B(n_1005),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1226),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1173),
.A2(n_1012),
.B(n_1113),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1159),
.A2(n_1146),
.B(n_1124),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1236),
.B(n_1116),
.Y(n_1351)
);

O2A1O1Ixp5_ASAP7_75t_SL g1352 ( 
.A1(n_1241),
.A2(n_1146),
.B(n_1113),
.C(n_1005),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1250),
.A2(n_1029),
.B(n_1006),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1177),
.A2(n_1257),
.B1(n_1178),
.B2(n_1283),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1300),
.A2(n_993),
.B(n_985),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1169),
.A2(n_1116),
.B(n_607),
.Y(n_1356)
);

BUFx8_ASAP7_75t_SL g1357 ( 
.A(n_1227),
.Y(n_1357)
);

A2O1A1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1252),
.A2(n_1116),
.B(n_606),
.C(n_27),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_SL g1359 ( 
.A1(n_1228),
.A2(n_1116),
.B(n_218),
.C(n_207),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1159),
.A2(n_1116),
.B(n_612),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1202),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1163),
.B(n_24),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1245),
.B(n_612),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1224),
.A2(n_25),
.B(n_28),
.C(n_29),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1275),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1168),
.B(n_25),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1177),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1254),
.A2(n_136),
.B(n_203),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1223),
.A2(n_612),
.B(n_202),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1271),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1229),
.A2(n_200),
.B(n_196),
.Y(n_1371)
);

NOR2xp67_ASAP7_75t_L g1372 ( 
.A(n_1211),
.B(n_195),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1224),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1218),
.B(n_36),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1262),
.A2(n_193),
.B(n_190),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1210),
.A2(n_188),
.B(n_156),
.Y(n_1376)
);

NOR2xp67_ASAP7_75t_L g1377 ( 
.A(n_1200),
.B(n_1280),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1167),
.A2(n_38),
.A3(n_39),
.B(n_40),
.Y(n_1378)
);

AO31x2_ASAP7_75t_L g1379 ( 
.A1(n_1167),
.A2(n_39),
.A3(n_42),
.B(n_44),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1181),
.A2(n_151),
.B(n_138),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1246),
.B(n_42),
.Y(n_1381)
);

AOI221xp5_ASAP7_75t_L g1382 ( 
.A1(n_1194),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.C(n_53),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1216),
.A2(n_135),
.B(n_133),
.Y(n_1383)
);

OR2x6_ASAP7_75t_L g1384 ( 
.A(n_1188),
.B(n_131),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1269),
.B(n_47),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1247),
.B(n_49),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1205),
.B(n_52),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1263),
.Y(n_1388)
);

BUFx12f_ASAP7_75t_L g1389 ( 
.A(n_1311),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1209),
.A2(n_128),
.B(n_119),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1166),
.A2(n_114),
.B(n_105),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1255),
.B(n_54),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1183),
.A2(n_100),
.B(n_99),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1240),
.B(n_57),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1259),
.B(n_57),
.Y(n_1395)
);

INVx6_ASAP7_75t_L g1396 ( 
.A(n_1217),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_SL g1397 ( 
.A(n_1222),
.Y(n_1397)
);

BUFx12f_ASAP7_75t_L g1398 ( 
.A(n_1312),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1265),
.A2(n_97),
.B(n_89),
.Y(n_1399)
);

INVx6_ASAP7_75t_SL g1400 ( 
.A(n_1222),
.Y(n_1400)
);

AO32x2_ASAP7_75t_L g1401 ( 
.A1(n_1303),
.A2(n_60),
.A3(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1188),
.B(n_62),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1260),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1187),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1273),
.B(n_88),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1268),
.A2(n_63),
.B(n_64),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1261),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_1407)
);

BUFx4f_ASAP7_75t_SL g1408 ( 
.A(n_1217),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1260),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1213),
.A2(n_1249),
.B(n_1225),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1219),
.B(n_1222),
.Y(n_1411)
);

AO31x2_ASAP7_75t_L g1412 ( 
.A1(n_1282),
.A2(n_65),
.A3(n_67),
.B(n_69),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1154),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1256),
.A2(n_69),
.B(n_70),
.Y(n_1414)
);

AOI221xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1248),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.C(n_75),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1308),
.B(n_71),
.Y(n_1416)
);

AO31x2_ASAP7_75t_L g1417 ( 
.A1(n_1282),
.A2(n_76),
.A3(n_77),
.B(n_86),
.Y(n_1417)
);

AO31x2_ASAP7_75t_L g1418 ( 
.A1(n_1228),
.A2(n_76),
.A3(n_1284),
.B(n_1299),
.Y(n_1418)
);

AO31x2_ASAP7_75t_L g1419 ( 
.A1(n_1284),
.A2(n_1299),
.A3(n_1274),
.B(n_1208),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1180),
.A2(n_1289),
.B(n_1280),
.C(n_1264),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1305),
.A2(n_1195),
.B(n_1191),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1298),
.B(n_1286),
.Y(n_1422)
);

AO32x2_ASAP7_75t_L g1423 ( 
.A1(n_1291),
.A2(n_1287),
.A3(n_1231),
.B1(n_1274),
.B2(n_1301),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1307),
.A2(n_1279),
.B(n_1293),
.Y(n_1424)
);

AO31x2_ASAP7_75t_L g1425 ( 
.A1(n_1248),
.A2(n_1264),
.A3(n_1277),
.B(n_1294),
.Y(n_1425)
);

NOR3xp33_ASAP7_75t_SL g1426 ( 
.A(n_1270),
.B(n_1237),
.C(n_1230),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1286),
.B(n_1187),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1199),
.B(n_1306),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1309),
.B(n_1272),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_1288),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1288),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1191),
.A2(n_1195),
.B(n_1162),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_SL g1433 ( 
.A1(n_1192),
.A2(n_1285),
.B(n_1278),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1296),
.A2(n_1302),
.B(n_1241),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1196),
.B(n_1214),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1184),
.A2(n_1220),
.B1(n_1186),
.B2(n_1204),
.Y(n_1436)
);

O2A1O1Ixp33_ASAP7_75t_SL g1437 ( 
.A1(n_1197),
.A2(n_1203),
.B(n_1267),
.C(n_1258),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1221),
.B(n_1154),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1156),
.A2(n_1158),
.B1(n_1170),
.B2(n_1174),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1295),
.A2(n_1253),
.B(n_1297),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1197),
.A2(n_1310),
.B(n_1304),
.Y(n_1441)
);

INVx5_ASAP7_75t_L g1442 ( 
.A(n_1156),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1290),
.A2(n_1276),
.B(n_1281),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1281),
.A2(n_1233),
.B(n_1231),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1170),
.B(n_1175),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1189),
.A2(n_1242),
.B(n_1182),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1206),
.A2(n_1175),
.B(n_1182),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1190),
.B(n_979),
.Y(n_1448)
);

INVx3_ASAP7_75t_SL g1449 ( 
.A(n_1190),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1157),
.Y(n_1450)
);

AO31x2_ASAP7_75t_L g1451 ( 
.A1(n_1198),
.A2(n_1159),
.A3(n_1051),
.B(n_1083),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1157),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1207),
.B(n_1077),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1234),
.A2(n_1165),
.B(n_1176),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1172),
.A2(n_1160),
.B(n_819),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1152),
.B(n_979),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1155),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1172),
.A2(n_804),
.B1(n_818),
.B2(n_1080),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1172),
.A2(n_1160),
.B(n_819),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1157),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1234),
.A2(n_1165),
.B(n_1176),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1155),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1157),
.Y(n_1463)
);

OAI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1172),
.A2(n_1031),
.B1(n_804),
.B2(n_1080),
.C(n_979),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1157),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1157),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1207),
.B(n_1077),
.Y(n_1467)
);

BUFx12f_ASAP7_75t_L g1468 ( 
.A(n_1164),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1173),
.A2(n_829),
.B(n_979),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1155),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1155),
.Y(n_1471)
);

AOI221x1_ASAP7_75t_L g1472 ( 
.A1(n_1172),
.A2(n_1030),
.B1(n_1071),
.B2(n_1010),
.C(n_1051),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1152),
.B(n_979),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1159),
.A2(n_1193),
.B(n_1161),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1207),
.B(n_1077),
.Y(n_1475)
);

AO31x2_ASAP7_75t_L g1476 ( 
.A1(n_1198),
.A2(n_1159),
.A3(n_1051),
.B(n_1083),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1188),
.B(n_1168),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1173),
.A2(n_829),
.B(n_1056),
.Y(n_1478)
);

AO31x2_ASAP7_75t_L g1479 ( 
.A1(n_1198),
.A2(n_1159),
.A3(n_1051),
.B(n_1083),
.Y(n_1479)
);

OAI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1458),
.A2(n_1464),
.B1(n_1367),
.B2(n_1473),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1427),
.Y(n_1481)
);

INVx8_ASAP7_75t_L g1482 ( 
.A(n_1389),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1427),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1464),
.A2(n_1382),
.B1(n_1374),
.B2(n_1385),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1327),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1377),
.A2(n_1453),
.B1(n_1475),
.B2(n_1467),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1403),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_SL g1488 ( 
.A1(n_1382),
.A2(n_1433),
.B(n_1407),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1398),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1357),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1409),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1411),
.A2(n_1429),
.B1(n_1336),
.B2(n_1354),
.Y(n_1492)
);

CKINVDCx11_ASAP7_75t_R g1493 ( 
.A(n_1329),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1456),
.A2(n_1473),
.B1(n_1428),
.B2(n_1354),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1367),
.A2(n_1459),
.B1(n_1455),
.B2(n_1456),
.Y(n_1495)
);

INVx8_ASAP7_75t_L g1496 ( 
.A(n_1342),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1397),
.A2(n_1387),
.B1(n_1459),
.B2(n_1455),
.Y(n_1497)
);

OAI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1362),
.A2(n_1395),
.B1(n_1381),
.B2(n_1386),
.Y(n_1498)
);

INVx5_ASAP7_75t_L g1499 ( 
.A(n_1384),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1342),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1314),
.A2(n_1366),
.B1(n_1397),
.B2(n_1414),
.Y(n_1501)
);

CKINVDCx11_ASAP7_75t_R g1502 ( 
.A(n_1316),
.Y(n_1502)
);

BUFx8_ASAP7_75t_SL g1503 ( 
.A(n_1468),
.Y(n_1503)
);

CKINVDCx11_ASAP7_75t_R g1504 ( 
.A(n_1365),
.Y(n_1504)
);

OAI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1381),
.A2(n_1392),
.B1(n_1386),
.B2(n_1395),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1392),
.A2(n_1416),
.B1(n_1394),
.B2(n_1406),
.Y(n_1506)
);

OAI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1472),
.A2(n_1416),
.B1(n_1384),
.B2(n_1433),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1327),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1315),
.Y(n_1509)
);

INVx6_ASAP7_75t_L g1510 ( 
.A(n_1342),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1420),
.A2(n_1318),
.B1(n_1322),
.B2(n_1449),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1338),
.A2(n_1322),
.B1(n_1318),
.B2(n_1400),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1400),
.A2(n_1347),
.B1(n_1332),
.B2(n_1402),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_SL g1514 ( 
.A1(n_1364),
.A2(n_1373),
.B(n_1358),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1457),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1347),
.A2(n_1332),
.B1(n_1396),
.B2(n_1471),
.Y(n_1516)
);

CKINVDCx6p67_ASAP7_75t_R g1517 ( 
.A(n_1348),
.Y(n_1517)
);

BUFx12f_ASAP7_75t_L g1518 ( 
.A(n_1361),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_1370),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1436),
.A2(n_1442),
.B1(n_1462),
.B2(n_1448),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1347),
.A2(n_1396),
.B1(n_1477),
.B2(n_1384),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1325),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1477),
.A2(n_1372),
.B1(n_1345),
.B2(n_1470),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1408),
.A2(n_1405),
.B1(n_1319),
.B2(n_1440),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1440),
.A2(n_1326),
.B1(n_1339),
.B2(n_1448),
.Y(n_1525)
);

INVx6_ASAP7_75t_L g1526 ( 
.A(n_1327),
.Y(n_1526)
);

INVx1_ASAP7_75t_SL g1527 ( 
.A(n_1331),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1404),
.Y(n_1528)
);

BUFx12f_ASAP7_75t_L g1529 ( 
.A(n_1340),
.Y(n_1529)
);

CKINVDCx10_ASAP7_75t_R g1530 ( 
.A(n_1319),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1431),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1442),
.A2(n_1339),
.B1(n_1426),
.B2(n_1435),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1313),
.A2(n_1317),
.B1(n_1466),
.B2(n_1465),
.Y(n_1533)
);

INVx6_ASAP7_75t_L g1534 ( 
.A(n_1330),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1450),
.A2(n_1452),
.B1(n_1463),
.B2(n_1460),
.Y(n_1535)
);

OAI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1422),
.A2(n_1435),
.B1(n_1344),
.B2(n_1442),
.Y(n_1536)
);

CKINVDCx11_ASAP7_75t_R g1537 ( 
.A(n_1330),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1446),
.A2(n_1438),
.B1(n_1422),
.B2(n_1443),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1430),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1405),
.B(n_1438),
.Y(n_1540)
);

BUFx4_ASAP7_75t_SL g1541 ( 
.A(n_1319),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1341),
.Y(n_1542)
);

BUFx10_ASAP7_75t_L g1543 ( 
.A(n_1415),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1446),
.A2(n_1376),
.B1(n_1432),
.B2(n_1443),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1351),
.A2(n_1439),
.B1(n_1344),
.B2(n_1320),
.Y(n_1545)
);

BUFx10_ASAP7_75t_L g1546 ( 
.A(n_1415),
.Y(n_1546)
);

NAND2x1p5_ASAP7_75t_L g1547 ( 
.A(n_1341),
.B(n_1388),
.Y(n_1547)
);

CKINVDCx16_ASAP7_75t_R g1548 ( 
.A(n_1351),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1474),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_SL g1550 ( 
.A1(n_1376),
.A2(n_1401),
.B1(n_1474),
.B2(n_1360),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1413),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1388),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1445),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1391),
.A2(n_1393),
.B1(n_1383),
.B2(n_1424),
.Y(n_1554)
);

BUFx4f_ASAP7_75t_SL g1555 ( 
.A(n_1412),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1371),
.A2(n_1380),
.B(n_1369),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_1363),
.Y(n_1557)
);

OAI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1401),
.A2(n_1350),
.B1(n_1363),
.B2(n_1445),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1432),
.A2(n_1444),
.B1(n_1469),
.B2(n_1335),
.Y(n_1559)
);

BUFx12f_ASAP7_75t_L g1560 ( 
.A(n_1412),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1444),
.A2(n_1447),
.B1(n_1350),
.B2(n_1355),
.Y(n_1561)
);

INVx6_ASAP7_75t_L g1562 ( 
.A(n_1447),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1378),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1434),
.Y(n_1564)
);

BUFx12f_ASAP7_75t_L g1565 ( 
.A(n_1412),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1418),
.B(n_1419),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1390),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1418),
.B(n_1419),
.Y(n_1568)
);

INVx6_ASAP7_75t_L g1569 ( 
.A(n_1437),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1378),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1478),
.A2(n_1349),
.B1(n_1324),
.B2(n_1334),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1390),
.A2(n_1337),
.B1(n_1368),
.B2(n_1375),
.Y(n_1572)
);

NAND4xp25_ASAP7_75t_SL g1573 ( 
.A(n_1352),
.B(n_1417),
.C(n_1378),
.D(n_1379),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1379),
.Y(n_1574)
);

OAI21xp33_ASAP7_75t_L g1575 ( 
.A1(n_1399),
.A2(n_1421),
.B(n_1343),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1417),
.B(n_1379),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1337),
.A2(n_1478),
.B1(n_1441),
.B2(n_1356),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1418),
.B(n_1419),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1417),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_SL g1580 ( 
.A1(n_1359),
.A2(n_1346),
.B1(n_1423),
.B2(n_1451),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1425),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1333),
.A2(n_1410),
.B1(n_1353),
.B2(n_1461),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1425),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1454),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1423),
.A2(n_1479),
.B1(n_1476),
.B2(n_1451),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1323),
.A2(n_1423),
.B1(n_1476),
.B2(n_1451),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1425),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1476),
.Y(n_1588)
);

BUFx4f_ASAP7_75t_L g1589 ( 
.A(n_1321),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1479),
.A2(n_1464),
.B1(n_1382),
.B2(n_1458),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1328),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1328),
.Y(n_1592)
);

CKINVDCx11_ASAP7_75t_R g1593 ( 
.A(n_1328),
.Y(n_1593)
);

BUFx2_ASAP7_75t_SL g1594 ( 
.A(n_1342),
.Y(n_1594)
);

INVx6_ASAP7_75t_L g1595 ( 
.A(n_1342),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1464),
.A2(n_1031),
.B1(n_1367),
.B2(n_625),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_1357),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1357),
.Y(n_1598)
);

CKINVDCx11_ASAP7_75t_R g1599 ( 
.A(n_1329),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1427),
.Y(n_1600)
);

CKINVDCx6p67_ASAP7_75t_R g1601 ( 
.A(n_1316),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1427),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_SL g1603 ( 
.A1(n_1464),
.A2(n_1031),
.B1(n_1367),
.B2(n_625),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1456),
.B(n_979),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1389),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1464),
.A2(n_1382),
.B1(n_1458),
.B2(n_1031),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1456),
.B(n_979),
.Y(n_1607)
);

CKINVDCx6p67_ASAP7_75t_R g1608 ( 
.A(n_1316),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1327),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1458),
.A2(n_1172),
.B(n_1464),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1357),
.Y(n_1611)
);

CKINVDCx11_ASAP7_75t_R g1612 ( 
.A(n_1329),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1327),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1427),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1357),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1342),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1357),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1427),
.Y(n_1618)
);

INVx6_ASAP7_75t_L g1619 ( 
.A(n_1342),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1325),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1464),
.A2(n_1382),
.B1(n_1458),
.B2(n_1031),
.Y(n_1621)
);

NAND2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1442),
.B(n_1068),
.Y(n_1622)
);

INVx4_ASAP7_75t_L g1623 ( 
.A(n_1342),
.Y(n_1623)
);

OA21x2_ASAP7_75t_L g1624 ( 
.A1(n_1324),
.A2(n_1459),
.B(n_1455),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1464),
.A2(n_1458),
.B1(n_1374),
.B2(n_804),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1427),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_SL g1627 ( 
.A1(n_1464),
.A2(n_1031),
.B1(n_1367),
.B2(n_625),
.Y(n_1627)
);

BUFx4f_ASAP7_75t_SL g1628 ( 
.A(n_1389),
.Y(n_1628)
);

CKINVDCx11_ASAP7_75t_R g1629 ( 
.A(n_1329),
.Y(n_1629)
);

OAI22x1_ASAP7_75t_L g1630 ( 
.A1(n_1458),
.A2(n_1374),
.B1(n_690),
.B2(n_1407),
.Y(n_1630)
);

BUFx4f_ASAP7_75t_SL g1631 ( 
.A(n_1389),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1458),
.A2(n_1464),
.B1(n_1172),
.B2(n_804),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1427),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_SL g1634 ( 
.A1(n_1464),
.A2(n_1031),
.B1(n_1367),
.B2(n_625),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1427),
.Y(n_1635)
);

CKINVDCx6p67_ASAP7_75t_R g1636 ( 
.A(n_1316),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1374),
.A2(n_804),
.B1(n_1031),
.B2(n_1080),
.Y(n_1637)
);

CKINVDCx20_ASAP7_75t_R g1638 ( 
.A(n_1357),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1315),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1464),
.A2(n_1382),
.B1(n_1458),
.B2(n_1031),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1458),
.A2(n_1464),
.B1(n_1172),
.B2(n_804),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1389),
.Y(n_1642)
);

BUFx6f_ASAP7_75t_SL g1643 ( 
.A(n_1342),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_SL g1644 ( 
.A1(n_1464),
.A2(n_1031),
.B1(n_1367),
.B2(n_625),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1427),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1458),
.A2(n_1464),
.B1(n_1172),
.B2(n_804),
.Y(n_1646)
);

OAI22x1_ASAP7_75t_L g1647 ( 
.A1(n_1458),
.A2(n_1374),
.B1(n_690),
.B2(n_1407),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_L g1648 ( 
.A(n_1327),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1357),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1592),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1498),
.B(n_1604),
.Y(n_1651)
);

OA21x2_ASAP7_75t_L g1652 ( 
.A1(n_1544),
.A2(n_1579),
.B(n_1570),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1563),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1606),
.A2(n_1640),
.B1(n_1621),
.B2(n_1634),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1576),
.B(n_1564),
.Y(n_1655)
);

OA21x2_ASAP7_75t_L g1656 ( 
.A1(n_1574),
.A2(n_1568),
.B(n_1566),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1578),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1499),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1559),
.A2(n_1582),
.B(n_1571),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1561),
.A2(n_1577),
.B(n_1587),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1637),
.A2(n_1641),
.B1(n_1632),
.B2(n_1646),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1610),
.B(n_1588),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1549),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1591),
.B(n_1624),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1562),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1624),
.B(n_1548),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1549),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1583),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1498),
.B(n_1607),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1560),
.Y(n_1670)
);

AOI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1630),
.A2(n_1647),
.B(n_1532),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1565),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1555),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1555),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1573),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1484),
.A2(n_1606),
.B1(n_1640),
.B2(n_1621),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1581),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1496),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1562),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1562),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1499),
.B(n_1553),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1585),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1499),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1497),
.B(n_1495),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1585),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1596),
.A2(n_1603),
.B1(n_1644),
.B2(n_1634),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1593),
.Y(n_1687)
);

OAI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1488),
.A2(n_1514),
.B1(n_1499),
.B2(n_1507),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1527),
.Y(n_1689)
);

NAND3xp33_ASAP7_75t_SL g1690 ( 
.A(n_1625),
.B(n_1484),
.C(n_1596),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1558),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1558),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1569),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1569),
.Y(n_1694)
);

BUFx12f_ASAP7_75t_L g1695 ( 
.A(n_1504),
.Y(n_1695)
);

AO21x1_ASAP7_75t_SL g1696 ( 
.A1(n_1590),
.A2(n_1506),
.B(n_1495),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1584),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1520),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1528),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1586),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_L g1701 ( 
.A(n_1603),
.B(n_1644),
.C(n_1627),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1586),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1481),
.B(n_1483),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1536),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1531),
.B(n_1509),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1497),
.B(n_1600),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1536),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1602),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1614),
.B(n_1618),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1626),
.Y(n_1710)
);

OAI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1627),
.A2(n_1506),
.B(n_1505),
.Y(n_1711)
);

AO21x1_ASAP7_75t_SL g1712 ( 
.A1(n_1590),
.A2(n_1554),
.B(n_1538),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1633),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1635),
.Y(n_1714)
);

INVx2_ASAP7_75t_SL g1715 ( 
.A(n_1496),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1645),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1487),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1491),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1538),
.Y(n_1719)
);

INVxp67_ASAP7_75t_L g1720 ( 
.A(n_1620),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1550),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1524),
.A2(n_1486),
.B1(n_1492),
.B2(n_1501),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1550),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1545),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1589),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1551),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1567),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1496),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1543),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1589),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1543),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1539),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1546),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1494),
.B(n_1505),
.Y(n_1734)
);

AO21x2_ASAP7_75t_L g1735 ( 
.A1(n_1575),
.A2(n_1507),
.B(n_1480),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1546),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1580),
.Y(n_1737)
);

OA21x2_ASAP7_75t_L g1738 ( 
.A1(n_1554),
.A2(n_1556),
.B(n_1525),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1580),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1525),
.B(n_1512),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1511),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1480),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1547),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1533),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1533),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1535),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1535),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1572),
.Y(n_1748)
);

NAND2x1p5_ASAP7_75t_L g1749 ( 
.A(n_1540),
.B(n_1609),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1516),
.B(n_1513),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1572),
.Y(n_1751)
);

AO21x2_ASAP7_75t_L g1752 ( 
.A1(n_1501),
.A2(n_1622),
.B(n_1557),
.Y(n_1752)
);

OAI21x1_ASAP7_75t_L g1753 ( 
.A1(n_1521),
.A2(n_1547),
.B(n_1523),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1515),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1639),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1541),
.Y(n_1756)
);

AOI31xp33_ASAP7_75t_L g1757 ( 
.A1(n_1611),
.A2(n_1615),
.A3(n_1617),
.B(n_1616),
.Y(n_1757)
);

OA21x2_ASAP7_75t_L g1758 ( 
.A1(n_1542),
.A2(n_1552),
.B(n_1541),
.Y(n_1758)
);

INVx4_ASAP7_75t_L g1759 ( 
.A(n_1613),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1485),
.B(n_1609),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1613),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1648),
.A2(n_1485),
.B(n_1508),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1648),
.Y(n_1763)
);

OAI21x1_ASAP7_75t_L g1764 ( 
.A1(n_1508),
.A2(n_1530),
.B(n_1643),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1648),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1526),
.Y(n_1766)
);

CKINVDCx20_ASAP7_75t_R g1767 ( 
.A(n_1490),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1623),
.B(n_1594),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1526),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1510),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1534),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1500),
.B(n_1623),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1510),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1510),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1595),
.Y(n_1775)
);

OAI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1628),
.A2(n_1631),
.B1(n_1608),
.B2(n_1601),
.Y(n_1776)
);

BUFx3_ASAP7_75t_L g1777 ( 
.A(n_1595),
.Y(n_1777)
);

INVx6_ASAP7_75t_L g1778 ( 
.A(n_1595),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1619),
.Y(n_1779)
);

NAND2x1p5_ASAP7_75t_L g1780 ( 
.A(n_1489),
.B(n_1605),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1619),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1642),
.B(n_1522),
.Y(n_1782)
);

INVx2_ASAP7_75t_SL g1783 ( 
.A(n_1619),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1537),
.B(n_1519),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1643),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1529),
.Y(n_1786)
);

O2A1O1Ixp33_ASAP7_75t_L g1787 ( 
.A1(n_1690),
.A2(n_1649),
.B(n_1638),
.C(n_1598),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1676),
.A2(n_1636),
.B1(n_1517),
.B2(n_1628),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1655),
.B(n_1502),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1655),
.B(n_1518),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1666),
.B(n_1482),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1666),
.B(n_1599),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1670),
.B(n_1597),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1651),
.B(n_1482),
.Y(n_1794)
);

AO32x2_ASAP7_75t_L g1795 ( 
.A1(n_1722),
.A2(n_1631),
.A3(n_1612),
.B1(n_1629),
.B2(n_1493),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1767),
.Y(n_1796)
);

AOI21x1_ASAP7_75t_L g1797 ( 
.A1(n_1729),
.A2(n_1503),
.B(n_1733),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1669),
.B(n_1716),
.Y(n_1798)
);

O2A1O1Ixp33_ASAP7_75t_SL g1799 ( 
.A1(n_1688),
.A2(n_1701),
.B(n_1711),
.C(n_1693),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1695),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1706),
.B(n_1687),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1670),
.B(n_1673),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1673),
.B(n_1674),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1661),
.B(n_1701),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1734),
.B(n_1708),
.Y(n_1805)
);

INVxp67_ASAP7_75t_SL g1806 ( 
.A(n_1663),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1654),
.A2(n_1686),
.B1(n_1684),
.B2(n_1741),
.Y(n_1807)
);

NOR2x1_ASAP7_75t_L g1808 ( 
.A(n_1729),
.B(n_1733),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1684),
.A2(n_1741),
.B1(n_1740),
.B2(n_1750),
.Y(n_1809)
);

OA21x2_ASAP7_75t_L g1810 ( 
.A1(n_1659),
.A2(n_1660),
.B(n_1748),
.Y(n_1810)
);

BUFx3_ASAP7_75t_L g1811 ( 
.A(n_1782),
.Y(n_1811)
);

BUFx3_ASAP7_75t_L g1812 ( 
.A(n_1782),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1708),
.B(n_1710),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1662),
.B(n_1664),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1662),
.B(n_1664),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1752),
.B(n_1750),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1782),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1736),
.B(n_1731),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1752),
.B(n_1698),
.Y(n_1819)
);

AO21x1_ASAP7_75t_L g1820 ( 
.A1(n_1675),
.A2(n_1694),
.B(n_1693),
.Y(n_1820)
);

NOR2x1p5_ASAP7_75t_L g1821 ( 
.A(n_1695),
.B(n_1725),
.Y(n_1821)
);

AND2x6_ASAP7_75t_L g1822 ( 
.A(n_1725),
.B(n_1694),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1754),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1727),
.B(n_1704),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1681),
.B(n_1672),
.Y(n_1825)
);

NOR2x1_ASAP7_75t_SL g1826 ( 
.A(n_1712),
.B(n_1696),
.Y(n_1826)
);

A2O1A1Ixp33_ASAP7_75t_L g1827 ( 
.A1(n_1724),
.A2(n_1740),
.B(n_1698),
.C(n_1742),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1754),
.Y(n_1828)
);

AO32x2_ASAP7_75t_L g1829 ( 
.A1(n_1759),
.A2(n_1682),
.A3(n_1685),
.B1(n_1783),
.B2(n_1739),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1681),
.B(n_1672),
.Y(n_1830)
);

NAND2x1p5_ASAP7_75t_L g1831 ( 
.A(n_1758),
.B(n_1658),
.Y(n_1831)
);

OA21x2_ASAP7_75t_L g1832 ( 
.A1(n_1659),
.A2(n_1660),
.B(n_1751),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1713),
.B(n_1714),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1749),
.B(n_1760),
.Y(n_1834)
);

AO32x2_ASAP7_75t_L g1835 ( 
.A1(n_1759),
.A2(n_1682),
.A3(n_1685),
.B1(n_1783),
.B2(n_1737),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1742),
.A2(n_1724),
.B1(n_1719),
.B2(n_1756),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1727),
.B(n_1704),
.Y(n_1837)
);

O2A1O1Ixp33_ASAP7_75t_L g1838 ( 
.A1(n_1689),
.A2(n_1699),
.B(n_1707),
.C(n_1732),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1761),
.B(n_1744),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1671),
.A2(n_1738),
.B(n_1719),
.Y(n_1840)
);

A2O1A1Ixp33_ASAP7_75t_L g1841 ( 
.A1(n_1696),
.A2(n_1753),
.B(n_1691),
.C(n_1692),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1744),
.A2(n_1747),
.B1(n_1746),
.B2(n_1745),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1745),
.B(n_1746),
.Y(n_1843)
);

CKINVDCx20_ASAP7_75t_R g1844 ( 
.A(n_1784),
.Y(n_1844)
);

AOI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1756),
.A2(n_1705),
.B1(n_1735),
.B2(n_1776),
.Y(n_1845)
);

OAI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1738),
.A2(n_1753),
.B(n_1748),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1747),
.B(n_1763),
.Y(n_1847)
);

NOR2x1_ASAP7_75t_SL g1848 ( 
.A(n_1658),
.B(n_1683),
.Y(n_1848)
);

OAI211xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1720),
.A2(n_1751),
.B(n_1785),
.C(n_1755),
.Y(n_1849)
);

OAI211xp5_ASAP7_75t_L g1850 ( 
.A1(n_1738),
.A2(n_1721),
.B(n_1723),
.C(n_1703),
.Y(n_1850)
);

A2O1A1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1764),
.A2(n_1730),
.B(n_1725),
.C(n_1785),
.Y(n_1851)
);

OA21x2_ASAP7_75t_L g1852 ( 
.A1(n_1653),
.A2(n_1667),
.B(n_1663),
.Y(n_1852)
);

OAI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1738),
.A2(n_1680),
.B(n_1679),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1765),
.B(n_1773),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1735),
.A2(n_1680),
.B(n_1679),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1679),
.A2(n_1697),
.B(n_1665),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1653),
.Y(n_1857)
);

A2O1A1Ixp33_ASAP7_75t_L g1858 ( 
.A1(n_1764),
.A2(n_1725),
.B(n_1683),
.C(n_1768),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1773),
.B(n_1775),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1735),
.A2(n_1782),
.B1(n_1786),
.B2(n_1758),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1773),
.B(n_1781),
.Y(n_1861)
);

A2O1A1Ixp33_ASAP7_75t_L g1862 ( 
.A1(n_1683),
.A2(n_1714),
.B(n_1709),
.C(n_1665),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1770),
.Y(n_1863)
);

AO32x2_ASAP7_75t_L g1864 ( 
.A1(n_1759),
.A2(n_1700),
.A3(n_1702),
.B1(n_1656),
.B2(n_1715),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1657),
.B(n_1718),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1823),
.Y(n_1866)
);

INVxp67_ASAP7_75t_SL g1867 ( 
.A(n_1838),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1852),
.Y(n_1868)
);

INVx1_ASAP7_75t_SL g1869 ( 
.A(n_1823),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1801),
.B(n_1667),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1852),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1857),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1802),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1816),
.B(n_1700),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1806),
.Y(n_1875)
);

AOI221xp5_ASAP7_75t_L g1876 ( 
.A1(n_1804),
.A2(n_1717),
.B1(n_1718),
.B2(n_1668),
.C(n_1757),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1814),
.B(n_1815),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1819),
.B(n_1668),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1804),
.A2(n_1758),
.B1(n_1665),
.B2(n_1772),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1798),
.B(n_1656),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1794),
.A2(n_1665),
.B1(n_1775),
.B2(n_1781),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1806),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1828),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1798),
.B(n_1656),
.Y(n_1884)
);

NOR2x1p5_ASAP7_75t_L g1885 ( 
.A(n_1797),
.B(n_1781),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1794),
.A2(n_1775),
.B1(n_1743),
.B2(n_1779),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1846),
.B(n_1652),
.Y(n_1887)
);

INVxp67_ASAP7_75t_SL g1888 ( 
.A(n_1838),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1846),
.B(n_1652),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1831),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1810),
.B(n_1652),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1848),
.B(n_1677),
.Y(n_1892)
);

BUFx2_ASAP7_75t_L g1893 ( 
.A(n_1831),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1864),
.B(n_1652),
.Y(n_1894)
);

INVxp67_ASAP7_75t_SL g1895 ( 
.A(n_1865),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_1864),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1828),
.Y(n_1897)
);

BUFx2_ASAP7_75t_L g1898 ( 
.A(n_1864),
.Y(n_1898)
);

HB1xp67_ASAP7_75t_L g1899 ( 
.A(n_1839),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_1808),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1845),
.A2(n_1743),
.B1(n_1779),
.B2(n_1770),
.Y(n_1901)
);

OAI21xp33_ASAP7_75t_L g1902 ( 
.A1(n_1807),
.A2(n_1827),
.B(n_1850),
.Y(n_1902)
);

INVx4_ASAP7_75t_L g1903 ( 
.A(n_1822),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1859),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1805),
.B(n_1843),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1813),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1805),
.B(n_1697),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1853),
.B(n_1650),
.Y(n_1908)
);

AOI22xp33_ASAP7_75t_L g1909 ( 
.A1(n_1849),
.A2(n_1774),
.B1(n_1777),
.B2(n_1770),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1849),
.A2(n_1774),
.B1(n_1777),
.B2(n_1778),
.Y(n_1910)
);

NOR2xp67_ASAP7_75t_L g1911 ( 
.A(n_1855),
.B(n_1726),
.Y(n_1911)
);

HB1xp67_ASAP7_75t_L g1912 ( 
.A(n_1861),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1810),
.B(n_1650),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1832),
.B(n_1650),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1847),
.Y(n_1915)
);

INVxp67_ASAP7_75t_L g1916 ( 
.A(n_1818),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1813),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1903),
.B(n_1825),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1877),
.B(n_1860),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1868),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1914),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1868),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1871),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1871),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1872),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1916),
.B(n_1841),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1902),
.A2(n_1812),
.B1(n_1817),
.B2(n_1811),
.Y(n_1927)
);

OAI321xp33_ASAP7_75t_L g1928 ( 
.A1(n_1902),
.A2(n_1850),
.A3(n_1827),
.B1(n_1840),
.B2(n_1836),
.C(n_1842),
.Y(n_1928)
);

HB1xp67_ASAP7_75t_L g1929 ( 
.A(n_1866),
.Y(n_1929)
);

AOI222xp33_ASAP7_75t_L g1930 ( 
.A1(n_1876),
.A2(n_1826),
.B1(n_1867),
.B2(n_1888),
.C1(n_1840),
.C2(n_1799),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1916),
.B(n_1841),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1876),
.A2(n_1809),
.B1(n_1788),
.B2(n_1787),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1877),
.B(n_1832),
.Y(n_1933)
);

AOI31xp33_ASAP7_75t_L g1934 ( 
.A1(n_1879),
.A2(n_1799),
.A3(n_1820),
.B(n_1792),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1914),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1905),
.B(n_1791),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1872),
.Y(n_1937)
);

OAI321xp33_ASAP7_75t_L g1938 ( 
.A1(n_1879),
.A2(n_1842),
.A3(n_1889),
.B1(n_1787),
.B2(n_1901),
.C(n_1887),
.Y(n_1938)
);

INVx1_ASAP7_75t_SL g1939 ( 
.A(n_1869),
.Y(n_1939)
);

INVxp67_ASAP7_75t_SL g1940 ( 
.A(n_1900),
.Y(n_1940)
);

BUFx3_ASAP7_75t_L g1941 ( 
.A(n_1892),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1904),
.B(n_1829),
.Y(n_1942)
);

OR2x6_ASAP7_75t_L g1943 ( 
.A(n_1903),
.B(n_1862),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1912),
.B(n_1829),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1895),
.B(n_1824),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1874),
.B(n_1829),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1875),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1874),
.B(n_1835),
.Y(n_1948)
);

OAI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1900),
.A2(n_1862),
.B(n_1858),
.Y(n_1949)
);

AOI221xp5_ASAP7_75t_L g1950 ( 
.A1(n_1896),
.A2(n_1818),
.B1(n_1851),
.B2(n_1856),
.C(n_1802),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1913),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1915),
.B(n_1835),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_SL g1953 ( 
.A1(n_1896),
.A2(n_1795),
.B1(n_1800),
.B2(n_1844),
.Y(n_1953)
);

NAND3xp33_ASAP7_75t_L g1954 ( 
.A(n_1889),
.B(n_1856),
.C(n_1837),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1886),
.A2(n_1821),
.B1(n_1881),
.B2(n_1789),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1883),
.Y(n_1956)
);

BUFx3_ASAP7_75t_L g1957 ( 
.A(n_1892),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1913),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1870),
.B(n_1835),
.Y(n_1959)
);

OAI211xp5_ASAP7_75t_SL g1960 ( 
.A1(n_1880),
.A2(n_1771),
.B(n_1769),
.C(n_1766),
.Y(n_1960)
);

OAI222xp33_ASAP7_75t_L g1961 ( 
.A1(n_1869),
.A2(n_1830),
.B1(n_1803),
.B2(n_1790),
.C1(n_1834),
.C2(n_1780),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1891),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1903),
.B(n_1803),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1897),
.B(n_1854),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1898),
.A2(n_1863),
.B1(n_1865),
.B2(n_1833),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1880),
.B(n_1833),
.Y(n_1966)
);

INVx3_ASAP7_75t_L g1967 ( 
.A(n_1892),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1882),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_1873),
.Y(n_1969)
);

AND4x1_ASAP7_75t_L g1970 ( 
.A(n_1930),
.B(n_1910),
.C(n_1909),
.D(n_1795),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1920),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1951),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1933),
.B(n_1898),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1933),
.B(n_1894),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1967),
.B(n_1894),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_R g1976 ( 
.A(n_1927),
.B(n_1796),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1920),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1951),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1966),
.B(n_1895),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1951),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1922),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1967),
.B(n_1958),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1958),
.Y(n_1983)
);

BUFx2_ASAP7_75t_L g1984 ( 
.A(n_1943),
.Y(n_1984)
);

INVx2_ASAP7_75t_SL g1985 ( 
.A(n_1941),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1966),
.B(n_1884),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1922),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1967),
.B(n_1887),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1940),
.B(n_1884),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1958),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1946),
.B(n_1906),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1946),
.B(n_1906),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1923),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1967),
.B(n_1890),
.Y(n_1994)
);

INVxp67_ASAP7_75t_L g1995 ( 
.A(n_1926),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1952),
.B(n_1890),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1952),
.B(n_1893),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1923),
.Y(n_1998)
);

HB1xp67_ASAP7_75t_L g1999 ( 
.A(n_1924),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1924),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1942),
.B(n_1893),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1947),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1948),
.B(n_1917),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1925),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1925),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1948),
.B(n_1945),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1937),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1945),
.B(n_1917),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1941),
.B(n_1911),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1962),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1931),
.B(n_1873),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1962),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1962),
.Y(n_2013)
);

OAI21x1_ASAP7_75t_L g2014 ( 
.A1(n_1921),
.A2(n_1891),
.B(n_1908),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1942),
.B(n_1908),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1921),
.B(n_1907),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1944),
.B(n_1899),
.Y(n_2017)
);

INVx6_ASAP7_75t_L g2018 ( 
.A(n_1943),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1919),
.B(n_1878),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1947),
.Y(n_2020)
);

INVx1_ASAP7_75t_SL g2021 ( 
.A(n_1939),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1999),
.Y(n_2022)
);

INVx1_ASAP7_75t_SL g2023 ( 
.A(n_2021),
.Y(n_2023)
);

OAI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_1984),
.A2(n_1934),
.B1(n_1928),
.B2(n_1938),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_2006),
.B(n_1954),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1999),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2002),
.Y(n_2027)
);

AND3x1_ASAP7_75t_L g2028 ( 
.A(n_2011),
.B(n_1950),
.C(n_1955),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2002),
.Y(n_2029)
);

OAI32xp33_ASAP7_75t_L g2030 ( 
.A1(n_1995),
.A2(n_1932),
.A3(n_1949),
.B1(n_1965),
.B2(n_1939),
.Y(n_2030)
);

NAND3xp33_ASAP7_75t_SL g2031 ( 
.A(n_1970),
.B(n_1930),
.C(n_1949),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1984),
.B(n_1941),
.Y(n_2032)
);

BUFx2_ASAP7_75t_L g2033 ( 
.A(n_1984),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2020),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_2021),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2020),
.Y(n_2036)
);

INVxp67_ASAP7_75t_L g2037 ( 
.A(n_2011),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1985),
.B(n_1957),
.Y(n_2038)
);

NAND2x1_ASAP7_75t_L g2039 ( 
.A(n_2018),
.B(n_1943),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_1995),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1977),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_2019),
.B(n_1919),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1977),
.Y(n_2043)
);

NOR2x1_ASAP7_75t_L g2044 ( 
.A(n_1989),
.B(n_1934),
.Y(n_2044)
);

INVx1_ASAP7_75t_SL g2045 ( 
.A(n_1976),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1970),
.B(n_1928),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1996),
.B(n_1957),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1977),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1996),
.B(n_1957),
.Y(n_2049)
);

NOR2x1p5_ASAP7_75t_SL g2050 ( 
.A(n_2010),
.B(n_1921),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1981),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2019),
.B(n_1929),
.Y(n_2052)
);

NAND2x1p5_ASAP7_75t_L g2053 ( 
.A(n_1985),
.B(n_1963),
.Y(n_2053)
);

NAND2xp33_ASAP7_75t_L g2054 ( 
.A(n_1976),
.B(n_1953),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1981),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1996),
.B(n_1959),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1981),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1987),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_1985),
.B(n_1963),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_2018),
.A2(n_1953),
.B1(n_1932),
.B2(n_1955),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_2019),
.Y(n_2061)
);

NAND3xp33_ASAP7_75t_L g2062 ( 
.A(n_1989),
.B(n_1954),
.C(n_1965),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1987),
.Y(n_2063)
);

HB1xp67_ASAP7_75t_L g2064 ( 
.A(n_2008),
.Y(n_2064)
);

BUFx2_ASAP7_75t_L g2065 ( 
.A(n_2018),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1982),
.Y(n_2066)
);

AOI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_2018),
.A2(n_1943),
.B1(n_1885),
.B2(n_1963),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2008),
.B(n_1956),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1987),
.Y(n_2069)
);

OAI33xp33_ASAP7_75t_L g2070 ( 
.A1(n_1979),
.A2(n_1971),
.A3(n_1993),
.B1(n_1998),
.B2(n_2000),
.B3(n_2006),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1979),
.B(n_1936),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_1986),
.B(n_1935),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2047),
.B(n_1973),
.Y(n_2073)
);

OAI31xp33_ASAP7_75t_L g2074 ( 
.A1(n_2024),
.A2(n_2046),
.A3(n_2060),
.B(n_2062),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2040),
.B(n_2015),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2035),
.Y(n_2076)
);

AOI31xp33_ASAP7_75t_L g2077 ( 
.A1(n_2046),
.A2(n_1780),
.A3(n_1793),
.B(n_1938),
.Y(n_2077)
);

NAND4xp25_ASAP7_75t_SL g2078 ( 
.A(n_2044),
.B(n_1973),
.C(n_1988),
.D(n_1997),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2037),
.B(n_2015),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2041),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2047),
.B(n_1973),
.Y(n_2081)
);

AND2x2_ASAP7_75t_SL g2082 ( 
.A(n_2054),
.B(n_1793),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2042),
.B(n_1986),
.Y(n_2083)
);

INVxp67_ASAP7_75t_L g2084 ( 
.A(n_2033),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2023),
.B(n_2015),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_2061),
.B(n_2025),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2025),
.B(n_2016),
.Y(n_2087)
);

AOI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_2031),
.A2(n_2018),
.B1(n_1943),
.B2(n_1885),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2071),
.B(n_2017),
.Y(n_2089)
);

HB1xp67_ASAP7_75t_L g2090 ( 
.A(n_2033),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2066),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2043),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2048),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2051),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_2045),
.B(n_1780),
.Y(n_2095)
);

BUFx2_ASAP7_75t_L g2096 ( 
.A(n_2053),
.Y(n_2096)
);

INVxp67_ASAP7_75t_L g2097 ( 
.A(n_2028),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2049),
.B(n_1997),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2049),
.B(n_1997),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2064),
.B(n_2017),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2055),
.Y(n_2101)
);

INVxp67_ASAP7_75t_L g2102 ( 
.A(n_2054),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2057),
.Y(n_2103)
);

OAI21xp5_ASAP7_75t_SL g2104 ( 
.A1(n_2067),
.A2(n_1961),
.B(n_1960),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2052),
.B(n_2017),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2053),
.B(n_2001),
.Y(n_2106)
);

OR2x2_ASAP7_75t_L g2107 ( 
.A(n_2068),
.B(n_2016),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_2030),
.B(n_2018),
.Y(n_2108)
);

NAND4xp25_ASAP7_75t_L g2109 ( 
.A(n_2065),
.B(n_1988),
.C(n_2001),
.D(n_1975),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2032),
.B(n_2001),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2058),
.Y(n_2111)
);

AND2x4_ASAP7_75t_L g2112 ( 
.A(n_2059),
.B(n_2009),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2090),
.Y(n_2113)
);

OAI22xp33_ASAP7_75t_L g2114 ( 
.A1(n_2077),
.A2(n_2039),
.B1(n_2018),
.B2(n_2065),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2093),
.Y(n_2115)
);

OAI21xp33_ASAP7_75t_L g2116 ( 
.A1(n_2097),
.A2(n_2102),
.B(n_2078),
.Y(n_2116)
);

OAI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_2074),
.A2(n_2039),
.B(n_2032),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2093),
.Y(n_2118)
);

OAI22x1_ASAP7_75t_L g2119 ( 
.A1(n_2088),
.A2(n_2059),
.B1(n_2038),
.B2(n_2026),
.Y(n_2119)
);

NAND2xp33_ASAP7_75t_R g2120 ( 
.A(n_2108),
.B(n_2038),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2112),
.Y(n_2121)
);

OR2x2_ASAP7_75t_L g2122 ( 
.A(n_2085),
.B(n_2072),
.Y(n_2122)
);

INVx1_ASAP7_75t_SL g2123 ( 
.A(n_2082),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2076),
.B(n_2056),
.Y(n_2124)
);

NAND3xp33_ASAP7_75t_L g2125 ( 
.A(n_2084),
.B(n_2022),
.C(n_2063),
.Y(n_2125)
);

INVx1_ASAP7_75t_SL g2126 ( 
.A(n_2082),
.Y(n_2126)
);

OAI22xp33_ASAP7_75t_L g2127 ( 
.A1(n_2104),
.A2(n_1795),
.B1(n_2072),
.B2(n_2066),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2110),
.B(n_2056),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2098),
.B(n_2059),
.Y(n_2129)
);

NAND3xp33_ASAP7_75t_L g2130 ( 
.A(n_2086),
.B(n_2069),
.C(n_2029),
.Y(n_2130)
);

OR2x2_ASAP7_75t_L g2131 ( 
.A(n_2086),
.B(n_2027),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_2096),
.Y(n_2132)
);

OAI22xp33_ASAP7_75t_SL g2133 ( 
.A1(n_2096),
.A2(n_2038),
.B1(n_2036),
.B2(n_2034),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2110),
.B(n_1991),
.Y(n_2134)
);

A2O1A1Ixp33_ASAP7_75t_L g2135 ( 
.A1(n_2095),
.A2(n_2050),
.B(n_2014),
.C(n_2009),
.Y(n_2135)
);

OAI211xp5_ASAP7_75t_SL g2136 ( 
.A1(n_2079),
.A2(n_2075),
.B(n_2100),
.C(n_2083),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2112),
.Y(n_2137)
);

OAI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_2089),
.A2(n_2105),
.B1(n_2099),
.B2(n_2098),
.Y(n_2138)
);

OAI21xp33_ASAP7_75t_L g2139 ( 
.A1(n_2109),
.A2(n_2050),
.B(n_1988),
.Y(n_2139)
);

HB1xp67_ASAP7_75t_L g2140 ( 
.A(n_2087),
.Y(n_2140)
);

AOI221xp5_ASAP7_75t_L g2141 ( 
.A1(n_2080),
.A2(n_2070),
.B1(n_2111),
.B2(n_2094),
.C(n_2092),
.Y(n_2141)
);

OAI22xp5_ASAP7_75t_L g2142 ( 
.A1(n_2127),
.A2(n_2106),
.B1(n_2099),
.B2(n_2073),
.Y(n_2142)
);

AOI22xp5_ASAP7_75t_L g2143 ( 
.A1(n_2127),
.A2(n_2106),
.B1(n_2112),
.B2(n_2081),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2140),
.Y(n_2144)
);

OAI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_2117),
.A2(n_2087),
.B(n_2101),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2140),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2129),
.B(n_2123),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2116),
.B(n_2073),
.Y(n_2148)
);

OAI32xp33_ASAP7_75t_L g2149 ( 
.A1(n_2120),
.A2(n_2081),
.A3(n_2083),
.B1(n_2107),
.B2(n_2103),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2113),
.B(n_2107),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2115),
.Y(n_2151)
);

OAI21xp5_ASAP7_75t_L g2152 ( 
.A1(n_2125),
.A2(n_2101),
.B(n_2091),
.Y(n_2152)
);

AOI221xp5_ASAP7_75t_L g2153 ( 
.A1(n_2136),
.A2(n_2091),
.B1(n_2010),
.B2(n_2012),
.C(n_2013),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2132),
.B(n_2121),
.Y(n_2154)
);

INVx5_ASAP7_75t_L g2155 ( 
.A(n_2137),
.Y(n_2155)
);

O2A1O1Ixp33_ASAP7_75t_L g2156 ( 
.A1(n_2133),
.A2(n_2012),
.B(n_2010),
.C(n_2013),
.Y(n_2156)
);

OAI22xp5_ASAP7_75t_SL g2157 ( 
.A1(n_2126),
.A2(n_2009),
.B1(n_1994),
.B2(n_1963),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2118),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2119),
.B(n_1994),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2131),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2124),
.B(n_1991),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2130),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2122),
.Y(n_2163)
);

OAI22xp33_ASAP7_75t_L g2164 ( 
.A1(n_2120),
.A2(n_1992),
.B1(n_2003),
.B2(n_1969),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2128),
.Y(n_2165)
);

AOI22xp5_ASAP7_75t_SL g2166 ( 
.A1(n_2162),
.A2(n_2138),
.B1(n_2009),
.B2(n_2134),
.Y(n_2166)
);

OAI221xp5_ASAP7_75t_L g2167 ( 
.A1(n_2145),
.A2(n_2136),
.B1(n_2139),
.B2(n_2141),
.C(n_2135),
.Y(n_2167)
);

NAND5xp2_ASAP7_75t_L g2168 ( 
.A(n_2145),
.B(n_2114),
.C(n_1772),
.D(n_1975),
.E(n_1974),
.Y(n_2168)
);

AOI21xp33_ASAP7_75t_SL g2169 ( 
.A1(n_2149),
.A2(n_2114),
.B(n_2009),
.Y(n_2169)
);

XNOR2x1_ASAP7_75t_L g2170 ( 
.A(n_2147),
.B(n_1918),
.Y(n_2170)
);

OAI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_2143),
.A2(n_2142),
.B1(n_2148),
.B2(n_2146),
.Y(n_2171)
);

XNOR2xp5_ASAP7_75t_L g2172 ( 
.A(n_2165),
.B(n_1918),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_2164),
.B(n_2009),
.Y(n_2173)
);

AOI221xp5_ASAP7_75t_L g2174 ( 
.A1(n_2152),
.A2(n_2010),
.B1(n_2012),
.B2(n_2013),
.C(n_1993),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2144),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2160),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2155),
.B(n_1974),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2150),
.Y(n_2178)
);

A2O1A1Ixp33_ASAP7_75t_L g2179 ( 
.A1(n_2156),
.A2(n_2014),
.B(n_1994),
.C(n_1974),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2155),
.B(n_1992),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2171),
.B(n_2155),
.Y(n_2181)
);

INVx1_ASAP7_75t_SL g2182 ( 
.A(n_2166),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2175),
.Y(n_2183)
);

INVx1_ASAP7_75t_SL g2184 ( 
.A(n_2170),
.Y(n_2184)
);

NOR3xp33_ASAP7_75t_L g2185 ( 
.A(n_2167),
.B(n_2154),
.C(n_2163),
.Y(n_2185)
);

NOR2x1_ASAP7_75t_L g2186 ( 
.A(n_2176),
.B(n_2151),
.Y(n_2186)
);

HB1xp67_ASAP7_75t_L g2187 ( 
.A(n_2177),
.Y(n_2187)
);

INVx2_ASAP7_75t_SL g2188 ( 
.A(n_2172),
.Y(n_2188)
);

NAND4xp25_ASAP7_75t_SL g2189 ( 
.A(n_2169),
.B(n_2159),
.C(n_2152),
.D(n_2161),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_L g2190 ( 
.A(n_2178),
.B(n_2158),
.Y(n_2190)
);

OAI211xp5_ASAP7_75t_SL g2191 ( 
.A1(n_2171),
.A2(n_2179),
.B(n_2173),
.C(n_2174),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2180),
.B(n_2155),
.Y(n_2192)
);

AOI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_2189),
.A2(n_2157),
.B1(n_2153),
.B2(n_2168),
.Y(n_2193)
);

AOI221xp5_ASAP7_75t_L g2194 ( 
.A1(n_2191),
.A2(n_2013),
.B1(n_2012),
.B2(n_1994),
.C(n_1993),
.Y(n_2194)
);

OR2x2_ASAP7_75t_L g2195 ( 
.A(n_2187),
.B(n_2003),
.Y(n_2195)
);

INVxp33_ASAP7_75t_SL g2196 ( 
.A(n_2181),
.Y(n_2196)
);

AOI221xp5_ASAP7_75t_L g2197 ( 
.A1(n_2191),
.A2(n_1994),
.B1(n_2000),
.B2(n_1998),
.C(n_1971),
.Y(n_2197)
);

O2A1O1Ixp33_ASAP7_75t_L g2198 ( 
.A1(n_2182),
.A2(n_1983),
.B(n_1972),
.C(n_1980),
.Y(n_2198)
);

OAI221xp5_ASAP7_75t_SL g2199 ( 
.A1(n_2185),
.A2(n_2016),
.B1(n_1975),
.B2(n_1982),
.C(n_1978),
.Y(n_2199)
);

OAI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_2196),
.A2(n_2184),
.B(n_2186),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2195),
.B(n_2192),
.Y(n_2201)
);

BUFx6f_ASAP7_75t_L g2202 ( 
.A(n_2199),
.Y(n_2202)
);

OAI211xp5_ASAP7_75t_SL g2203 ( 
.A1(n_2193),
.A2(n_2188),
.B(n_2183),
.C(n_2190),
.Y(n_2203)
);

NAND4xp25_ASAP7_75t_SL g2204 ( 
.A(n_2197),
.B(n_1982),
.C(n_1972),
.D(n_1978),
.Y(n_2204)
);

OAI211xp5_ASAP7_75t_SL g2205 ( 
.A1(n_2194),
.A2(n_1964),
.B(n_2000),
.C(n_1998),
.Y(n_2205)
);

AOI221xp5_ASAP7_75t_L g2206 ( 
.A1(n_2198),
.A2(n_1994),
.B1(n_2005),
.B2(n_2007),
.C(n_1972),
.Y(n_2206)
);

NOR2x1_ASAP7_75t_L g2207 ( 
.A(n_2200),
.B(n_1774),
.Y(n_2207)
);

NAND4xp75_ASAP7_75t_L g2208 ( 
.A(n_2206),
.B(n_1728),
.C(n_1678),
.D(n_1715),
.Y(n_2208)
);

NAND2x1p5_ASAP7_75t_SL g2209 ( 
.A(n_2203),
.B(n_1678),
.Y(n_2209)
);

NAND2xp33_ASAP7_75t_L g2210 ( 
.A(n_2201),
.B(n_2004),
.Y(n_2210)
);

INVx2_ASAP7_75t_SL g2211 ( 
.A(n_2202),
.Y(n_2211)
);

NOR3xp33_ASAP7_75t_L g2212 ( 
.A(n_2211),
.B(n_2204),
.C(n_2205),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2207),
.B(n_1972),
.Y(n_2213)
);

OAI211xp5_ASAP7_75t_SL g2214 ( 
.A1(n_2210),
.A2(n_1728),
.B(n_1766),
.C(n_1771),
.Y(n_2214)
);

AOI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_2212),
.A2(n_2208),
.B1(n_2209),
.B2(n_1778),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2215),
.Y(n_2216)
);

NAND3xp33_ASAP7_75t_SL g2217 ( 
.A(n_2216),
.B(n_2213),
.C(n_2214),
.Y(n_2217)
);

AOI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_2216),
.A2(n_1983),
.B1(n_1978),
.B2(n_1980),
.Y(n_2218)
);

BUFx2_ASAP7_75t_L g2219 ( 
.A(n_2218),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2217),
.Y(n_2220)
);

AOI221xp5_ASAP7_75t_L g2221 ( 
.A1(n_2220),
.A2(n_2004),
.B1(n_1980),
.B2(n_1990),
.C(n_1983),
.Y(n_2221)
);

HB1xp67_ASAP7_75t_L g2222 ( 
.A(n_2219),
.Y(n_2222)
);

AOI21xp5_ASAP7_75t_L g2223 ( 
.A1(n_2222),
.A2(n_2221),
.B(n_1978),
.Y(n_2223)
);

AOI21xp5_ASAP7_75t_L g2224 ( 
.A1(n_2223),
.A2(n_1980),
.B(n_1990),
.Y(n_2224)
);

OAI22xp33_ASAP7_75t_L g2225 ( 
.A1(n_2224),
.A2(n_1990),
.B1(n_1983),
.B2(n_2005),
.Y(n_2225)
);

AOI221xp5_ASAP7_75t_L g2226 ( 
.A1(n_2225),
.A2(n_2007),
.B1(n_2005),
.B2(n_1990),
.C(n_1968),
.Y(n_2226)
);

AOI211xp5_ASAP7_75t_L g2227 ( 
.A1(n_2226),
.A2(n_1777),
.B(n_1762),
.C(n_1769),
.Y(n_2227)
);


endmodule