module fake_jpeg_27464_n_199 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_SL g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_16),
.B(n_0),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_23),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_29),
.C(n_18),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_60),
.B(n_42),
.C(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_52),
.Y(n_74)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_27),
.B1(n_21),
.B2(n_26),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_43),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_27),
.B1(n_21),
.B2(n_28),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_61),
.B1(n_41),
.B2(n_24),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_27),
.B1(n_19),
.B2(n_22),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_28),
.B1(n_30),
.B2(n_22),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_41),
.B1(n_24),
.B2(n_19),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_48),
.B1(n_51),
.B2(n_30),
.Y(n_92)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_51),
.B1(n_42),
.B2(n_35),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_73),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_63),
.B1(n_48),
.B2(n_55),
.Y(n_87)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_33),
.A3(n_32),
.B1(n_17),
.B2(n_30),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_31),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_1),
.B(n_2),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_31),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_79),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_13),
.C(n_15),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_82),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_47),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_25),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_72),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_83),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_46),
.C(n_45),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_77),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_87),
.B1(n_92),
.B2(n_102),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_58),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_89),
.B(n_99),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_74),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_50),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_93),
.B(n_96),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_37),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_25),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_28),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_17),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_62),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_72),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_51),
.B1(n_36),
.B2(n_35),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_101),
.A2(n_81),
.B1(n_75),
.B2(n_64),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_36),
.B1(n_32),
.B2(n_29),
.Y(n_102)
);

AOI22x1_ASAP7_75t_SL g104 ( 
.A1(n_99),
.A2(n_89),
.B1(n_93),
.B2(n_84),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_104),
.A2(n_114),
.B(n_1),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_115),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_69),
.B1(n_77),
.B2(n_67),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_111),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_62),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_117),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_75),
.B1(n_65),
.B2(n_36),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_95),
.B1(n_94),
.B2(n_101),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_11),
.B(n_14),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_37),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_12),
.B(n_10),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_98),
.B(n_2),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_72),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_65),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_120),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_125),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_126),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_103),
.C(n_94),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_118),
.C(n_115),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_97),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_137),
.Y(n_142)
);

AOI22x1_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_62),
.B1(n_47),
.B2(n_64),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_107),
.B1(n_110),
.B2(n_108),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_106),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_104),
.B1(n_106),
.B2(n_122),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_145),
.Y(n_155)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_149),
.C(n_54),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_105),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_152),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_138),
.B(n_127),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_107),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_54),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_148),
.C(n_149),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_128),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_164),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_132),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_159),
.B(n_146),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_154),
.A2(n_133),
.B1(n_123),
.B2(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_163),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_123),
.B(n_129),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_162),
.A2(n_142),
.B(n_6),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_150),
.A2(n_129),
.B1(n_130),
.B2(n_134),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_3),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_153),
.C(n_151),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_166),
.C(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_147),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_172),
.Y(n_180)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_161),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_152),
.B(n_142),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_176),
.B(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_175),
.B(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_178),
.B(n_179),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_170),
.B(n_162),
.Y(n_181)
);

OAI221xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_168),
.B1(n_170),
.B2(n_167),
.C(n_8),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_5),
.B(n_6),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_168),
.B1(n_173),
.B2(n_174),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_176),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_185),
.Y(n_193)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_187),
.A2(n_7),
.B(n_8),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_189),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_7),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_178),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_186),
.C(n_54),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_195),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_191),
.B(n_9),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_197),
.Y(n_199)
);


endmodule