module fake_netlist_5_1816_n_1712 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1712);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1712;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_53),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_24),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_41),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_46),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_113),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_77),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_43),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_29),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_1),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_5),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_101),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_97),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_75),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

BUFx2_ASAP7_75t_SL g173 ( 
.A(n_151),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_58),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_4),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_7),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_78),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_39),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_132),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_130),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_25),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_34),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_93),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_23),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_76),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_89),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_10),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_119),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_62),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_102),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_103),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_152),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_81),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_146),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_42),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_1),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_117),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_28),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_18),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_41),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_107),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_30),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_42),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_13),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_143),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_96),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_106),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_59),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_84),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_67),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_35),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_60),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_21),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_23),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_128),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_121),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_55),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_144),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_82),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_126),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_50),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_3),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_10),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_74),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_155),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_145),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_50),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_95),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_142),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_3),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_131),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_105),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_122),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_9),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_129),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_49),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_9),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_153),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_17),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_71),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_92),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_98),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_17),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_21),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_45),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_118),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_7),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_120),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_40),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_46),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_13),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_111),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_22),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_14),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_64),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_20),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_88),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_43),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_147),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_44),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_53),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_94),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_66),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_123),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_31),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_134),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_63),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_108),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_38),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_137),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_16),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_61),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_79),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_73),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_133),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_44),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_112),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_39),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_30),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_27),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_2),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_19),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_100),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_36),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_6),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_114),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_140),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_4),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_127),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_139),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_33),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_85),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_47),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_25),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_148),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_57),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_52),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_104),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_27),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_37),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_51),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_15),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_26),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_56),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_72),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_215),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_157),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_193),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_195),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_157),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_196),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_157),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_234),
.B(n_0),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_229),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_191),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_186),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_157),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_157),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_215),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_215),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_198),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_156),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_218),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_199),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_0),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_198),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_203),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_303),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_207),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_219),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_156),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_205),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_234),
.B(n_2),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_176),
.B(n_183),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_L g343 ( 
.A(n_165),
.B(n_5),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_164),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_250),
.B(n_8),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_281),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_281),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_285),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_209),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_210),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_259),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_217),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_194),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_221),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_222),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_237),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_185),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_205),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_201),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_240),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_158),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_202),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_165),
.B(n_8),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_248),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_257),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_264),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_268),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_269),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_204),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_197),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_200),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_206),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_235),
.B(n_11),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_235),
.B(n_11),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_213),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_216),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_180),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_159),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_224),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_223),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_247),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_309),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_309),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_312),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_312),
.Y(n_385)
);

OR2x6_ASAP7_75t_L g386 ( 
.A(n_316),
.B(n_173),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_314),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_159),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_317),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_314),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_320),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_344),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_320),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_319),
.A2(n_339),
.B(n_323),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_344),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_161),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_322),
.B(n_180),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_344),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_374),
.B(n_161),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_321),
.B(n_162),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_344),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_344),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_308),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_308),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_323),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_324),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_322),
.B(n_346),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_324),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_346),
.B(n_220),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_L g415 ( 
.A(n_341),
.B(n_258),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_329),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_347),
.B(n_162),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_343),
.B(n_220),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_332),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_332),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_370),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_333),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_347),
.B(n_169),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_333),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_336),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_359),
.B(n_169),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_336),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_340),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_341),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_340),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_342),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_342),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_343),
.B(n_265),
.Y(n_437)
);

OA21x2_ASAP7_75t_L g438 ( 
.A1(n_359),
.A2(n_239),
.B(n_232),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_362),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_362),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_369),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_369),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_372),
.B(n_170),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_380),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_363),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_337),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_328),
.B(n_170),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_438),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_396),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_420),
.Y(n_453)
);

BUFx6f_ASAP7_75t_SL g454 ( 
.A(n_386),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_396),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_447),
.B(n_164),
.Y(n_456)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_391),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_447),
.B(n_449),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_411),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_420),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_411),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_420),
.Y(n_462)
);

INVx4_ASAP7_75t_SL g463 ( 
.A(n_398),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_391),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_420),
.B(n_310),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_396),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_420),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_425),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_411),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_398),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_418),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_418),
.Y(n_472)
);

INVx8_ASAP7_75t_L g473 ( 
.A(n_386),
.Y(n_473)
);

OAI22xp33_ASAP7_75t_L g474 ( 
.A1(n_450),
.A2(n_348),
.B1(n_163),
.B2(n_182),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_420),
.B(n_311),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_447),
.B(n_172),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_433),
.B(n_371),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_449),
.B(n_437),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_425),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_433),
.B(n_388),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_449),
.B(n_172),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_423),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_450),
.B(n_313),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_399),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_423),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_437),
.B(n_208),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_399),
.Y(n_489)
);

OR2x6_ASAP7_75t_L g490 ( 
.A(n_386),
.B(n_258),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_389),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_398),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_391),
.Y(n_493)
);

OR2x6_ASAP7_75t_L g494 ( 
.A(n_386),
.B(n_265),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_437),
.B(n_327),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_399),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_437),
.B(n_331),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_437),
.B(n_334),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_437),
.B(n_349),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_399),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_400),
.B(n_350),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_382),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_433),
.B(n_400),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_439),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_403),
.B(n_352),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_403),
.B(n_354),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_388),
.B(n_355),
.Y(n_507)
);

BUFx10_ASAP7_75t_L g508 ( 
.A(n_386),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_425),
.B(n_375),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_440),
.B(n_208),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_382),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_386),
.A2(n_364),
.B1(n_356),
.B2(n_360),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_419),
.B(n_366),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_404),
.B(n_367),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_382),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_385),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_389),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_385),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_385),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_448),
.B(n_361),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_387),
.Y(n_521)
);

BUFx4f_ASAP7_75t_L g522 ( 
.A(n_438),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_419),
.B(n_368),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_448),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_427),
.B(n_325),
.Y(n_525)
);

BUFx4f_ASAP7_75t_L g526 ( 
.A(n_438),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_391),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_387),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_386),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_440),
.B(n_270),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_439),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_404),
.B(n_376),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_446),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_446),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_446),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_427),
.B(n_379),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_401),
.B(n_168),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_387),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_383),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_391),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_391),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_415),
.A2(n_365),
.B1(n_378),
.B2(n_353),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_393),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_430),
.B(n_315),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_413),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_L g546 ( 
.A(n_409),
.B(n_186),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_394),
.Y(n_547)
);

AND2x4_ASAP7_75t_SL g548 ( 
.A(n_413),
.B(n_318),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_393),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_394),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_394),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_440),
.B(n_270),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_393),
.Y(n_553)
);

OAI22xp33_ASAP7_75t_L g554 ( 
.A1(n_430),
.A2(n_189),
.B1(n_345),
.B2(n_252),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_395),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_415),
.A2(n_256),
.B1(n_245),
.B2(n_249),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_444),
.B(n_381),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_383),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_402),
.B(n_214),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_444),
.B(n_338),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_384),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_409),
.B(n_186),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_402),
.B(n_274),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_384),
.Y(n_564)
);

BUFx10_ASAP7_75t_L g565 ( 
.A(n_409),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_401),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_390),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_390),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_402),
.B(n_274),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_L g570 ( 
.A(n_409),
.B(n_186),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_441),
.B(n_358),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_402),
.B(n_405),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_395),
.Y(n_573)
);

INVxp67_ASAP7_75t_SL g574 ( 
.A(n_393),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_440),
.B(n_188),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_441),
.B(n_326),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_392),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_392),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_441),
.B(n_351),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_438),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_438),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_438),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_395),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_405),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_441),
.B(n_335),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_393),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_397),
.Y(n_587)
);

INVx8_ASAP7_75t_L g588 ( 
.A(n_440),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_397),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_405),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_410),
.Y(n_591)
);

AND2x6_ASAP7_75t_L g592 ( 
.A(n_406),
.B(n_211),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_406),
.B(n_212),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_440),
.B(n_226),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_412),
.B(n_247),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_459),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_520),
.B(n_158),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_501),
.B(n_397),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_506),
.B(n_440),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_525),
.B(n_536),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_451),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_485),
.B(n_440),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_581),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_482),
.B(n_171),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_581),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_513),
.B(n_443),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_523),
.B(n_443),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_524),
.B(n_160),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_505),
.B(n_503),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_557),
.B(n_171),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_502),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_479),
.B(n_560),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_461),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_469),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_503),
.B(n_443),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_544),
.B(n_174),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_502),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_566),
.B(n_576),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_507),
.B(n_443),
.Y(n_619)
);

AND2x6_ASAP7_75t_SL g620 ( 
.A(n_509),
.B(n_253),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_471),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_532),
.B(n_514),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_545),
.B(n_174),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_480),
.B(n_443),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_458),
.B(n_443),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_579),
.B(n_177),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_458),
.B(n_443),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_585),
.A2(n_192),
.B1(n_190),
.B2(n_187),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_453),
.B(n_406),
.Y(n_629)
);

INVxp67_ASAP7_75t_SL g630 ( 
.A(n_470),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_511),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_SL g632 ( 
.A(n_468),
.B(n_246),
.C(n_238),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_481),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_472),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_548),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_484),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_460),
.B(n_409),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_554),
.B(n_177),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_571),
.B(n_595),
.Y(n_639)
);

NOR3xp33_ASAP7_75t_L g640 ( 
.A(n_517),
.B(n_241),
.C(n_236),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_511),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_491),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_460),
.B(n_409),
.Y(n_643)
);

OAI221xp5_ASAP7_75t_L g644 ( 
.A1(n_556),
.A2(n_284),
.B1(n_260),
.B2(n_255),
.C(n_282),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_462),
.B(n_409),
.Y(n_645)
);

O2A1O1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_580),
.A2(n_445),
.B(n_442),
.C(n_271),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_515),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_462),
.B(n_409),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_465),
.B(n_179),
.Y(n_649)
);

BUFx12f_ASAP7_75t_SL g650 ( 
.A(n_494),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_522),
.B(n_186),
.Y(n_651)
);

A2O1A1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_522),
.A2(n_231),
.B(n_227),
.C(n_230),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_467),
.B(n_408),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_477),
.B(n_179),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_582),
.A2(n_287),
.B1(n_290),
.B2(n_299),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_495),
.B(n_181),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_497),
.B(n_181),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_487),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_522),
.B(n_186),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_498),
.B(n_184),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_481),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_548),
.B(n_412),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_542),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_504),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_537),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_467),
.B(n_408),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_526),
.B(n_186),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_533),
.B(n_408),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_470),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_515),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_537),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_534),
.B(n_442),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_531),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_535),
.B(n_442),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_470),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_539),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_537),
.B(n_412),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_558),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_516),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_499),
.B(n_184),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_561),
.B(n_442),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_470),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_474),
.B(n_187),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_564),
.B(n_567),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_568),
.B(n_445),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_456),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_577),
.B(n_190),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_526),
.B(n_186),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_578),
.Y(n_689)
);

INVx5_ASAP7_75t_L g690 ( 
.A(n_588),
.Y(n_690)
);

AOI221xp5_ASAP7_75t_L g691 ( 
.A1(n_512),
.A2(n_286),
.B1(n_283),
.B2(n_293),
.C(n_225),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_508),
.B(n_529),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_516),
.Y(n_693)
);

NAND2x1p5_ASAP7_75t_L g694 ( 
.A(n_526),
.B(n_243),
.Y(n_694)
);

BUFx8_ASAP7_75t_L g695 ( 
.A(n_454),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_518),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_518),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_508),
.B(n_192),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_519),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_454),
.A2(n_228),
.B1(n_272),
.B2(n_275),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_456),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_559),
.B(n_490),
.Y(n_702)
);

AO22x2_ASAP7_75t_L g703 ( 
.A1(n_587),
.A2(n_306),
.B1(n_254),
.B2(n_261),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_587),
.A2(n_267),
.B1(n_266),
.B2(n_307),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_519),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_508),
.B(n_272),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_475),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_529),
.B(n_475),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_529),
.B(n_266),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_475),
.B(n_275),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_589),
.A2(n_266),
.B1(n_291),
.B2(n_244),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_490),
.B(n_279),
.Y(n_712)
);

O2A1O1Ixp5_ASAP7_75t_L g713 ( 
.A1(n_488),
.A2(n_478),
.B(n_483),
.C(n_510),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_L g714 ( 
.A(n_473),
.B(n_266),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_490),
.B(n_414),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_583),
.B(n_445),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_492),
.B(n_445),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_521),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_521),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_584),
.B(n_407),
.Y(n_720)
);

INVx8_ASAP7_75t_L g721 ( 
.A(n_473),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_475),
.B(n_279),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_528),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_490),
.B(n_414),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_589),
.A2(n_266),
.B1(n_276),
.B2(n_298),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_590),
.B(n_494),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_473),
.B(n_292),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_494),
.Y(n_728)
);

CKINVDCx16_ASAP7_75t_R g729 ( 
.A(n_454),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_478),
.B(n_414),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_574),
.B(n_407),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_528),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_488),
.B(n_407),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_538),
.Y(n_734)
);

BUFx4_ASAP7_75t_L g735 ( 
.A(n_593),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_483),
.Y(n_736)
);

BUFx5_ASAP7_75t_L g737 ( 
.A(n_565),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_541),
.B(n_407),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_494),
.B(n_160),
.Y(n_739)
);

NOR2xp67_ASAP7_75t_SL g740 ( 
.A(n_493),
.B(n_393),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_563),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_569),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_541),
.B(n_417),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_538),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_541),
.B(n_417),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_473),
.A2(n_266),
.B1(n_277),
.B2(n_289),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_575),
.A2(n_594),
.B1(n_592),
.B2(n_572),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_547),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_594),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_549),
.B(n_417),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_547),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_549),
.B(n_417),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_550),
.B(n_266),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_549),
.B(n_417),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_586),
.B(n_417),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_550),
.B(n_292),
.Y(n_756)
);

INVx8_ASAP7_75t_L g757 ( 
.A(n_592),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_551),
.B(n_266),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_551),
.B(n_294),
.Y(n_759)
);

AO22x1_ASAP7_75t_L g760 ( 
.A1(n_592),
.A2(n_166),
.B1(n_167),
.B2(n_175),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_555),
.B(n_393),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_598),
.A2(n_466),
.B(n_452),
.Y(n_762)
);

OAI321xp33_ASAP7_75t_L g763 ( 
.A1(n_616),
.A2(n_530),
.A3(n_510),
.B1(n_552),
.B2(n_416),
.C(n_426),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_642),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_611),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_690),
.A2(n_588),
.B(n_540),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_622),
.B(n_639),
.Y(n_767)
);

NOR2x1_ASAP7_75t_L g768 ( 
.A(n_612),
.B(n_555),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_622),
.B(n_573),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_690),
.A2(n_607),
.B(n_606),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_600),
.B(n_463),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_690),
.A2(n_588),
.B(n_553),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_609),
.B(n_573),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_611),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_704),
.A2(n_530),
.B1(n_552),
.B2(n_586),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_610),
.B(n_586),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_616),
.A2(n_546),
.B(n_562),
.C(n_570),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_690),
.A2(n_588),
.B(n_476),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_610),
.B(n_452),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_599),
.A2(n_476),
.B(n_464),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_602),
.A2(n_476),
.B(n_464),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_704),
.A2(n_294),
.B1(n_297),
.B2(n_527),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_605),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_605),
.B(n_463),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_605),
.B(n_463),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_619),
.A2(n_464),
.B(n_540),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_662),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_633),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_721),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_596),
.A2(n_546),
.B(n_570),
.C(n_562),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_626),
.B(n_455),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_661),
.Y(n_792)
);

AO21x1_ASAP7_75t_L g793 ( 
.A1(n_626),
.A2(n_540),
.B(n_553),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_741),
.B(n_455),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_618),
.B(n_543),
.Y(n_795)
);

NOR3xp33_ASAP7_75t_L g796 ( 
.A(n_632),
.B(n_297),
.C(n_262),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_677),
.B(n_466),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_617),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_702),
.A2(n_592),
.B1(n_543),
.B2(n_553),
.Y(n_799)
);

O2A1O1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_613),
.A2(n_614),
.B(n_659),
.C(n_651),
.Y(n_800)
);

AND2x2_ASAP7_75t_SL g801 ( 
.A(n_714),
.B(n_543),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_637),
.A2(n_493),
.B(n_527),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_691),
.B(n_251),
.C(n_263),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_643),
.A2(n_648),
.B(n_645),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_623),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_624),
.A2(n_527),
.B(n_457),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_702),
.A2(n_654),
.B1(n_660),
.B2(n_657),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_635),
.Y(n_808)
);

A2O1A1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_604),
.A2(n_657),
.B(n_660),
.C(n_736),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_665),
.B(n_233),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_651),
.A2(n_489),
.B(n_486),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_731),
.A2(n_457),
.B(n_393),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_659),
.A2(n_489),
.B(n_486),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_604),
.A2(n_496),
.B(n_500),
.C(n_591),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_630),
.A2(n_457),
.B(n_500),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_667),
.A2(n_591),
.B(n_496),
.C(n_428),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_671),
.B(n_416),
.Y(n_817)
);

INVxp67_ASAP7_75t_L g818 ( 
.A(n_623),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_675),
.A2(n_457),
.B(n_565),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_655),
.A2(n_592),
.B1(n_305),
.B2(n_301),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_667),
.A2(n_426),
.B(n_428),
.C(n_434),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_688),
.A2(n_426),
.B(n_428),
.C(n_434),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_737),
.B(n_233),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_726),
.A2(n_592),
.B1(n_431),
.B2(n_434),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_715),
.B(n_431),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_695),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_724),
.B(n_621),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_686),
.A2(n_431),
.B(n_432),
.C(n_435),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_688),
.A2(n_435),
.B(n_432),
.C(n_410),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_597),
.B(n_166),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_663),
.B(n_167),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_629),
.A2(n_457),
.B(n_565),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_713),
.A2(n_410),
.B(n_435),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_717),
.A2(n_424),
.B(n_435),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_701),
.A2(n_410),
.B(n_432),
.C(n_429),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_653),
.A2(n_432),
.B(n_429),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_601),
.B(n_421),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_726),
.A2(n_421),
.B(n_429),
.C(n_424),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_601),
.B(n_421),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_638),
.B(n_175),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_737),
.B(n_233),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_R g842 ( 
.A(n_650),
.B(n_178),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_669),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_603),
.B(n_421),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_666),
.A2(n_429),
.B(n_424),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_631),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_615),
.A2(n_627),
.B(n_625),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_608),
.B(n_286),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_603),
.B(n_436),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_742),
.A2(n_436),
.B(n_422),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_728),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_683),
.B(n_178),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_694),
.A2(n_225),
.B(n_273),
.Y(n_853)
);

BUFx8_ASAP7_75t_L g854 ( 
.A(n_739),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_631),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_641),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_707),
.A2(n_436),
.B(n_422),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_737),
.B(n_242),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_641),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_628),
.B(n_305),
.Y(n_860)
);

NOR2xp67_ASAP7_75t_L g861 ( 
.A(n_700),
.B(n_634),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_707),
.A2(n_436),
.B(n_422),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_709),
.A2(n_242),
.B(n_288),
.C(n_278),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_636),
.B(n_658),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_712),
.B(n_664),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_721),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_673),
.B(n_676),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_709),
.A2(n_436),
.B(n_422),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_712),
.B(n_283),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_733),
.A2(n_436),
.B(n_422),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_669),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_649),
.B(n_301),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_761),
.A2(n_436),
.B(n_422),
.Y(n_873)
);

NOR2x1_ASAP7_75t_R g874 ( 
.A(n_698),
.B(n_273),
.Y(n_874)
);

AOI33xp33_ASAP7_75t_L g875 ( 
.A1(n_655),
.A2(n_278),
.A3(n_280),
.B1(n_293),
.B2(n_295),
.B3(n_242),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_669),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_678),
.B(n_295),
.Y(n_877)
);

INVxp67_ASAP7_75t_SL g878 ( 
.A(n_669),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_694),
.A2(n_280),
.B(n_288),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_721),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_757),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_708),
.A2(n_436),
.B(n_422),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_757),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_737),
.B(n_684),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_708),
.A2(n_422),
.B(n_417),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_695),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_743),
.A2(n_417),
.B(n_115),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_SL g888 ( 
.A1(n_652),
.A2(n_288),
.B(n_14),
.C(n_15),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_687),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_745),
.A2(n_154),
.B(n_150),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_750),
.A2(n_149),
.B(n_136),
.Y(n_891)
);

AND2x2_ASAP7_75t_SL g892 ( 
.A(n_746),
.B(n_135),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_647),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_757),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_689),
.B(n_12),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_737),
.B(n_125),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_647),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_687),
.A2(n_12),
.B(n_16),
.C(n_18),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_752),
.A2(n_124),
.B(n_116),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_749),
.A2(n_110),
.B1(n_90),
.B2(n_87),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_682),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_682),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_670),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_730),
.B(n_19),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_646),
.A2(n_20),
.B(n_22),
.C(n_24),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_656),
.B(n_26),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_723),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_747),
.A2(n_86),
.B(n_83),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_711),
.A2(n_80),
.B1(n_70),
.B2(n_69),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_680),
.B(n_28),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_670),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_756),
.A2(n_65),
.B1(n_31),
.B2(n_32),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_754),
.A2(n_29),
.B(n_32),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_755),
.A2(n_33),
.B(n_35),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_738),
.A2(n_36),
.B(n_37),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_679),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_SL g917 ( 
.A(n_729),
.B(n_38),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_679),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_737),
.A2(n_40),
.B(n_45),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_756),
.B(n_47),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_640),
.B(n_706),
.Y(n_921)
);

NOR2x1_ASAP7_75t_L g922 ( 
.A(n_692),
.B(n_727),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_759),
.B(n_48),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_760),
.B(n_54),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_681),
.A2(n_48),
.B(n_49),
.Y(n_925)
);

AOI21x1_ASAP7_75t_L g926 ( 
.A1(n_761),
.A2(n_51),
.B(n_52),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_735),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_693),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_SL g929 ( 
.A1(n_753),
.A2(n_54),
.B(n_758),
.C(n_710),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_723),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_693),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_753),
.A2(n_758),
.B(n_644),
.C(n_716),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_697),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_697),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_759),
.B(n_685),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_719),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_672),
.A2(n_674),
.B(n_720),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_668),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_719),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_732),
.B(n_751),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_696),
.A2(n_748),
.B(n_699),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_732),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_767),
.B(n_734),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_866),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_805),
.B(n_620),
.Y(n_945)
);

BUFx4f_ASAP7_75t_L g946 ( 
.A(n_866),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_936),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_770),
.A2(n_722),
.B(n_746),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_889),
.B(n_751),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_783),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_892),
.A2(n_725),
.B1(n_711),
.B2(n_703),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_764),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_SL g953 ( 
.A1(n_809),
.A2(n_705),
.B(n_718),
.C(n_744),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_SL g954 ( 
.A1(n_892),
.A2(n_703),
.B1(n_734),
.B2(n_725),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_827),
.B(n_703),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_884),
.A2(n_740),
.B(n_769),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_873),
.A2(n_804),
.B(n_786),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_SL g958 ( 
.A1(n_923),
.A2(n_935),
.B(n_818),
.C(n_805),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_788),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_935),
.B(n_807),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_923),
.A2(n_818),
.B1(n_920),
.B2(n_908),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_831),
.B(n_787),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_938),
.B(n_865),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_869),
.A2(n_827),
.B1(n_921),
.B2(n_861),
.Y(n_964)
);

NOR3xp33_ASAP7_75t_L g965 ( 
.A(n_831),
.B(n_860),
.C(n_840),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_787),
.B(n_840),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_825),
.B(n_864),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_825),
.B(n_867),
.Y(n_968)
);

AO21x1_ASAP7_75t_L g969 ( 
.A1(n_800),
.A2(n_919),
.B(n_879),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_801),
.A2(n_773),
.B(n_772),
.Y(n_970)
);

AO32x1_ASAP7_75t_L g971 ( 
.A1(n_775),
.A2(n_909),
.A3(n_900),
.B1(n_924),
.B2(n_782),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_866),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_801),
.A2(n_778),
.B(n_766),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_852),
.A2(n_910),
.B(n_906),
.C(n_800),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_866),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_852),
.A2(n_898),
.B(n_803),
.C(n_853),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_872),
.B(n_792),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_847),
.A2(n_777),
.B(n_937),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_783),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_811),
.A2(n_813),
.B(n_833),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_904),
.A2(n_820),
.B1(n_912),
.B2(n_779),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_794),
.B(n_817),
.Y(n_982)
);

BUFx4f_ASAP7_75t_L g983 ( 
.A(n_880),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_780),
.A2(n_781),
.B(n_776),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_820),
.A2(n_895),
.B1(n_791),
.B2(n_878),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_855),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_817),
.B(n_795),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_856),
.Y(n_988)
);

AND2x6_ASAP7_75t_L g989 ( 
.A(n_880),
.B(n_881),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_939),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_797),
.A2(n_802),
.B(n_790),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_880),
.Y(n_992)
);

OR2x6_ASAP7_75t_L g993 ( 
.A(n_927),
.B(n_880),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_851),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_790),
.A2(n_849),
.B(n_878),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_854),
.Y(n_996)
);

BUFx12f_ASAP7_75t_L g997 ( 
.A(n_854),
.Y(n_997)
);

NOR2xp67_ASAP7_75t_SL g998 ( 
.A(n_789),
.B(n_881),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_808),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_837),
.A2(n_839),
.B(n_844),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_922),
.B(n_796),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_789),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_762),
.A2(n_806),
.B(n_819),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_939),
.B(n_859),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_893),
.B(n_897),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_830),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_877),
.B(n_875),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_SL g1008 ( 
.A1(n_917),
.A2(n_848),
.B1(n_925),
.B2(n_913),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_832),
.A2(n_940),
.B(n_896),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_768),
.B(n_911),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_SL g1011 ( 
.A1(n_771),
.A2(n_928),
.B(n_931),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_765),
.B(n_774),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_842),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_881),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_824),
.A2(n_803),
.B1(n_934),
.B2(n_933),
.Y(n_1015)
);

NOR3xp33_ASAP7_75t_L g1016 ( 
.A(n_874),
.B(n_810),
.C(n_796),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_798),
.B(n_942),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_SL g1018 ( 
.A1(n_863),
.A2(n_763),
.B(n_932),
.C(n_843),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_863),
.B(n_930),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_823),
.A2(n_841),
.B(n_858),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_932),
.A2(n_784),
.B(n_785),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_905),
.A2(n_888),
.B(n_929),
.C(n_838),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_907),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_812),
.A2(n_799),
.B(n_815),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_902),
.A2(n_941),
.B(n_814),
.Y(n_1025)
);

BUFx12f_ASAP7_75t_L g1026 ( 
.A(n_826),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_846),
.A2(n_918),
.B1(n_916),
.B2(n_903),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_901),
.B(n_886),
.Y(n_1028)
);

NAND2xp33_ASAP7_75t_SL g1029 ( 
.A(n_881),
.B(n_894),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_907),
.B(n_930),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_930),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_907),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_816),
.A2(n_821),
.B(n_822),
.C(n_905),
.Y(n_1033)
);

CKINVDCx8_ASAP7_75t_R g1034 ( 
.A(n_883),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_901),
.A2(n_857),
.B(n_862),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_843),
.B(n_876),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_883),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_828),
.A2(n_835),
.B(n_915),
.C(n_914),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_871),
.A2(n_876),
.B(n_850),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_871),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_883),
.B(n_894),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_SL g1042 ( 
.A(n_890),
.B(n_899),
.C(n_891),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_834),
.A2(n_885),
.B(n_882),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_822),
.B(n_836),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_926),
.B(n_894),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_883),
.A2(n_894),
.B1(n_845),
.B2(n_829),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_870),
.A2(n_868),
.B(n_829),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_793),
.B(n_887),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_770),
.A2(n_690),
.B(n_460),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_SL g1050 ( 
.A1(n_831),
.A2(n_633),
.B1(n_481),
.B2(n_661),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_939),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_770),
.A2(n_690),
.B(n_460),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_809),
.A2(n_600),
.B(n_616),
.C(n_610),
.Y(n_1053)
);

AO32x1_ASAP7_75t_L g1054 ( 
.A1(n_775),
.A2(n_587),
.A3(n_589),
.B1(n_909),
.B2(n_900),
.Y(n_1054)
);

AND2x4_ASAP7_75t_SL g1055 ( 
.A(n_866),
.B(n_880),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_767),
.B(n_622),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_764),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_831),
.B(n_639),
.Y(n_1058)
);

AO21x1_ASAP7_75t_L g1059 ( 
.A1(n_923),
.A2(n_807),
.B(n_908),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_788),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_809),
.A2(n_600),
.B(n_616),
.C(n_610),
.Y(n_1061)
);

OR2x6_ASAP7_75t_SL g1062 ( 
.A(n_920),
.B(n_661),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_787),
.Y(n_1063)
);

OAI21xp33_ASAP7_75t_SL g1064 ( 
.A1(n_892),
.A2(n_704),
.B(n_807),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_807),
.A2(n_600),
.B1(n_622),
.B2(n_616),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_939),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_767),
.B(n_889),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_936),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_805),
.B(n_600),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_770),
.A2(n_690),
.B(n_460),
.Y(n_1070)
);

AND2x2_ASAP7_75t_SL g1071 ( 
.A(n_892),
.B(n_704),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_807),
.A2(n_600),
.B1(n_622),
.B2(n_616),
.Y(n_1072)
);

OR2x4_ASAP7_75t_L g1073 ( 
.A(n_831),
.B(n_632),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_767),
.B(n_622),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_L g1075 ( 
.A(n_807),
.B(n_610),
.C(n_616),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_770),
.A2(n_690),
.B(n_460),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_767),
.B(n_889),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_764),
.Y(n_1078)
);

O2A1O1Ixp5_ASAP7_75t_L g1079 ( 
.A1(n_793),
.A2(n_600),
.B(n_809),
.C(n_923),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_SL g1080 ( 
.A(n_892),
.B(n_923),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_767),
.B(n_622),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_787),
.Y(n_1082)
);

OAI21xp33_ASAP7_75t_SL g1083 ( 
.A1(n_892),
.A2(n_704),
.B(n_807),
.Y(n_1083)
);

OAI21xp33_ASAP7_75t_L g1084 ( 
.A1(n_869),
.A2(n_616),
.B(n_610),
.Y(n_1084)
);

INVx4_ASAP7_75t_L g1085 ( 
.A(n_866),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1058),
.B(n_962),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_965),
.B(n_966),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_947),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_978),
.A2(n_984),
.B(n_970),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1071),
.A2(n_1072),
.B1(n_1065),
.B2(n_1075),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_957),
.A2(n_1035),
.B(n_973),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_952),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_1028),
.B(n_993),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_1057),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_1084),
.B(n_1056),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1043),
.A2(n_1025),
.B(n_1003),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_1047),
.A2(n_991),
.B(n_1039),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_1074),
.B(n_1081),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_960),
.B(n_1069),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_977),
.B(n_963),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1067),
.B(n_1077),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_978),
.A2(n_1009),
.B(n_1076),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1064),
.A2(n_1083),
.B(n_1075),
.C(n_1053),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1049),
.A2(n_1052),
.B(n_1070),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1024),
.A2(n_1048),
.B(n_948),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1020),
.A2(n_1061),
.B(n_956),
.Y(n_1106)
);

AOI221xp5_ASAP7_75t_L g1107 ( 
.A1(n_976),
.A2(n_961),
.B1(n_974),
.B2(n_981),
.C(n_1080),
.Y(n_1107)
);

AO31x2_ASAP7_75t_L g1108 ( 
.A1(n_1059),
.A2(n_969),
.A3(n_961),
.B(n_1033),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_951),
.A2(n_981),
.A3(n_995),
.B(n_985),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1044),
.A2(n_1000),
.B(n_1042),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1068),
.Y(n_1111)
);

CKINVDCx8_ASAP7_75t_R g1112 ( 
.A(n_996),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_967),
.B(n_968),
.Y(n_1113)
);

NAND3x1_ASAP7_75t_L g1114 ( 
.A(n_1016),
.B(n_945),
.C(n_964),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_987),
.A2(n_1080),
.B(n_953),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_SL g1116 ( 
.A1(n_951),
.A2(n_958),
.B(n_1018),
.C(n_1001),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_982),
.B(n_943),
.Y(n_1117)
);

NAND2x1_ASAP7_75t_L g1118 ( 
.A(n_989),
.B(n_998),
.Y(n_1118)
);

CKINVDCx11_ASAP7_75t_R g1119 ( 
.A(n_997),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1046),
.A2(n_980),
.B(n_1021),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1006),
.B(n_1007),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1046),
.A2(n_971),
.B(n_1054),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1063),
.B(n_1082),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_985),
.B(n_1008),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1008),
.B(n_949),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_1079),
.A2(n_1022),
.B(n_1019),
.C(n_1038),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_986),
.Y(n_1127)
);

AND3x4_ASAP7_75t_L g1128 ( 
.A(n_959),
.B(n_1060),
.C(n_1050),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1015),
.A2(n_954),
.B(n_1011),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1015),
.A2(n_971),
.A3(n_1054),
.B(n_1010),
.Y(n_1130)
);

NOR2x1_ASAP7_75t_R g1131 ( 
.A(n_1026),
.B(n_1085),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1057),
.B(n_988),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_994),
.A2(n_1078),
.B(n_1013),
.C(n_955),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1005),
.B(n_955),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_971),
.A2(n_1054),
.B(n_1029),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_999),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1005),
.A2(n_1045),
.B(n_1030),
.C(n_1004),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_990),
.A2(n_1051),
.B1(n_1066),
.B2(n_1040),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1004),
.A2(n_1012),
.B(n_1041),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_993),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_946),
.A2(n_983),
.B(n_1036),
.Y(n_1141)
);

BUFx12f_ASAP7_75t_L g1142 ( 
.A(n_993),
.Y(n_1142)
);

AOI221xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1027),
.A2(n_1031),
.B1(n_944),
.B2(n_972),
.C(n_975),
.Y(n_1143)
);

CKINVDCx8_ASAP7_75t_R g1144 ( 
.A(n_944),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_SL g1145 ( 
.A1(n_1023),
.A2(n_1032),
.B(n_950),
.C(n_979),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1073),
.A2(n_979),
.B(n_950),
.C(n_1062),
.Y(n_1146)
);

NOR2xp67_ASAP7_75t_L g1147 ( 
.A(n_1085),
.B(n_1002),
.Y(n_1147)
);

AO31x2_ASAP7_75t_L g1148 ( 
.A1(n_1073),
.A2(n_989),
.A3(n_1034),
.B(n_946),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_983),
.B(n_1002),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_944),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_972),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1055),
.A2(n_1002),
.B(n_1014),
.C(n_1037),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_989),
.A2(n_1014),
.A3(n_1037),
.B(n_992),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_972),
.B(n_975),
.Y(n_1154)
);

BUFx8_ASAP7_75t_SL g1155 ( 
.A(n_975),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1037),
.A2(n_992),
.B(n_989),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_992),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_978),
.A2(n_690),
.B(n_770),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1075),
.A2(n_1084),
.B(n_1061),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1075),
.A2(n_1083),
.B(n_1064),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1071),
.A2(n_1072),
.B1(n_1065),
.B2(n_1075),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1028),
.B(n_827),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_978),
.A2(n_690),
.B(n_770),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_947),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1084),
.B(n_600),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1056),
.B(n_1074),
.Y(n_1166)
);

CKINVDCx11_ASAP7_75t_R g1167 ( 
.A(n_997),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_1059),
.A2(n_969),
.A3(n_793),
.B(n_1048),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1028),
.B(n_827),
.Y(n_1169)
);

NAND3x1_ASAP7_75t_L g1170 ( 
.A(n_965),
.B(n_803),
.C(n_860),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_947),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1056),
.B(n_1074),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_SL g1173 ( 
.A(n_997),
.B(n_1034),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_965),
.B(n_1084),
.C(n_600),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_965),
.A2(n_600),
.B(n_1084),
.C(n_974),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_978),
.A2(n_690),
.B(n_770),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1056),
.B(n_1074),
.Y(n_1177)
);

AO22x2_ASAP7_75t_L g1178 ( 
.A1(n_961),
.A2(n_965),
.B1(n_1075),
.B2(n_951),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1056),
.B(n_1074),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1075),
.A2(n_1083),
.B(n_1064),
.Y(n_1180)
);

OA21x2_ASAP7_75t_L g1181 ( 
.A1(n_978),
.A2(n_1048),
.B(n_980),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_978),
.A2(n_690),
.B(n_770),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1017),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_965),
.A2(n_600),
.B(n_1084),
.C(n_974),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_978),
.A2(n_690),
.B(n_770),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1059),
.A2(n_969),
.A3(n_793),
.B(n_1048),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1056),
.B(n_1074),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1075),
.A2(n_1084),
.B(n_1061),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1028),
.B(n_827),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_978),
.A2(n_690),
.B(n_770),
.Y(n_1190)
);

BUFx10_ASAP7_75t_L g1191 ( 
.A(n_945),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_944),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_978),
.A2(n_690),
.B(n_770),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1058),
.B(n_962),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1059),
.A2(n_969),
.A3(n_793),
.B(n_1048),
.Y(n_1195)
);

CKINVDCx16_ASAP7_75t_R g1196 ( 
.A(n_1050),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1084),
.A2(n_1083),
.B(n_1064),
.C(n_1075),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_1059),
.A2(n_969),
.A3(n_793),
.B(n_1048),
.Y(n_1198)
);

AOI211x1_ASAP7_75t_L g1199 ( 
.A1(n_1075),
.A2(n_1059),
.B(n_1084),
.C(n_960),
.Y(n_1199)
);

NOR2xp67_ASAP7_75t_SL g1200 ( 
.A(n_997),
.B(n_1034),
.Y(n_1200)
);

OA21x2_ASAP7_75t_L g1201 ( 
.A1(n_978),
.A2(n_1048),
.B(n_980),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1071),
.A2(n_1072),
.B1(n_1065),
.B2(n_1075),
.Y(n_1202)
);

CKINVDCx11_ASAP7_75t_R g1203 ( 
.A(n_997),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_957),
.A2(n_1035),
.B(n_973),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1017),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_978),
.A2(n_690),
.B(n_770),
.Y(n_1206)
);

OA21x2_ASAP7_75t_L g1207 ( 
.A1(n_978),
.A2(n_1048),
.B(n_980),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_947),
.Y(n_1208)
);

AO22x1_ASAP7_75t_L g1209 ( 
.A1(n_965),
.A2(n_831),
.B1(n_616),
.B2(n_610),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1028),
.B(n_827),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1080),
.A2(n_965),
.B1(n_1071),
.B2(n_1084),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_978),
.A2(n_690),
.B(n_770),
.Y(n_1212)
);

O2A1O1Ixp5_ASAP7_75t_SL g1213 ( 
.A1(n_961),
.A2(n_600),
.B(n_1001),
.C(n_879),
.Y(n_1213)
);

AO32x2_ASAP7_75t_L g1214 ( 
.A1(n_961),
.A2(n_981),
.A3(n_985),
.B1(n_951),
.B2(n_1015),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1056),
.B(n_1074),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_957),
.A2(n_1035),
.B(n_973),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_957),
.A2(n_1035),
.B(n_973),
.Y(n_1217)
);

NOR4xp25_ASAP7_75t_L g1218 ( 
.A(n_1084),
.B(n_1075),
.C(n_976),
.D(n_974),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1028),
.B(n_827),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_957),
.A2(n_1035),
.B(n_973),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_957),
.A2(n_1035),
.B(n_973),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_957),
.A2(n_1035),
.B(n_973),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1034),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_978),
.A2(n_690),
.B(n_770),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1058),
.B(n_962),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_978),
.A2(n_690),
.B(n_770),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1056),
.B(n_1074),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_957),
.A2(n_1035),
.B(n_973),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_978),
.A2(n_690),
.B(n_770),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1127),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1088),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1170),
.A2(n_1100),
.B1(n_1099),
.B2(n_1211),
.Y(n_1232)
);

BUFx10_ASAP7_75t_L g1233 ( 
.A(n_1162),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_SL g1234 ( 
.A1(n_1090),
.A2(n_1202),
.B1(n_1161),
.B2(n_1087),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1166),
.B(n_1172),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1211),
.A2(n_1098),
.B1(n_1227),
.B2(n_1177),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1155),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1179),
.A2(n_1215),
.B1(n_1187),
.B2(n_1095),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1209),
.A2(n_1114),
.B1(n_1174),
.B2(n_1165),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1107),
.A2(n_1178),
.B1(n_1159),
.B2(n_1188),
.Y(n_1240)
);

BUFx8_ASAP7_75t_SL g1241 ( 
.A(n_1092),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1178),
.A2(n_1160),
.B1(n_1180),
.B2(n_1124),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1164),
.Y(n_1243)
);

BUFx12f_ASAP7_75t_L g1244 ( 
.A(n_1119),
.Y(n_1244)
);

INVx6_ASAP7_75t_L g1245 ( 
.A(n_1142),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1160),
.A2(n_1180),
.B1(n_1129),
.B2(n_1225),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1113),
.B(n_1086),
.Y(n_1247)
);

NAND2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1118),
.B(n_1173),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1109),
.Y(n_1249)
);

BUFx2_ASAP7_75t_SL g1250 ( 
.A(n_1144),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1126),
.A2(n_1094),
.B1(n_1134),
.B2(n_1101),
.Y(n_1251)
);

CKINVDCx9p33_ASAP7_75t_R g1252 ( 
.A(n_1140),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1171),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1150),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1196),
.A2(n_1132),
.B1(n_1121),
.B2(n_1117),
.Y(n_1255)
);

BUFx12f_ASAP7_75t_L g1256 ( 
.A(n_1167),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1094),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1183),
.B(n_1205),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1109),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1199),
.A2(n_1197),
.B1(n_1125),
.B2(n_1103),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1111),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1203),
.Y(n_1262)
);

CKINVDCx11_ASAP7_75t_R g1263 ( 
.A(n_1112),
.Y(n_1263)
);

INVx3_ASAP7_75t_SL g1264 ( 
.A(n_1223),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1191),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1115),
.A2(n_1208),
.B1(n_1191),
.B2(n_1123),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1218),
.A2(n_1223),
.B1(n_1214),
.B2(n_1122),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1199),
.A2(n_1175),
.B1(n_1184),
.B2(n_1138),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1192),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1093),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1139),
.Y(n_1271)
);

BUFx2_ASAP7_75t_SL g1272 ( 
.A(n_1147),
.Y(n_1272)
);

OAI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1218),
.A2(n_1136),
.B1(n_1135),
.B2(n_1141),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1153),
.Y(n_1274)
);

CKINVDCx14_ASAP7_75t_R g1275 ( 
.A(n_1162),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1157),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1106),
.A2(n_1128),
.B1(n_1105),
.B2(n_1093),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1145),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1192),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1154),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1181),
.A2(n_1201),
.B1(n_1207),
.B2(n_1110),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1192),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_1149),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1133),
.A2(n_1137),
.B1(n_1169),
.B2(n_1189),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_SL g1285 ( 
.A1(n_1146),
.A2(n_1219),
.B(n_1210),
.Y(n_1285)
);

INVx4_ASAP7_75t_L g1286 ( 
.A(n_1131),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1152),
.A2(n_1147),
.B1(n_1151),
.B2(n_1229),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1181),
.A2(n_1207),
.B1(n_1201),
.B2(n_1089),
.Y(n_1288)
);

BUFx12f_ASAP7_75t_L g1289 ( 
.A(n_1131),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1148),
.B(n_1200),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1156),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1148),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1214),
.A2(n_1102),
.B1(n_1120),
.B2(n_1116),
.Y(n_1293)
);

BUFx12f_ASAP7_75t_L g1294 ( 
.A(n_1213),
.Y(n_1294)
);

INVx6_ASAP7_75t_L g1295 ( 
.A(n_1143),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1158),
.A2(n_1190),
.B1(n_1212),
.B2(n_1206),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1163),
.A2(n_1176),
.B1(n_1224),
.B2(n_1193),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_1143),
.Y(n_1298)
);

CKINVDCx11_ASAP7_75t_R g1299 ( 
.A(n_1108),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1108),
.B(n_1214),
.Y(n_1300)
);

CKINVDCx6p67_ASAP7_75t_R g1301 ( 
.A(n_1168),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1182),
.A2(n_1226),
.B1(n_1185),
.B2(n_1109),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1168),
.B(n_1198),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1168),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1104),
.A2(n_1198),
.B1(n_1186),
.B2(n_1195),
.Y(n_1305)
);

CKINVDCx6p67_ASAP7_75t_R g1306 ( 
.A(n_1186),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1096),
.A2(n_1097),
.B1(n_1130),
.B2(n_1198),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1091),
.A2(n_1217),
.B1(n_1222),
.B2(n_1204),
.Y(n_1308)
);

BUFx2_ASAP7_75t_SL g1309 ( 
.A(n_1195),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1130),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1216),
.A2(n_1220),
.B1(n_1221),
.B2(n_1228),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1127),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1090),
.A2(n_965),
.B1(n_1084),
.B2(n_1075),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1119),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1090),
.A2(n_965),
.B1(n_1084),
.B2(n_1075),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1150),
.Y(n_1316)
);

CKINVDCx11_ASAP7_75t_R g1317 ( 
.A(n_1119),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1090),
.A2(n_965),
.B1(n_1084),
.B2(n_1075),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1094),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1086),
.B(n_1194),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_SL g1321 ( 
.A(n_1162),
.Y(n_1321)
);

CKINVDCx11_ASAP7_75t_R g1322 ( 
.A(n_1119),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1092),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1211),
.A2(n_1080),
.B1(n_1072),
.B2(n_1065),
.Y(n_1324)
);

INVx6_ASAP7_75t_L g1325 ( 
.A(n_1142),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1150),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1092),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1092),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1090),
.A2(n_965),
.B1(n_1084),
.B2(n_1075),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1094),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1119),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1094),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1170),
.A2(n_1071),
.B1(n_1072),
.B2(n_1065),
.Y(n_1333)
);

INVx6_ASAP7_75t_L g1334 ( 
.A(n_1142),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1170),
.A2(n_1071),
.B1(n_1072),
.B2(n_1065),
.Y(n_1335)
);

CKINVDCx6p67_ASAP7_75t_R g1336 ( 
.A(n_1119),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1150),
.Y(n_1337)
);

CKINVDCx11_ASAP7_75t_R g1338 ( 
.A(n_1119),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1304),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1236),
.B(n_1240),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1271),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1300),
.B(n_1310),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1274),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1249),
.B(n_1259),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1249),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1296),
.A2(n_1297),
.B(n_1308),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1234),
.A2(n_1315),
.B1(n_1313),
.B2(n_1318),
.Y(n_1347)
);

OAI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1239),
.A2(n_1333),
.B1(n_1335),
.B2(n_1324),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1242),
.B(n_1267),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1303),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1308),
.A2(n_1311),
.B(n_1302),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1298),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1309),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1301),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1231),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1311),
.A2(n_1302),
.B(n_1288),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1295),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1240),
.B(n_1238),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1306),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1292),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1305),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1295),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1230),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1295),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1242),
.B(n_1267),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1293),
.B(n_1246),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1278),
.A2(n_1232),
.B(n_1268),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1293),
.B(n_1288),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1312),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1246),
.B(n_1234),
.Y(n_1370)
);

BUFx12f_ASAP7_75t_L g1371 ( 
.A(n_1338),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1294),
.Y(n_1372)
);

BUFx12f_ASAP7_75t_L g1373 ( 
.A(n_1338),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1281),
.B(n_1260),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1281),
.A2(n_1277),
.B(n_1266),
.Y(n_1375)
);

NAND3xp33_ASAP7_75t_L g1376 ( 
.A(n_1313),
.B(n_1329),
.C(n_1318),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_R g1377 ( 
.A(n_1263),
.B(n_1265),
.Y(n_1377)
);

AOI21xp33_ASAP7_75t_L g1378 ( 
.A1(n_1324),
.A2(n_1315),
.B(n_1329),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1287),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1299),
.B(n_1307),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1277),
.A2(n_1266),
.B(n_1284),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1307),
.B(n_1243),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1253),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1252),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1251),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1273),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1255),
.B(n_1247),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1273),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1320),
.B(n_1290),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1248),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1255),
.A2(n_1291),
.B1(n_1235),
.B2(n_1283),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1261),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1280),
.B(n_1276),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1257),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1319),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1258),
.A2(n_1282),
.A3(n_1326),
.B(n_1327),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1330),
.A2(n_1332),
.B1(n_1264),
.B2(n_1285),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1275),
.A2(n_1321),
.B1(n_1250),
.B2(n_1334),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1252),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1321),
.A2(n_1270),
.B1(n_1275),
.B2(n_1334),
.Y(n_1400)
);

AOI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1323),
.A2(n_1328),
.B(n_1272),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1245),
.A2(n_1325),
.B1(n_1334),
.B2(n_1256),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1264),
.Y(n_1403)
);

OAI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1286),
.A2(n_1336),
.B1(n_1325),
.B2(n_1245),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1279),
.A2(n_1325),
.B(n_1245),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1254),
.B(n_1337),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1314),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1233),
.B(n_1286),
.Y(n_1408)
);

AOI221xp5_ASAP7_75t_L g1409 ( 
.A1(n_1376),
.A2(n_1237),
.B1(n_1262),
.B2(n_1331),
.C(n_1269),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1376),
.A2(n_1316),
.B(n_1269),
.C(n_1263),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1356),
.A2(n_1346),
.B(n_1351),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1405),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1378),
.A2(n_1316),
.B(n_1289),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1347),
.A2(n_1378),
.B(n_1348),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1342),
.B(n_1314),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1345),
.Y(n_1416)
);

OAI211xp5_ASAP7_75t_L g1417 ( 
.A1(n_1347),
.A2(n_1322),
.B(n_1317),
.C(n_1241),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1369),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1363),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_SL g1420 ( 
.A1(n_1348),
.A2(n_1358),
.B(n_1340),
.C(n_1404),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1387),
.B(n_1322),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1370),
.A2(n_1244),
.B1(n_1340),
.B2(n_1358),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1370),
.A2(n_1387),
.B1(n_1391),
.B2(n_1397),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1405),
.B(n_1354),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1342),
.B(n_1389),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_SL g1426 ( 
.A(n_1407),
.B(n_1371),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1403),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1391),
.A2(n_1381),
.B(n_1385),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1381),
.A2(n_1367),
.B(n_1397),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1381),
.A2(n_1349),
.B(n_1365),
.C(n_1379),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1398),
.A2(n_1357),
.B1(n_1364),
.B2(n_1400),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1351),
.A2(n_1356),
.B(n_1388),
.Y(n_1432)
);

OR2x6_ASAP7_75t_L g1433 ( 
.A(n_1375),
.B(n_1405),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1349),
.A2(n_1365),
.B(n_1379),
.C(n_1375),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1399),
.B(n_1396),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1396),
.B(n_1384),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1394),
.B(n_1395),
.Y(n_1437)
);

NAND4xp25_ASAP7_75t_L g1438 ( 
.A(n_1386),
.B(n_1402),
.C(n_1355),
.D(n_1393),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1349),
.A2(n_1365),
.B(n_1375),
.C(n_1366),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1374),
.B(n_1346),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1396),
.B(n_1384),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1395),
.B(n_1393),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1346),
.A2(n_1351),
.B(n_1356),
.Y(n_1443)
);

A2O1A1Ixp33_ASAP7_75t_L g1444 ( 
.A1(n_1366),
.A2(n_1374),
.B(n_1357),
.C(n_1364),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1396),
.B(n_1406),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1393),
.B(n_1392),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1366),
.A2(n_1374),
.B(n_1357),
.C(n_1364),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1361),
.A2(n_1367),
.B(n_1353),
.Y(n_1448)
);

AO32x1_ASAP7_75t_L g1449 ( 
.A1(n_1350),
.A2(n_1339),
.A3(n_1343),
.B1(n_1361),
.B2(n_1360),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1377),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1342),
.B(n_1382),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1392),
.B(n_1355),
.Y(n_1452)
);

AO21x2_ASAP7_75t_L g1453 ( 
.A1(n_1353),
.A2(n_1359),
.B(n_1339),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1404),
.A2(n_1400),
.B1(n_1402),
.B2(n_1398),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1372),
.A2(n_1362),
.B(n_1408),
.C(n_1390),
.Y(n_1455)
);

AOI221xp5_ASAP7_75t_L g1456 ( 
.A1(n_1372),
.A2(n_1382),
.B1(n_1362),
.B2(n_1380),
.C(n_1383),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1432),
.B(n_1368),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1453),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1451),
.B(n_1382),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1432),
.B(n_1440),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1419),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1418),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1416),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1440),
.B(n_1368),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1425),
.B(n_1368),
.Y(n_1465)
);

BUFx12f_ASAP7_75t_L g1466 ( 
.A(n_1450),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1412),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1414),
.A2(n_1380),
.B1(n_1362),
.B2(n_1373),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1424),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1445),
.B(n_1360),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1422),
.A2(n_1373),
.B1(n_1371),
.B2(n_1362),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1449),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1448),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1452),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1446),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1442),
.B(n_1439),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1433),
.B(n_1341),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_SL g1478 ( 
.A(n_1433),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1433),
.B(n_1344),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1453),
.Y(n_1480)
);

INVx6_ASAP7_75t_L g1481 ( 
.A(n_1466),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1469),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1463),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1473),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1476),
.B(n_1421),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1459),
.B(n_1411),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1459),
.B(n_1411),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1466),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1459),
.B(n_1411),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1473),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1479),
.B(n_1435),
.Y(n_1491)
);

AOI221xp5_ASAP7_75t_L g1492 ( 
.A1(n_1476),
.A2(n_1420),
.B1(n_1439),
.B2(n_1430),
.C(n_1434),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1474),
.B(n_1434),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1463),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1479),
.B(n_1443),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1464),
.B(n_1436),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1473),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1464),
.B(n_1441),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1464),
.B(n_1465),
.Y(n_1499)
);

OAI31xp33_ASAP7_75t_L g1500 ( 
.A1(n_1471),
.A2(n_1420),
.A3(n_1430),
.B(n_1417),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1468),
.A2(n_1423),
.B1(n_1422),
.B2(n_1444),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1465),
.B(n_1470),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1475),
.B(n_1437),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1468),
.A2(n_1428),
.B(n_1429),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1461),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1462),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1462),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1506),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1484),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1486),
.B(n_1460),
.Y(n_1510)
);

AND2x2_ASAP7_75t_SL g1511 ( 
.A(n_1492),
.B(n_1380),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1494),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1486),
.B(n_1460),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1486),
.B(n_1460),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1484),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1487),
.B(n_1472),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1506),
.B(n_1507),
.Y(n_1517)
);

NAND2x1p5_ASAP7_75t_L g1518 ( 
.A(n_1482),
.B(n_1467),
.Y(n_1518)
);

INVxp67_ASAP7_75t_SL g1519 ( 
.A(n_1494),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1484),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1484),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1490),
.Y(n_1522)
);

NOR2x1_ASAP7_75t_L g1523 ( 
.A(n_1488),
.B(n_1467),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1506),
.B(n_1472),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1490),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1492),
.A2(n_1421),
.B1(n_1471),
.B2(n_1409),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1482),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1497),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1507),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1489),
.B(n_1477),
.Y(n_1530)
);

INVx1_ASAP7_75t_SL g1531 ( 
.A(n_1482),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1507),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1499),
.B(n_1495),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1483),
.B(n_1472),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1505),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1499),
.B(n_1477),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1527),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1508),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1511),
.B(n_1485),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1508),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1527),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1527),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1527),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1527),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1511),
.B(n_1485),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1508),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1529),
.Y(n_1547)
);

NAND2xp33_ASAP7_75t_L g1548 ( 
.A(n_1526),
.B(n_1450),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1533),
.B(n_1499),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1529),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1534),
.B(n_1493),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1529),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1528),
.Y(n_1553)
);

OAI21xp33_ASAP7_75t_L g1554 ( 
.A1(n_1511),
.A2(n_1504),
.B(n_1501),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1534),
.B(n_1493),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1532),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1532),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1532),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1517),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1533),
.B(n_1496),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1517),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1517),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1511),
.A2(n_1501),
.B1(n_1504),
.B2(n_1454),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1511),
.B(n_1500),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1523),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1531),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1536),
.B(n_1503),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1535),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1533),
.B(n_1496),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1533),
.B(n_1496),
.Y(n_1570)
);

NAND4xp75_ASAP7_75t_L g1571 ( 
.A(n_1523),
.B(n_1500),
.C(n_1415),
.D(n_1413),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1535),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1534),
.B(n_1457),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1535),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1528),
.Y(n_1575)
);

AOI21xp33_ASAP7_75t_L g1576 ( 
.A1(n_1526),
.A2(n_1455),
.B(n_1431),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1523),
.B(n_1488),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1536),
.B(n_1498),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1551),
.B(n_1531),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1542),
.B(n_1531),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1578),
.B(n_1536),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1554),
.B(n_1536),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1539),
.B(n_1498),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1538),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1571),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1578),
.B(n_1530),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1538),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1566),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1545),
.B(n_1498),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1563),
.B(n_1502),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1551),
.B(n_1524),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1564),
.A2(n_1519),
.B(n_1410),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1540),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1555),
.B(n_1502),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1555),
.B(n_1524),
.Y(n_1595)
);

INVx3_ASAP7_75t_SL g1596 ( 
.A(n_1577),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1548),
.B(n_1371),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1542),
.B(n_1544),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1540),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1576),
.B(n_1502),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1566),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1544),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1560),
.B(n_1569),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1560),
.B(n_1530),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1567),
.B(n_1524),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1577),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1571),
.B(n_1537),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1546),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1537),
.B(n_1503),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1569),
.B(n_1570),
.Y(n_1610)
);

OAI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1565),
.A2(n_1481),
.B1(n_1457),
.B2(n_1488),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1541),
.B(n_1491),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1546),
.Y(n_1613)
);

NAND3xp33_ASAP7_75t_SL g1614 ( 
.A(n_1585),
.B(n_1377),
.C(n_1426),
.Y(n_1614)
);

OAI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1592),
.A2(n_1410),
.B1(n_1481),
.B2(n_1488),
.C(n_1565),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1587),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1587),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_1598),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1608),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1596),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1607),
.A2(n_1577),
.B(n_1519),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1588),
.B(n_1541),
.Y(n_1622)
);

OAI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1596),
.A2(n_1481),
.B1(n_1457),
.B2(n_1438),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1608),
.Y(n_1624)
);

OAI21xp33_ASAP7_75t_SL g1625 ( 
.A1(n_1582),
.A2(n_1606),
.B(n_1590),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1598),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1600),
.A2(n_1478),
.B1(n_1481),
.B2(n_1543),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1613),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1601),
.B(n_1543),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1597),
.A2(n_1573),
.B(n_1512),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_SL g1631 ( 
.A1(n_1606),
.A2(n_1415),
.B1(n_1512),
.B2(n_1352),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1613),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1601),
.A2(n_1481),
.B1(n_1456),
.B2(n_1573),
.C(n_1447),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1598),
.Y(n_1634)
);

OAI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1583),
.A2(n_1481),
.B1(n_1518),
.B2(n_1480),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1611),
.A2(n_1480),
.B(n_1458),
.C(n_1518),
.Y(n_1636)
);

OAI32xp33_ASAP7_75t_L g1637 ( 
.A1(n_1579),
.A2(n_1518),
.A3(n_1516),
.B1(n_1570),
.B2(n_1559),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1609),
.A2(n_1518),
.B(n_1458),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1616),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1614),
.B(n_1373),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1617),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1619),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1624),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1620),
.B(n_1603),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1615),
.A2(n_1602),
.B1(n_1612),
.B2(n_1589),
.Y(n_1645)
);

AOI21xp33_ASAP7_75t_L g1646 ( 
.A1(n_1625),
.A2(n_1602),
.B(n_1579),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1631),
.B(n_1603),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1615),
.A2(n_1591),
.B1(n_1595),
.B2(n_1481),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1628),
.Y(n_1649)
);

AOI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1621),
.A2(n_1637),
.B1(n_1623),
.B2(n_1633),
.C(n_1630),
.Y(n_1650)
);

AOI22x1_ASAP7_75t_L g1651 ( 
.A1(n_1621),
.A2(n_1580),
.B1(n_1466),
.B2(n_1595),
.Y(n_1651)
);

AOI222xp33_ASAP7_75t_L g1652 ( 
.A1(n_1633),
.A2(n_1622),
.B1(n_1638),
.B2(n_1629),
.C1(n_1635),
.C2(n_1632),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1634),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1626),
.B(n_1610),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1618),
.B(n_1610),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_L g1656 ( 
.A(n_1627),
.B(n_1634),
.C(n_1636),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1634),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1653),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1644),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1657),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1657),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1647),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1650),
.A2(n_1580),
.B(n_1584),
.Y(n_1663)
);

NOR2x1_ASAP7_75t_L g1664 ( 
.A(n_1640),
.B(n_1580),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1654),
.B(n_1594),
.Y(n_1665)
);

OAI22xp33_ASAP7_75t_SL g1666 ( 
.A1(n_1651),
.A2(n_1591),
.B1(n_1593),
.B2(n_1599),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1639),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1641),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1664),
.B(n_1655),
.Y(n_1669)
);

NAND3xp33_ASAP7_75t_SL g1670 ( 
.A(n_1662),
.B(n_1652),
.C(n_1663),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1660),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1666),
.B(n_1648),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1661),
.B(n_1645),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1659),
.B(n_1666),
.Y(n_1674)
);

NOR3xp33_ASAP7_75t_SL g1675 ( 
.A(n_1658),
.B(n_1656),
.C(n_1648),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1665),
.A2(n_1646),
.B1(n_1649),
.B2(n_1643),
.Y(n_1676)
);

NOR4xp25_ASAP7_75t_L g1677 ( 
.A(n_1667),
.B(n_1646),
.C(n_1642),
.D(n_1605),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1668),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1660),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1670),
.A2(n_1605),
.B(n_1553),
.C(n_1575),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_SL g1681 ( 
.A(n_1677),
.B(n_1604),
.C(n_1581),
.Y(n_1681)
);

AOI222xp33_ASAP7_75t_L g1682 ( 
.A1(n_1672),
.A2(n_1604),
.B1(n_1586),
.B2(n_1581),
.C1(n_1575),
.C2(n_1553),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1674),
.A2(n_1586),
.B1(n_1466),
.B2(n_1549),
.Y(n_1683)
);

NOR4xp75_ASAP7_75t_L g1684 ( 
.A(n_1673),
.B(n_1549),
.C(n_1510),
.D(n_1514),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1669),
.Y(n_1685)
);

OAI221xp5_ASAP7_75t_SL g1686 ( 
.A1(n_1683),
.A2(n_1676),
.B1(n_1671),
.B2(n_1679),
.C(n_1678),
.Y(n_1686)
);

OAI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1685),
.A2(n_1675),
.B1(n_1518),
.B2(n_1559),
.C(n_1562),
.Y(n_1687)
);

NOR4xp25_ASAP7_75t_L g1688 ( 
.A(n_1680),
.B(n_1675),
.C(n_1561),
.D(n_1562),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_SL g1689 ( 
.A1(n_1681),
.A2(n_1408),
.B1(n_1427),
.B2(n_1558),
.Y(n_1689)
);

AOI32xp33_ASAP7_75t_L g1690 ( 
.A1(n_1684),
.A2(n_1514),
.A3(n_1510),
.B1(n_1513),
.B2(n_1561),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1682),
.A2(n_1550),
.B(n_1547),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1689),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1686),
.Y(n_1693)
);

XNOR2xp5_ASAP7_75t_L g1694 ( 
.A(n_1688),
.B(n_1352),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1687),
.A2(n_1691),
.B1(n_1690),
.B2(n_1516),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1687),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1693),
.A2(n_1692),
.B1(n_1696),
.B2(n_1694),
.Y(n_1697)
);

OAI322xp33_ASAP7_75t_L g1698 ( 
.A1(n_1695),
.A2(n_1574),
.A3(n_1572),
.B1(n_1568),
.B2(n_1557),
.C1(n_1556),
.C2(n_1552),
.Y(n_1698)
);

AOI21xp33_ASAP7_75t_SL g1699 ( 
.A1(n_1695),
.A2(n_1550),
.B(n_1547),
.Y(n_1699)
);

OAI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1697),
.A2(n_1574),
.B1(n_1572),
.B2(n_1568),
.C(n_1557),
.Y(n_1700)
);

AO22x2_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1699),
.B1(n_1698),
.B2(n_1556),
.Y(n_1701)
);

OAI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1552),
.B1(n_1516),
.B2(n_1528),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1701),
.Y(n_1703)
);

NAND3xp33_ASAP7_75t_SL g1704 ( 
.A(n_1703),
.B(n_1516),
.C(n_1515),
.Y(n_1704)
);

AO22x2_ASAP7_75t_L g1705 ( 
.A1(n_1702),
.A2(n_1528),
.B1(n_1509),
.B2(n_1515),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1704),
.A2(n_1510),
.B1(n_1513),
.B2(n_1514),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1705),
.A2(n_1513),
.B(n_1510),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1706),
.B(n_1513),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1708),
.B(n_1707),
.Y(n_1709)
);

XNOR2xp5_ASAP7_75t_L g1710 ( 
.A(n_1709),
.B(n_1401),
.Y(n_1710)
);

AOI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1710),
.A2(n_1525),
.B1(n_1520),
.B2(n_1509),
.C(n_1521),
.Y(n_1711)
);

AOI211xp5_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1352),
.B(n_1514),
.C(n_1522),
.Y(n_1712)
);


endmodule