module fake_jpeg_18855_n_209 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_209);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_12),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_44),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_48),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_17),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_34),
.Y(n_57)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_43),
.B1(n_36),
.B2(n_45),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_23),
.B1(n_26),
.B2(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_53),
.B1(n_56),
.B2(n_63),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_26),
.B1(n_23),
.B2(n_39),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_16),
.B1(n_30),
.B2(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_0),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_71),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_21),
.B1(n_20),
.B2(n_25),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_64),
.B1(n_47),
.B2(n_46),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_19),
.B1(n_28),
.B2(n_24),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_34),
.B1(n_50),
.B2(n_27),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_17),
.C(n_28),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_44),
.B(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_12),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_78),
.Y(n_104)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_58),
.B(n_17),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_24),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_80),
.Y(n_123)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_11),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_69),
.B1(n_49),
.B2(n_4),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_8),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_88),
.Y(n_118)
);

INVx5_ASAP7_75t_SL g89 ( 
.A(n_68),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_14),
.Y(n_90)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_13),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_99),
.B1(n_102),
.B2(n_59),
.Y(n_106)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

CKINVDCx12_ASAP7_75t_R g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_0),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_98),
.Y(n_121)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_69),
.B(n_50),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_103),
.B1(n_18),
.B2(n_6),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_81),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_115),
.B1(n_102),
.B2(n_77),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_18),
.B1(n_27),
.B2(n_5),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_87),
.B1(n_89),
.B2(n_122),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_82),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_131),
.B1(n_138),
.B2(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_84),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_112),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_84),
.C(n_75),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_135),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_93),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_132),
.B(n_110),
.Y(n_142)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_122),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_80),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_116),
.B(n_107),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_107),
.C(n_112),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_108),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_98),
.B1(n_91),
.B2(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_114),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_120),
.B(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_149),
.Y(n_168)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_135),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_124),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_152),
.B(n_151),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_118),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_131),
.B1(n_133),
.B2(n_125),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_152),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_130),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_157),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_134),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_165),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_138),
.B1(n_134),
.B2(n_137),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_162),
.B1(n_120),
.B2(n_76),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_153),
.B(n_150),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_167),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_128),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_139),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_170),
.A2(n_156),
.B1(n_160),
.B2(n_114),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_163),
.B(n_164),
.C(n_165),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_171),
.B(n_180),
.Y(n_183)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_173),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_153),
.B1(n_150),
.B2(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_158),
.B(n_118),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_179),
.Y(n_185)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_114),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_174),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_187),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_5),
.B(n_6),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_178),
.B(n_7),
.Y(n_188)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_188),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_105),
.B(n_85),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_176),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_188),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_176),
.B1(n_113),
.B2(n_7),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_191),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_184),
.C(n_182),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_181),
.B1(n_186),
.B2(n_183),
.Y(n_201)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_194),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_199),
.B(n_183),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_203),
.A2(n_200),
.B(n_186),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_204),
.B(n_195),
.Y(n_207)
);

A2O1A1O1Ixp25_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_195),
.B(n_113),
.C(n_105),
.D(n_100),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_85),
.Y(n_209)
);


endmodule