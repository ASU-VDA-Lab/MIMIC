module fake_netlist_1_2905_n_13 (n_3, n_1, n_2, n_0, n_13);
input n_3;
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
BUFx10_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
NAND2xp33_ASAP7_75t_R g5 ( .A(n_2), .B(n_3), .Y(n_5) );
NOR2xp33_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .Y(n_6) );
BUFx10_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_7), .B(n_4), .Y(n_8) );
INVxp67_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
AOI221xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_8), .B1(n_7), .B2(n_4), .C(n_5), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
OAI22xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_12) );
AOI22xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_13) );
endmodule