module fake_jpeg_25587_n_167 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_28),
.Y(n_48)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_1),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_18),
.B1(n_28),
.B2(n_23),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_29),
.B1(n_27),
.B2(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_48),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_31),
.B1(n_25),
.B2(n_30),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_31),
.A2(n_30),
.B1(n_21),
.B2(n_27),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_19),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_58),
.B(n_61),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_62),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_54),
.B1(n_47),
.B2(n_51),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_46),
.B1(n_53),
.B2(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_66),
.B(n_71),
.Y(n_82)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_37),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_16),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_35),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_17),
.B1(n_20),
.B2(n_16),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_87),
.B(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_64),
.B1(n_74),
.B2(n_53),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_17),
.B1(n_20),
.B2(n_46),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_35),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_71),
.C(n_70),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_95),
.C(n_101),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_67),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_102),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_86),
.B1(n_80),
.B2(n_78),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_67),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_105),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_69),
.C(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_91),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_65),
.B1(n_64),
.B2(n_43),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_109),
.A2(n_85),
.B1(n_93),
.B2(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_110),
.B(n_112),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_116),
.B1(n_119),
.B2(n_121),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_122),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_99),
.B1(n_104),
.B2(n_106),
.Y(n_124)
);

NAND2x1_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_88),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_77),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_77),
.B(n_87),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_123),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_134),
.B1(n_22),
.B2(n_38),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_111),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_115),
.B1(n_34),
.B2(n_38),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_96),
.C(n_43),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_52),
.C(n_38),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_34),
.B1(n_43),
.B2(n_52),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_131),
.A2(n_124),
.B1(n_129),
.B2(n_126),
.Y(n_137)
);

OAI321xp33_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_113),
.A3(n_111),
.B1(n_121),
.B2(n_116),
.C(n_112),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_136),
.A2(n_125),
.B(n_133),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_140),
.B(n_142),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_143),
.Y(n_146)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_128),
.C(n_125),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_132),
.A2(n_2),
.B(n_3),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_22),
.B1(n_38),
.B2(n_9),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_3),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_145),
.B(n_149),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_150),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_141),
.C(n_139),
.Y(n_149)
);

AOI321xp33_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_130),
.A3(n_12),
.B1(n_11),
.B2(n_10),
.C(n_7),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_143),
.B1(n_140),
.B2(n_12),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_136),
.C(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_154),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_4),
.C(n_5),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_153),
.A2(n_147),
.B1(n_146),
.B2(n_6),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_158),
.C(n_152),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_4),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_5),
.C(n_6),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_162),
.B(n_163),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_4),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_162),
.A2(n_5),
.B(n_7),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_7),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_164),
.Y(n_167)
);


endmodule