module fake_jpeg_27297_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx8_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_0),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_14),
.Y(n_40)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_29),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_37),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_21),
.B1(n_22),
.B2(n_20),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_16),
.B1(n_11),
.B2(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_19),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_17),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_26),
.B1(n_28),
.B2(n_27),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_36),
.B1(n_28),
.B2(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_23),
.B1(n_22),
.B2(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_16),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

AND2x4_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_29),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_29),
.B(n_11),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_36),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_49),
.B1(n_44),
.B2(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_49),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_63),
.B(n_50),
.Y(n_66)
);

XNOR2x1_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_13),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_49),
.B(n_45),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_63),
.B(n_64),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_67),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_57),
.C(n_54),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_47),
.B1(n_43),
.B2(n_15),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_73),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_47),
.B1(n_43),
.B2(n_15),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_69),
.B(n_53),
.Y(n_76)
);

OAI322xp33_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_70),
.A3(n_13),
.B1(n_8),
.B2(n_10),
.C1(n_56),
.C2(n_7),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_75),
.B(n_77),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_73),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_SL g83 ( 
.A(n_80),
.B(n_59),
.C(n_68),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_84),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_87),
.B1(n_55),
.B2(n_13),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_78),
.C(n_77),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_55),
.C(n_2),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_91),
.A2(n_56),
.B(n_2),
.Y(n_96)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVxp33_ASAP7_75t_SL g95 ( 
.A(n_92),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_88),
.B1(n_79),
.B2(n_70),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_97),
.C(n_1),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_90),
.B(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_95),
.B(n_89),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_99),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_6),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_3),
.C(n_6),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_101),
.A2(n_102),
.B(n_7),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_74),
.Y(n_104)
);


endmodule