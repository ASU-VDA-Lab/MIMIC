module fake_ariane_1639_n_1197 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1197);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1197;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1137;
wire n_646;
wire n_1174;
wire n_640;
wire n_197;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_176;
wire n_404;
wire n_172;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_183;
wire n_469;
wire n_1046;
wire n_726;
wire n_479;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_1029;
wire n_205;
wire n_341;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_690;
wire n_416;
wire n_1180;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_528;
wire n_584;
wire n_424;
wire n_1154;
wire n_1166;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_940;
wire n_756;
wire n_466;
wire n_1016;
wire n_346;
wire n_1138;
wire n_214;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_1196;
wire n_670;
wire n_607;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_1181;
wire n_515;
wire n_379;
wire n_445;
wire n_807;
wire n_1131;
wire n_765;
wire n_1187;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1167;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_186;
wire n_801;
wire n_1184;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_754;
wire n_336;
wire n_731;
wire n_779;
wire n_903;
wire n_871;
wire n_315;
wire n_1073;
wire n_594;
wire n_1173;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_557;
wire n_405;
wire n_1107;
wire n_173;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_1134;
wire n_1185;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_721;
wire n_433;
wire n_600;
wire n_840;
wire n_481;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_839;
wire n_218;
wire n_928;
wire n_1099;
wire n_1153;
wire n_271;
wire n_507;
wire n_465;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_240;
wire n_369;
wire n_1192;
wire n_224;
wire n_894;
wire n_787;
wire n_1105;
wire n_547;
wire n_1195;
wire n_420;
wire n_562;
wire n_518;
wire n_604;
wire n_677;
wire n_614;
wire n_439;
wire n_1172;
wire n_478;
wire n_703;
wire n_222;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_1160;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_1080;
wire n_576;
wire n_843;
wire n_206;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_192;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_1188;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_233;
wire n_728;
wire n_957;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_685;
wire n_911;
wire n_321;
wire n_459;
wire n_221;
wire n_1136;
wire n_361;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_181;
wire n_1142;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_1140;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_262;
wire n_209;
wire n_743;
wire n_1194;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_747;
wire n_741;
wire n_847;
wire n_939;
wire n_1135;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_673;
wire n_452;
wire n_1114;
wire n_676;
wire n_178;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_1038;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_571;
wire n_680;
wire n_414;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_212;
wire n_1043;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_1193;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_171;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_1081;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_774;
wire n_407;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_1157;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_664;
wire n_629;
wire n_1075;
wire n_215;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_1182;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_991;
wire n_834;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_179;
wire n_1126;
wire n_395;
wire n_621;
wire n_1178;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_998;
wire n_999;
wire n_967;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_174;
wire n_275;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_1148;
wire n_751;
wire n_1027;
wire n_615;
wire n_1070;
wire n_204;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1139;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_1051;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_1102;
wire n_360;
wire n_1101;
wire n_975;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1189;
wire n_1124;
wire n_250;
wire n_932;
wire n_1183;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_815;
wire n_542;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1191;
wire n_1071;
wire n_484;
wire n_411;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_1164;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_191;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_211;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_934;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_8),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_163),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_110),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_64),
.Y(n_176)
);

INVxp33_ASAP7_75t_SL g177 ( 
.A(n_84),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_26),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_111),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_36),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_88),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_93),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_12),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_62),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_18),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_15),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_35),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_71),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_103),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_118),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_60),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_138),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_122),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_73),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_47),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_58),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_23),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_33),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_98),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_40),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_6),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_12),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_143),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_8),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_169),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_120),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_125),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_128),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_41),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_89),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_28),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_13),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_75),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_114),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_81),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_115),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_217),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_193),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_178),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_216),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_207),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_216),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_170),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_173),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_187),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_202),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_183),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_183),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_208),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_190),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_196),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_234),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_174),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_175),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_237),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_225),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

BUFx8_ASAP7_75t_SL g268 ( 
.A(n_243),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_230),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_248),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_233),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_231),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_241),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_228),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_238),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_245),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_238),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_240),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_242),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_242),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_247),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_244),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_251),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_235),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_235),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_243),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_234),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_234),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_243),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_268),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_260),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_268),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_253),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_260),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_274),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_254),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_288),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_267),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_262),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_262),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_288),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_272),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_258),
.Y(n_317)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_292),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_275),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_264),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_270),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_277),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_300),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_286),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_271),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_276),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_283),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_274),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_295),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_298),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_299),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_284),
.Y(n_344)
);

INVxp33_ASAP7_75t_SL g345 ( 
.A(n_287),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_295),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_337),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_337),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_322),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_344),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_305),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_344),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_308),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_308),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_321),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_338),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_309),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g359 ( 
.A(n_310),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_338),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_336),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_331),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_293),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_307),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_341),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_318),
.B(n_293),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_341),
.Y(n_368)
);

INVxp33_ASAP7_75t_SL g369 ( 
.A(n_315),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_347),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_315),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_347),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_311),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_312),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_318),
.B(n_294),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_345),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_345),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_306),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_302),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_303),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_302),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_323),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_313),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_313),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_257),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_352),
.B(n_327),
.Y(n_390)
);

OA21x2_ASAP7_75t_L g391 ( 
.A1(n_358),
.A2(n_317),
.B(n_309),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_348),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_381),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_360),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_375),
.A2(n_330),
.B1(n_332),
.B2(n_333),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_328),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_379),
.Y(n_398)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_385),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_374),
.Y(n_401)
);

OAI22x1_ASAP7_75t_R g402 ( 
.A1(n_366),
.A2(n_304),
.B1(n_301),
.B2(n_291),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_377),
.Y(n_403)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

BUFx8_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_314),
.Y(n_406)
);

NAND2xp33_ASAP7_75t_R g407 ( 
.A(n_371),
.B(n_257),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_383),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_370),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_349),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_356),
.B(n_263),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_351),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_364),
.A2(n_294),
.B1(n_263),
.B2(n_255),
.Y(n_415)
);

BUFx12f_ASAP7_75t_L g416 ( 
.A(n_380),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_372),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_378),
.B(n_314),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_363),
.B(n_316),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_362),
.B(n_282),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_354),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_355),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_353),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_371),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_353),
.Y(n_426)
);

AND2x6_ASAP7_75t_L g427 ( 
.A(n_359),
.B(n_334),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_376),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_376),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_382),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_380),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_359),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_382),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_369),
.B(n_282),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_369),
.B(n_282),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_357),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_385),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_350),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_367),
.B(n_296),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_348),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_370),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_358),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_358),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_350),
.Y(n_447)
);

AND2x6_ASAP7_75t_L g448 ( 
.A(n_381),
.B(n_335),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_350),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_348),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_350),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_350),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_L g453 ( 
.A(n_348),
.B(n_282),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_350),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_358),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_370),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_367),
.A2(n_282),
.B1(n_343),
.B2(n_342),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_381),
.Y(n_458)
);

NOR2x1_ASAP7_75t_L g459 ( 
.A(n_361),
.B(n_339),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_350),
.B(n_326),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_357),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_388),
.B(n_265),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_419),
.B(n_340),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_387),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_419),
.B(n_346),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_387),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_440),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_399),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_442),
.B(n_413),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_445),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_399),
.B(n_303),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_409),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_401),
.B(n_403),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_446),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_394),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_403),
.B(n_256),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_394),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_408),
.B(n_259),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_408),
.B(n_273),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_409),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_458),
.Y(n_485)
);

OR2x6_ASAP7_75t_L g486 ( 
.A(n_400),
.B(n_320),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_458),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_437),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_399),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_398),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_391),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_437),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_398),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_399),
.B(n_404),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_441),
.B(n_320),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_447),
.Y(n_496)
);

BUFx8_ASAP7_75t_L g497 ( 
.A(n_416),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_404),
.B(n_320),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_415),
.B(n_291),
.Y(n_499)
);

AND2x2_ASAP7_75t_SL g500 ( 
.A(n_453),
.B(n_199),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_444),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_497),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_497),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_497),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_467),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_497),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_501),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_462),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_475),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_404),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_496),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_475),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_488),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_488),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_496),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_492),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_492),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_469),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_468),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_483),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_467),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_490),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_490),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_468),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_499),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_493),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_484),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_476),
.B(n_418),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_489),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_489),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_494),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_494),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_472),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_494),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_489),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_471),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_493),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_471),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_471),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_500),
.B(n_435),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_471),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_536),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_511),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_509),
.B(n_476),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_505),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_515),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_522),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_541),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_508),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_510),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_505),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_523),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_538),
.Y(n_553)
);

INVxp33_ASAP7_75t_L g554 ( 
.A(n_528),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_521),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_512),
.B(n_444),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_521),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_540),
.B(n_500),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_525),
.A2(n_301),
.B1(n_500),
.B2(n_434),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_526),
.B(n_456),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_513),
.B(n_456),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_533),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_537),
.B(n_464),
.Y(n_563)
);

AND2x2_ASAP7_75t_SL g564 ( 
.A(n_510),
.B(n_453),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_533),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_514),
.B(n_436),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_510),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_535),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_507),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_539),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_516),
.B(n_463),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_517),
.B(n_465),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_524),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_531),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_532),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_535),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_534),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_529),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_529),
.B(n_411),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_519),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_530),
.Y(n_581)
);

BUFx10_ASAP7_75t_L g582 ( 
.A(n_502),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_530),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_527),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_518),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_520),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_503),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_525),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_504),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_506),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_511),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_509),
.B(n_449),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_511),
.Y(n_593)
);

AND2x6_ASAP7_75t_L g594 ( 
.A(n_510),
.B(n_491),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_505),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_509),
.B(n_451),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_510),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_505),
.Y(n_598)
);

INVxp33_ASAP7_75t_L g599 ( 
.A(n_528),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_505),
.Y(n_600)
);

AND3x2_ASAP7_75t_L g601 ( 
.A(n_510),
.B(n_395),
.C(n_389),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_536),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_511),
.B(n_464),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_536),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_511),
.B(n_466),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_527),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_535),
.Y(n_607)
);

BUFx10_ASAP7_75t_L g608 ( 
.A(n_502),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_511),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_511),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_508),
.B(n_443),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_510),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_511),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_540),
.B(n_471),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_508),
.B(n_443),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_509),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_511),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_511),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_535),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_510),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_573),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_543),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_550),
.Y(n_623)
);

INVx8_ASAP7_75t_L g624 ( 
.A(n_549),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_620),
.B(n_498),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_579),
.B(n_411),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_546),
.Y(n_627)
);

BUFx4f_ASAP7_75t_L g628 ( 
.A(n_587),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_587),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_549),
.B(n_392),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_547),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_578),
.B(n_434),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_583),
.B(n_404),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_552),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_611),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_550),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_594),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_591),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_615),
.B(n_392),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_593),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_573),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_579),
.B(n_411),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_578),
.B(n_425),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_616),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_609),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_610),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_559),
.A2(n_482),
.B1(n_480),
.B2(n_410),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_560),
.B(n_466),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_573),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_606),
.B(n_393),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_583),
.B(n_485),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_586),
.B(n_393),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_571),
.B(n_450),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_567),
.B(n_485),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_603),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_568),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_567),
.B(n_485),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_613),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_617),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_618),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_594),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_587),
.Y(n_662)
);

INVx6_ASAP7_75t_L g663 ( 
.A(n_582),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_542),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_603),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_587),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_572),
.A2(n_304),
.B1(n_425),
.B2(n_281),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_582),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_550),
.Y(n_669)
);

INVx4_ASAP7_75t_SL g670 ( 
.A(n_594),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_556),
.B(n_450),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_542),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_605),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_605),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_582),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_608),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_560),
.B(n_421),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_563),
.Y(n_678)
);

BUFx4f_ASAP7_75t_L g679 ( 
.A(n_584),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_581),
.B(n_426),
.Y(n_680)
);

BUFx4f_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_563),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_569),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_542),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_545),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_561),
.B(n_422),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_620),
.B(n_498),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_568),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_592),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_596),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_588),
.B(n_422),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_588),
.B(n_426),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_548),
.B(n_411),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_545),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_551),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_550),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_553),
.B(n_438),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_608),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_553),
.B(n_438),
.Y(n_699)
);

AND2x6_ASAP7_75t_L g700 ( 
.A(n_597),
.B(n_498),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_602),
.B(n_412),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_551),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_555),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_555),
.Y(n_704)
);

AND2x6_ASAP7_75t_L g705 ( 
.A(n_597),
.B(n_498),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_663),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_686),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_631),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_631),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_622),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_623),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_670),
.B(n_602),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_627),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_689),
.B(n_690),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_665),
.B(n_580),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_670),
.B(n_604),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_647),
.A2(n_407),
.B1(n_558),
.B2(n_427),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_635),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_638),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_624),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_634),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_673),
.B(n_570),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_702),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_640),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_621),
.B(n_604),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_645),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_678),
.B(n_570),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_664),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_623),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_624),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_646),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_653),
.A2(n_407),
.B1(n_558),
.B2(n_427),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_658),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_637),
.B(n_594),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_659),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_682),
.B(n_544),
.Y(n_736)
);

OAI221xp5_ASAP7_75t_L g737 ( 
.A1(n_667),
.A2(n_429),
.B1(n_421),
.B2(n_396),
.C(n_428),
.Y(n_737)
);

NOR2x1p5_ASAP7_75t_L g738 ( 
.A(n_676),
.B(n_585),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_621),
.B(n_641),
.Y(n_739)
);

AND2x6_ASAP7_75t_L g740 ( 
.A(n_637),
.B(n_597),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_688),
.Y(n_741)
);

AO22x2_ASAP7_75t_L g742 ( 
.A1(n_694),
.A2(n_562),
.B1(n_565),
.B2(n_557),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_641),
.B(n_649),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_637),
.B(n_661),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_688),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_671),
.A2(n_427),
.B1(n_564),
.B2(n_566),
.Y(n_746)
);

NAND2x1p5_ASAP7_75t_L g747 ( 
.A(n_628),
.B(n_681),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_660),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_683),
.B(n_576),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_679),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_655),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_674),
.Y(n_752)
);

INVx4_ASAP7_75t_SL g753 ( 
.A(n_663),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_648),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_694),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_695),
.Y(n_756)
);

NAND3x1_ASAP7_75t_L g757 ( 
.A(n_697),
.B(n_590),
.C(n_589),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_695),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_685),
.Y(n_759)
);

NAND3x1_ASAP7_75t_L g760 ( 
.A(n_699),
.B(n_575),
.C(n_574),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_703),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_656),
.B(n_644),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_623),
.Y(n_763)
);

AO22x2_ASAP7_75t_L g764 ( 
.A1(n_704),
.A2(n_562),
.B1(n_565),
.B2(n_557),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_677),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_672),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_675),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_656),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_632),
.B(n_585),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_691),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_661),
.B(n_594),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_684),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_661),
.B(n_594),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_636),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_643),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_692),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_680),
.B(n_701),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_636),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_636),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_693),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_L g781 ( 
.A(n_737),
.B(n_566),
.C(n_626),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_754),
.B(n_662),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_717),
.A2(n_599),
.B1(n_554),
.B2(n_410),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_708),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_724),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_726),
.B(n_614),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_762),
.B(n_666),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_707),
.B(n_668),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_732),
.A2(n_639),
.B(n_652),
.C(n_650),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_718),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_780),
.B(n_614),
.C(n_577),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_733),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_706),
.B(n_698),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_757),
.B(n_412),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_766),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_750),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_765),
.B(n_629),
.Y(n_797)
);

AND2x6_ASAP7_75t_SL g798 ( 
.A(n_714),
.B(n_630),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_770),
.B(n_720),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_735),
.B(n_736),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_721),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_722),
.B(n_576),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_727),
.B(n_568),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_710),
.B(n_607),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_764),
.Y(n_805)
);

O2A1O1Ixp5_ASAP7_75t_L g806 ( 
.A1(n_725),
.A2(n_642),
.B(n_633),
.C(n_619),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_710),
.B(n_607),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_709),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_712),
.B(n_633),
.Y(n_809)
);

AND2x4_ASAP7_75t_SL g810 ( 
.A(n_712),
.B(n_608),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_766),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_730),
.B(n_412),
.Y(n_812)
);

INVx5_ASAP7_75t_L g813 ( 
.A(n_740),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_713),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_777),
.B(n_607),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_767),
.B(n_412),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_719),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_731),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_734),
.B(n_669),
.Y(n_819)
);

NOR2xp67_ASAP7_75t_L g820 ( 
.A(n_768),
.B(n_772),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_775),
.B(n_669),
.Y(n_821)
);

INVx4_ASAP7_75t_L g822 ( 
.A(n_753),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_747),
.B(n_414),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_L g824 ( 
.A(n_760),
.B(n_414),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_772),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_739),
.A2(n_564),
.B(n_651),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_764),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_753),
.B(n_414),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_716),
.B(n_669),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_738),
.B(n_651),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_748),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_746),
.B(n_414),
.Y(n_832)
);

BUFx4_ASAP7_75t_L g833 ( 
.A(n_778),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_716),
.B(n_696),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_776),
.B(n_619),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_749),
.B(n_619),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_715),
.B(n_554),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_SL g838 ( 
.A(n_740),
.B(n_696),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_769),
.B(n_599),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_728),
.B(n_696),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_751),
.B(n_601),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_752),
.B(n_778),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_723),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_742),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_759),
.B(n_654),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_755),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_741),
.B(n_423),
.Y(n_847)
);

O2A1O1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_743),
.A2(n_429),
.B(n_432),
.C(n_433),
.Y(n_848)
);

AND2x4_ASAP7_75t_SL g849 ( 
.A(n_711),
.B(n_597),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_741),
.B(n_424),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_761),
.B(n_756),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_758),
.B(n_654),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_779),
.B(n_657),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_734),
.B(n_771),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_742),
.Y(n_855)
);

NAND2x1_ASAP7_75t_L g856 ( 
.A(n_745),
.B(n_657),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_745),
.B(n_595),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_771),
.A2(n_410),
.B1(n_400),
.B2(n_405),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_773),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_711),
.Y(n_860)
);

AND2x2_ASAP7_75t_SL g861 ( 
.A(n_773),
.B(n_612),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_844),
.Y(n_862)
);

BUFx4f_ASAP7_75t_L g863 ( 
.A(n_796),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_846),
.B(n_711),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_784),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_808),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_851),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_822),
.Y(n_868)
);

BUFx12f_ASAP7_75t_L g869 ( 
.A(n_790),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_814),
.B(n_729),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_836),
.B(n_729),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_836),
.B(n_729),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_781),
.A2(n_410),
.B1(n_400),
.B2(n_405),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_796),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_813),
.B(n_763),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_817),
.B(n_763),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_794),
.A2(n_423),
.B(n_402),
.C(n_744),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_818),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_824),
.A2(n_214),
.B(n_209),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_832),
.A2(n_783),
.B1(n_841),
.B2(n_791),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_796),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_813),
.B(n_763),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_855),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_831),
.B(n_774),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_813),
.B(n_774),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_SL g886 ( 
.A1(n_805),
.A2(n_740),
.B1(n_744),
.B2(n_423),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_822),
.B(n_774),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_800),
.B(n_740),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_786),
.B(n_595),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_795),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_827),
.A2(n_400),
.B1(n_405),
.B2(n_423),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_786),
.B(n_598),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_798),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_785),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_792),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_842),
.Y(n_896)
);

NOR2x2_ASAP7_75t_L g897 ( 
.A(n_798),
.B(n_416),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_802),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_799),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_789),
.A2(n_620),
.B1(n_612),
.B2(n_461),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_801),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_815),
.B(n_598),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_804),
.B(n_600),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_843),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_787),
.B(n_417),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_835),
.B(n_600),
.Y(n_906)
);

OAI21xp33_ASAP7_75t_SL g907 ( 
.A1(n_820),
.A2(n_431),
.B(n_433),
.Y(n_907)
);

NAND3xp33_ASAP7_75t_L g908 ( 
.A(n_791),
.B(n_424),
.C(n_430),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_839),
.A2(n_473),
.B1(n_477),
.B2(n_472),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_857),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_806),
.A2(n_620),
.B(n_612),
.Y(n_911)
);

OR2x6_ASAP7_75t_L g912 ( 
.A(n_826),
.B(n_612),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_858),
.A2(n_477),
.B1(n_478),
.B2(n_473),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_833),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_821),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_795),
.B(n_424),
.Y(n_916)
);

O2A1O1Ixp5_ASAP7_75t_L g917 ( 
.A1(n_788),
.A2(n_431),
.B(n_479),
.C(n_470),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_847),
.Y(n_918)
);

AOI21x1_ASAP7_75t_L g919 ( 
.A1(n_890),
.A2(n_850),
.B(n_782),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_900),
.A2(n_809),
.B(n_829),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_896),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_893),
.A2(n_828),
.B(n_823),
.C(n_848),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_914),
.B(n_811),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_900),
.A2(n_907),
.B(n_877),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_908),
.A2(n_834),
.B(n_856),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_880),
.A2(n_845),
.B1(n_861),
.B2(n_853),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_L g927 ( 
.A(n_910),
.B(n_807),
.C(n_803),
.Y(n_927)
);

AOI21x1_ASAP7_75t_L g928 ( 
.A1(n_905),
.A2(n_860),
.B(n_857),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_869),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_867),
.B(n_837),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_879),
.A2(n_838),
.B(n_854),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_879),
.A2(n_816),
.B(n_812),
.C(n_830),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_868),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_912),
.B(n_854),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_918),
.B(n_811),
.Y(n_935)
);

AOI21x1_ASAP7_75t_L g936 ( 
.A1(n_916),
.A2(n_797),
.B(n_840),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_898),
.B(n_825),
.Y(n_937)
);

OAI22x1_ASAP7_75t_L g938 ( 
.A1(n_897),
.A2(n_793),
.B1(n_859),
.B2(n_819),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_917),
.A2(n_825),
.B(n_852),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_878),
.B(n_810),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_865),
.B(n_819),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_912),
.A2(n_838),
.B(n_849),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_866),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_874),
.B(n_918),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_903),
.B(n_424),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_912),
.A2(n_431),
.B(n_430),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_899),
.B(n_868),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_874),
.B(n_430),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_862),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_903),
.B(n_430),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_874),
.B(n_439),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_906),
.B(n_218),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_889),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_863),
.A2(n_486),
.B(n_418),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_870),
.B(n_625),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_864),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_889),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_915),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_863),
.A2(n_486),
.B(n_418),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_870),
.B(n_625),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_876),
.B(n_625),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_876),
.A2(n_177),
.B(n_420),
.C(n_213),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_884),
.B(n_687),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_873),
.A2(n_911),
.B(n_888),
.C(n_881),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_871),
.A2(n_457),
.B1(n_479),
.B2(n_470),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_892),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_892),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_918),
.B(n_487),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_887),
.A2(n_486),
.B(n_474),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_875),
.A2(n_885),
.B(n_882),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_884),
.B(n_687),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_864),
.A2(n_486),
.B(n_474),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_902),
.B(n_487),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_891),
.A2(n_176),
.B(n_474),
.C(n_459),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_894),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_872),
.B(n_687),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_883),
.B(n_700),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_895),
.B(n_0),
.Y(n_978)
);

OAI21xp33_ASAP7_75t_L g979 ( 
.A1(n_886),
.A2(n_454),
.B(n_452),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_913),
.A2(n_474),
.B(n_406),
.C(n_180),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_901),
.B(n_904),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_909),
.B(n_700),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_869),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_900),
.A2(n_427),
.B(n_700),
.Y(n_984)
);

NOR2xp67_ASAP7_75t_L g985 ( 
.A(n_938),
.B(n_0),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_921),
.B(n_1),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_929),
.B(n_1),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_924),
.A2(n_406),
.B(n_180),
.C(n_495),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_978),
.A2(n_926),
.B1(n_984),
.B2(n_979),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_983),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_934),
.B(n_970),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_943),
.B(n_2),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_984),
.A2(n_427),
.B1(n_705),
.B2(n_406),
.Y(n_993)
);

NAND2xp33_ASAP7_75t_SL g994 ( 
.A(n_923),
.B(n_2),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_930),
.B(n_3),
.Y(n_995)
);

INVxp67_ASAP7_75t_L g996 ( 
.A(n_947),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_945),
.A2(n_705),
.B1(n_495),
.B2(n_448),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_964),
.A2(n_920),
.B(n_925),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_934),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_952),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_SL g1001 ( 
.A(n_931),
.B(n_705),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_956),
.B(n_3),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_932),
.A2(n_479),
.B1(n_481),
.B2(n_470),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_975),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_936),
.Y(n_1005)
);

BUFx4f_ASAP7_75t_L g1006 ( 
.A(n_1000),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_998),
.A2(n_962),
.B(n_922),
.C(n_946),
.Y(n_1007)
);

AO32x2_ASAP7_75t_L g1008 ( 
.A1(n_1003),
.A2(n_956),
.A3(n_958),
.B1(n_965),
.B2(n_928),
.Y(n_1008)
);

BUFx2_ASAP7_75t_SL g1009 ( 
.A(n_985),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_1002),
.B(n_950),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_996),
.B(n_933),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_SL g1012 ( 
.A1(n_987),
.A2(n_933),
.B(n_948),
.C(n_939),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_990),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_1000),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_999),
.B(n_935),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_992),
.B(n_951),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_989),
.A2(n_927),
.B1(n_940),
.B2(n_944),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_999),
.A2(n_919),
.B(n_937),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_1000),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_991),
.B(n_942),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_1004),
.Y(n_1021)
);

NOR2x1_ASAP7_75t_L g1022 ( 
.A(n_986),
.B(n_941),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_1005),
.A2(n_949),
.B(n_953),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_995),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_997),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_SL g1026 ( 
.A(n_994),
.B(n_968),
.C(n_960),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_988),
.B(n_957),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_1001),
.A2(n_974),
.B(n_980),
.C(n_967),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_993),
.A2(n_966),
.B(n_973),
.C(n_954),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_998),
.A2(n_961),
.B(n_963),
.C(n_955),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_1013),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_1013),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1024),
.B(n_971),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1021),
.Y(n_1034)
);

AOI222xp33_ASAP7_75t_L g1035 ( 
.A1(n_1007),
.A2(n_982),
.B1(n_981),
.B2(n_977),
.C1(n_180),
.C2(n_460),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1014),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_1006),
.B(n_976),
.Y(n_1037)
);

AO21x2_ASAP7_75t_L g1038 ( 
.A1(n_1036),
.A2(n_1020),
.B(n_1012),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_1037),
.A2(n_1026),
.B1(n_1019),
.B2(n_1017),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_1038),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_1039),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_1038),
.A2(n_1009),
.B1(n_1035),
.B2(n_1014),
.Y(n_1042)
);

AOI22x1_ASAP7_75t_L g1043 ( 
.A1(n_1040),
.A2(n_1031),
.B1(n_1032),
.B2(n_1011),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1042),
.A2(n_1032),
.B(n_1018),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_1041),
.B(n_1031),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_SL g1046 ( 
.A1(n_1044),
.A2(n_1045),
.B1(n_1043),
.B2(n_1034),
.Y(n_1046)
);

INVx5_ASAP7_75t_L g1047 ( 
.A(n_1045),
.Y(n_1047)
);

OA21x2_ASAP7_75t_L g1048 ( 
.A1(n_1046),
.A2(n_1023),
.B(n_1011),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_1047),
.Y(n_1049)
);

BUFx10_ASAP7_75t_L g1050 ( 
.A(n_1049),
.Y(n_1050)
);

INVxp67_ASAP7_75t_SL g1051 ( 
.A(n_1048),
.Y(n_1051)
);

NAND2x1p5_ASAP7_75t_L g1052 ( 
.A(n_1050),
.B(n_1031),
.Y(n_1052)
);

CKINVDCx6p67_ASAP7_75t_R g1053 ( 
.A(n_1051),
.Y(n_1053)
);

OA21x2_ASAP7_75t_L g1054 ( 
.A1(n_1053),
.A2(n_1033),
.B(n_1016),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1052),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_1054),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1054),
.B(n_1055),
.Y(n_1057)
);

AOI21xp33_ASAP7_75t_SL g1058 ( 
.A1(n_1057),
.A2(n_1056),
.B(n_1035),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1056),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_1057),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1060),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_1059),
.B(n_1015),
.Y(n_1062)
);

INVxp67_ASAP7_75t_SL g1063 ( 
.A(n_1058),
.Y(n_1063)
);

AND2x2_ASAP7_75t_SL g1064 ( 
.A(n_1061),
.B(n_1027),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1063),
.B(n_1022),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1064),
.B(n_1062),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1065),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1066),
.B(n_1008),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1067),
.B(n_1008),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_1069),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_1068),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1070),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1071),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1072),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_1073),
.B(n_1010),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1075),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1074),
.B(n_4),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1074),
.B(n_4),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_1076),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1077),
.B(n_1008),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1078),
.Y(n_1081)
);

XNOR2xp5_ASAP7_75t_L g1082 ( 
.A(n_1079),
.B(n_5),
.Y(n_1082)
);

XOR2x2_ASAP7_75t_L g1083 ( 
.A(n_1081),
.B(n_5),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1083),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_1082),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1084),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1085),
.B(n_1080),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1086),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1087),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1089),
.Y(n_1090)
);

AOI21xp33_ASAP7_75t_SL g1091 ( 
.A1(n_1088),
.A2(n_181),
.B(n_179),
.Y(n_1091)
);

OAI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1090),
.A2(n_1091),
.B1(n_180),
.B2(n_188),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1090),
.B(n_6),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1093),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1092),
.B(n_7),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1092),
.B(n_7),
.Y(n_1096)
);

NOR3xp33_ASAP7_75t_L g1097 ( 
.A(n_1094),
.B(n_191),
.C(n_184),
.Y(n_1097)
);

NAND4xp25_ASAP7_75t_L g1098 ( 
.A(n_1096),
.B(n_1030),
.C(n_1025),
.D(n_11),
.Y(n_1098)
);

AOI321xp33_ASAP7_75t_L g1099 ( 
.A1(n_1095),
.A2(n_1029),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.C(n_14),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_1097),
.A2(n_192),
.B(n_224),
.C(n_195),
.Y(n_1100)
);

AO22x1_ASAP7_75t_L g1101 ( 
.A1(n_1099),
.A2(n_206),
.B1(n_197),
.B2(n_200),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1101),
.Y(n_1102)
);

NAND4xp25_ASAP7_75t_L g1103 ( 
.A(n_1100),
.B(n_1098),
.C(n_10),
.D(n_14),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1102),
.A2(n_204),
.B(n_201),
.Y(n_1104)
);

NOR2x1_ASAP7_75t_L g1105 ( 
.A(n_1103),
.B(n_194),
.Y(n_1105)
);

AOI221xp5_ASAP7_75t_L g1106 ( 
.A1(n_1104),
.A2(n_215),
.B1(n_223),
.B2(n_222),
.C(n_221),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1105),
.A2(n_194),
.B1(n_205),
.B2(n_211),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1107),
.B(n_194),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1106),
.A2(n_194),
.B1(n_212),
.B2(n_959),
.Y(n_1109)
);

NAND4xp25_ASAP7_75t_L g1110 ( 
.A(n_1108),
.B(n_1109),
.C(n_194),
.D(n_16),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_1108),
.B(n_981),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_1110),
.B(n_194),
.Y(n_1112)
);

NAND4xp75_ASAP7_75t_L g1113 ( 
.A(n_1111),
.B(n_390),
.C(n_397),
.D(n_194),
.Y(n_1113)
);

NOR2x1_ASAP7_75t_L g1114 ( 
.A(n_1110),
.B(n_9),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_1112),
.B(n_9),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1114),
.B(n_15),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1113),
.A2(n_1028),
.B1(n_17),
.B2(n_18),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1116),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1115),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1119),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1118),
.B(n_1117),
.Y(n_1121)
);

AOI211xp5_ASAP7_75t_L g1122 ( 
.A1(n_1120),
.A2(n_16),
.B(n_17),
.C(n_19),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_SL g1123 ( 
.A(n_1121),
.B(n_19),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_1123),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_SL g1125 ( 
.A1(n_1122),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1124),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1125),
.A2(n_20),
.B(n_21),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_1126),
.B(n_22),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1127),
.B(n_23),
.Y(n_1129)
);

XOR2x1_ASAP7_75t_L g1130 ( 
.A(n_1129),
.B(n_24),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1128),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1128),
.Y(n_1132)
);

XOR2x1_ASAP7_75t_L g1133 ( 
.A(n_1131),
.B(n_24),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_1132),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1130),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_SL g1136 ( 
.A1(n_1134),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1133),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1137),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1136),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1138),
.B(n_1135),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1139),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1140),
.Y(n_1142)
);

OAI332xp33_ASAP7_75t_L g1143 ( 
.A1(n_1141),
.A2(n_29),
.A3(n_30),
.B1(n_31),
.B2(n_32),
.B3(n_34),
.C1(n_37),
.C2(n_38),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1142),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1143),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1144),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1145),
.Y(n_1147)
);

INVxp33_ASAP7_75t_L g1148 ( 
.A(n_1144),
.Y(n_1148)
);

OAI331xp33_ASAP7_75t_L g1149 ( 
.A1(n_1148),
.A2(n_48),
.A3(n_49),
.B1(n_50),
.B2(n_51),
.B3(n_52),
.C1(n_53),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1147),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1146),
.A2(n_54),
.B(n_55),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1148),
.B(n_56),
.Y(n_1152)
);

OAI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1150),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1149),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1152),
.A2(n_68),
.B(n_70),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1151),
.A2(n_72),
.B(n_74),
.Y(n_1156)
);

AOI222xp33_ASAP7_75t_L g1157 ( 
.A1(n_1154),
.A2(n_1153),
.B1(n_1155),
.B2(n_1156),
.C1(n_79),
.C2(n_80),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1155),
.A2(n_76),
.B(n_77),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1155),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1155),
.A2(n_78),
.B(n_82),
.Y(n_1160)
);

OAI221xp5_ASAP7_75t_L g1161 ( 
.A1(n_1155),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.C(n_87),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_SL g1162 ( 
.A1(n_1155),
.A2(n_90),
.B(n_91),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1155),
.A2(n_92),
.B(n_94),
.Y(n_1163)
);

AOI222xp33_ASAP7_75t_L g1164 ( 
.A1(n_1154),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.C1(n_99),
.C2(n_100),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1155),
.Y(n_1165)
);

AOI221xp5_ASAP7_75t_L g1166 ( 
.A1(n_1155),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.C(n_106),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1155),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_1167)
);

XOR2xp5_ASAP7_75t_L g1168 ( 
.A(n_1155),
.B(n_112),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1159),
.A2(n_113),
.B(n_116),
.C(n_117),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1165),
.B(n_119),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1164),
.Y(n_1171)
);

AOI221xp5_ASAP7_75t_L g1172 ( 
.A1(n_1162),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.C(n_126),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1160),
.A2(n_969),
.B(n_129),
.Y(n_1173)
);

INVxp67_ASAP7_75t_SL g1174 ( 
.A(n_1157),
.Y(n_1174)
);

INVxp67_ASAP7_75t_L g1175 ( 
.A(n_1166),
.Y(n_1175)
);

OA21x2_ASAP7_75t_L g1176 ( 
.A1(n_1161),
.A2(n_1163),
.B(n_1158),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1168),
.A2(n_127),
.B(n_130),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1175),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1174),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1176),
.B(n_1167),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1171),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1170),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_1172),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1169),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1178),
.Y(n_1185)
);

AOI222xp33_ASAP7_75t_L g1186 ( 
.A1(n_1179),
.A2(n_1177),
.B1(n_1173),
.B2(n_139),
.C1(n_140),
.C2(n_141),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1180),
.A2(n_135),
.B(n_137),
.Y(n_1187)
);

AO21x2_ASAP7_75t_L g1188 ( 
.A1(n_1183),
.A2(n_142),
.B(n_144),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_1185),
.A2(n_1181),
.B(n_1182),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_SL g1190 ( 
.A1(n_1189),
.A2(n_1187),
.B1(n_1188),
.B2(n_1186),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1190),
.A2(n_1184),
.B1(n_146),
.B2(n_148),
.Y(n_1191)
);

NAND3xp33_ASAP7_75t_L g1192 ( 
.A(n_1191),
.B(n_145),
.C(n_149),
.Y(n_1192)
);

OAI221xp5_ASAP7_75t_L g1193 ( 
.A1(n_1192),
.A2(n_150),
.B1(n_151),
.B2(n_154),
.C(n_155),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1193),
.A2(n_972),
.B(n_158),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1194),
.A2(n_156),
.B(n_159),
.Y(n_1195)
);

AOI211xp5_ASAP7_75t_L g1196 ( 
.A1(n_1195),
.A2(n_160),
.B(n_162),
.C(n_164),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1196),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_1197)
);


endmodule