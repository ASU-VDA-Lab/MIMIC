module fake_aes_8466_n_735 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_735);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_735;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_17), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_6), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_58), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_12), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_7), .Y(n_84) );
INVxp67_ASAP7_75t_L g85 ( .A(n_33), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_9), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_55), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_54), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_14), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_31), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_69), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_38), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_74), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_3), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_8), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_43), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_19), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_22), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_78), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_27), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_51), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_75), .Y(n_102) );
CKINVDCx14_ASAP7_75t_R g103 ( .A(n_39), .Y(n_103) );
BUFx2_ASAP7_75t_L g104 ( .A(n_20), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_24), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_64), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_18), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_77), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_9), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_44), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_46), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_79), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_13), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_50), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_34), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_8), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_16), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_76), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_32), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_26), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_65), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_40), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g124 ( .A(n_5), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_35), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_4), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_66), .B(n_41), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_53), .Y(n_128) );
INVxp67_ASAP7_75t_SL g129 ( .A(n_18), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_125), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_125), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_125), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_124), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_87), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_88), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_87), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_104), .B(n_0), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_125), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_125), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_104), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_82), .B(n_0), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_122), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_91), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_91), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_122), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_92), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_83), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
BUFx2_ASAP7_75t_L g152 ( .A(n_103), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_93), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_84), .B(n_1), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_84), .B(n_1), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_95), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_85), .B(n_2), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_95), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_86), .B(n_2), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_108), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_93), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_111), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_98), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_86), .B(n_3), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_111), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_99), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_98), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_118), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_105), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_105), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_94), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_100), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_152), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_166), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_152), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_130), .Y(n_177) );
NAND3xp33_ASAP7_75t_L g178 ( .A(n_141), .B(n_80), .C(n_117), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_155), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_166), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_150), .B(n_118), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_166), .Y(n_182) );
NAND3xp33_ASAP7_75t_L g183 ( .A(n_141), .B(n_81), .C(n_109), .Y(n_183) );
NOR3xp33_ASAP7_75t_L g184 ( .A(n_137), .B(n_129), .C(n_89), .Y(n_184) );
AOI22x1_ASAP7_75t_L g185 ( .A1(n_162), .A2(n_128), .B1(n_113), .B2(n_112), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_155), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_166), .Y(n_187) );
AND2x6_ASAP7_75t_L g188 ( .A(n_155), .B(n_128), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_130), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_163), .B(n_119), .Y(n_190) );
AND2x6_ASAP7_75t_L g191 ( .A(n_156), .B(n_110), .Y(n_191) );
OR2x2_ASAP7_75t_SL g192 ( .A(n_137), .B(n_126), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_141), .B(n_120), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_156), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_166), .Y(n_195) );
INVx1_ASAP7_75t_SL g196 ( .A(n_140), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_161), .B(n_115), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_135), .B(n_116), .Y(n_199) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_135), .A2(n_106), .B(n_123), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_160), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_166), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_150), .B(n_94), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_153), .B(n_126), .Y(n_204) );
BUFx2_ASAP7_75t_L g205 ( .A(n_157), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_153), .B(n_97), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_130), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_160), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_168), .Y(n_209) );
AO22x2_ASAP7_75t_L g210 ( .A1(n_160), .A2(n_97), .B1(n_107), .B2(n_114), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_130), .Y(n_211) );
AND2x2_ASAP7_75t_SL g212 ( .A(n_165), .B(n_102), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_165), .B(n_96), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_159), .Y(n_215) );
AND2x6_ASAP7_75t_L g216 ( .A(n_142), .B(n_101), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_168), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_162), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_162), .Y(n_219) );
BUFx8_ASAP7_75t_L g220 ( .A(n_142), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_143), .B(n_121), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_143), .B(n_4), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_144), .B(n_5), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_168), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_170), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_168), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_168), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_144), .B(n_127), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_130), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_146), .B(n_151), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_168), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_146), .B(n_6), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_147), .B(n_7), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_147), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_149), .B(n_10), .Y(n_235) );
INVx4_ASAP7_75t_L g236 ( .A(n_173), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_170), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_130), .Y(n_238) );
AO22x2_ASAP7_75t_L g239 ( .A1(n_149), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_170), .Y(n_240) );
OR2x6_ASAP7_75t_L g241 ( .A(n_210), .B(n_171), .Y(n_241) );
INVx1_ASAP7_75t_SL g242 ( .A(n_196), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_220), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_230), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_230), .B(n_167), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_209), .Y(n_246) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_220), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_230), .Y(n_248) );
AND3x1_ASAP7_75t_L g249 ( .A(n_184), .B(n_158), .C(n_133), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_203), .B(n_206), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_222), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_203), .B(n_171), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_218), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_203), .B(n_145), .Y(n_254) );
AND3x1_ASAP7_75t_SL g255 ( .A(n_179), .B(n_172), .C(n_164), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_209), .Y(n_256) );
NOR3xp33_ASAP7_75t_SL g257 ( .A(n_178), .B(n_134), .C(n_136), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_219), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_206), .B(n_148), .Y(n_259) );
NOR3xp33_ASAP7_75t_SL g260 ( .A(n_183), .B(n_158), .C(n_154), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_224), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_224), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_234), .A2(n_151), .B(n_164), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_225), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_226), .Y(n_265) );
NOR2xp33_ASAP7_75t_R g266 ( .A(n_220), .B(n_154), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_222), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_226), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_206), .B(n_169), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_212), .A2(n_169), .B1(n_139), .B2(n_132), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_227), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_237), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_240), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_222), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_227), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_234), .B(n_169), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_213), .B(n_169), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_176), .Y(n_278) );
INVx3_ASAP7_75t_L g279 ( .A(n_223), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_193), .B(n_48), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_223), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_174), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_231), .Y(n_283) );
OR2x6_ASAP7_75t_L g284 ( .A(n_210), .B(n_139), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_213), .B(n_139), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_188), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_223), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_186), .B(n_11), .Y(n_288) );
AND3x1_ASAP7_75t_SL g289 ( .A(n_194), .B(n_13), .C(n_14), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_188), .B(n_132), .Y(n_290) );
NAND3xp33_ASAP7_75t_L g291 ( .A(n_198), .B(n_138), .C(n_132), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_231), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_188), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_188), .B(n_131), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_175), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_175), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_188), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_197), .B(n_15), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_212), .A2(n_131), .B1(n_138), .B2(n_17), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_201), .B(n_15), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_233), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_208), .B(n_52), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_214), .B(n_49), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_176), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_174), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_182), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_188), .B(n_204), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_210), .B(n_131), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_182), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_205), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_187), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_204), .B(n_138), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_251), .Y(n_313) );
INVx4_ASAP7_75t_L g314 ( .A(n_241), .Y(n_314) );
INVx5_ASAP7_75t_L g315 ( .A(n_241), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_241), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_253), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_254), .B(n_215), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_293), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_244), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_244), .Y(n_321) );
O2A1O1Ixp5_ASAP7_75t_L g322 ( .A1(n_302), .A2(n_199), .B(n_190), .C(n_221), .Y(n_322) );
OAI21x1_ASAP7_75t_SL g323 ( .A1(n_307), .A2(n_232), .B(n_185), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_251), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_242), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_253), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_241), .Y(n_327) );
AOI222xp33_ASAP7_75t_L g328 ( .A1(n_282), .A2(n_181), .B1(n_205), .B2(n_215), .C1(n_210), .C2(n_236), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_258), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_258), .Y(n_330) );
BUFx2_ASAP7_75t_SL g331 ( .A(n_293), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_252), .B(n_191), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_251), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_252), .B(n_236), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_263), .A2(n_199), .B(n_200), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_252), .B(n_236), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_264), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_251), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_248), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_310), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_250), .B(n_181), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_248), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_284), .B(n_235), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_284), .A2(n_191), .B1(n_235), .B2(n_233), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_269), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_249), .A2(n_191), .B1(n_235), .B2(n_233), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_287), .A2(n_192), .B1(n_239), .B2(n_228), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_251), .Y(n_348) );
INVx5_ASAP7_75t_L g349 ( .A(n_284), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_284), .B(n_191), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_287), .A2(n_192), .B1(n_239), .B2(n_228), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_264), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_297), .Y(n_353) );
BUFx3_ASAP7_75t_L g354 ( .A(n_297), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_308), .A2(n_191), .B1(n_216), .B2(n_200), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_301), .A2(n_200), .B(n_187), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_310), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_301), .A2(n_202), .B(n_195), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_286), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_286), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_308), .A2(n_191), .B1(n_216), .B2(n_239), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_267), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_308), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_269), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_288), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_272), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_278), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_356), .A2(n_274), .B(n_279), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_317), .Y(n_369) );
AOI22xp33_ASAP7_75t_SL g370 ( .A1(n_325), .A2(n_266), .B1(n_243), .B2(n_247), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_343), .B(n_308), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_315), .B(n_304), .Y(n_372) );
AOI21xp33_ASAP7_75t_L g373 ( .A1(n_347), .A2(n_303), .B(n_280), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_337), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_337), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_367), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_328), .A2(n_288), .B1(n_300), .B2(n_298), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_317), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_326), .B(n_267), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_344), .A2(n_361), .B1(n_349), .B2(n_355), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_315), .B(n_304), .Y(n_381) );
INVx6_ASAP7_75t_L g382 ( .A(n_315), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_366), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_340), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_326), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_315), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_336), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_329), .Y(n_388) );
NAND2xp33_ASAP7_75t_R g389 ( .A(n_316), .B(n_243), .Y(n_389) );
OAI22xp33_ASAP7_75t_L g390 ( .A1(n_315), .A2(n_305), .B1(n_245), .B2(n_279), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_357), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_336), .Y(n_392) );
INVx5_ASAP7_75t_L g393 ( .A(n_314), .Y(n_393) );
NAND3xp33_ASAP7_75t_L g394 ( .A(n_351), .B(n_260), .C(n_299), .Y(n_394) );
OAI211xp5_ASAP7_75t_L g395 ( .A1(n_346), .A2(n_257), .B(n_259), .C(n_277), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_349), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_349), .A2(n_298), .B1(n_288), .B2(n_300), .Y(n_397) );
BUFx4f_ASAP7_75t_SL g398 ( .A(n_336), .Y(n_398) );
INVx3_ASAP7_75t_L g399 ( .A(n_314), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_343), .B(n_267), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_329), .B(n_279), .Y(n_401) );
OA21x2_ASAP7_75t_L g402 ( .A1(n_368), .A2(n_323), .B(n_322), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_397), .A2(n_318), .B1(n_334), .B2(n_255), .Y(n_403) );
INVx2_ASAP7_75t_SL g404 ( .A(n_393), .Y(n_404) );
OAI211xp5_ASAP7_75t_SL g405 ( .A1(n_370), .A2(n_364), .B(n_345), .C(n_285), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_377), .A2(n_298), .B1(n_300), .B2(n_334), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_376), .B(n_341), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_369), .B(n_341), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_397), .A2(n_349), .B1(n_314), .B2(n_327), .Y(n_409) );
AOI21x1_ASAP7_75t_L g410 ( .A1(n_368), .A2(n_323), .B(n_335), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_369), .B(n_365), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_380), .A2(n_350), .B1(n_316), .B2(n_327), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_378), .Y(n_413) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_395), .A2(n_332), .B1(n_270), .B2(n_281), .C(n_320), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_378), .B(n_321), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_385), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_384), .Y(n_417) );
A2O1A1Ixp33_ASAP7_75t_L g418 ( .A1(n_394), .A2(n_366), .B(n_352), .C(n_330), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_393), .B(n_349), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_385), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_380), .A2(n_350), .B1(n_352), .B2(n_330), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_394), .A2(n_281), .B1(n_363), .B2(n_216), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_389), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_388), .Y(n_424) );
OAI22xp33_ASAP7_75t_L g425 ( .A1(n_398), .A2(n_363), .B1(n_281), .B2(n_339), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_400), .A2(n_216), .B1(n_342), .B2(n_239), .Y(n_426) );
A2O1A1Ixp33_ASAP7_75t_L g427 ( .A1(n_373), .A2(n_272), .B(n_273), .C(n_358), .Y(n_427) );
OAI21x1_ASAP7_75t_L g428 ( .A1(n_374), .A2(n_324), .B(n_294), .Y(n_428) );
OAI22xp33_ASAP7_75t_L g429 ( .A1(n_391), .A2(n_360), .B1(n_359), .B2(n_273), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_392), .A2(n_289), .B1(n_216), .B2(n_362), .Y(n_430) );
NOR5xp2_ASAP7_75t_SL g431 ( .A(n_409), .B(n_373), .C(n_19), .D(n_20), .E(n_16), .Y(n_431) );
INVx2_ASAP7_75t_SL g432 ( .A(n_419), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_413), .B(n_374), .Y(n_433) );
BUFx10_ASAP7_75t_L g434 ( .A(n_419), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_416), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_407), .B(n_388), .Y(n_436) );
OAI33xp33_ASAP7_75t_L g437 ( .A1(n_405), .A2(n_390), .A3(n_312), .B1(n_291), .B2(n_379), .B3(n_401), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_406), .A2(n_374), .B1(n_375), .B2(n_383), .Y(n_438) );
NOR2xp33_ASAP7_75t_R g439 ( .A(n_423), .B(n_393), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_420), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_424), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_421), .B(n_375), .Y(n_442) );
OR2x6_ASAP7_75t_L g443 ( .A(n_404), .B(n_386), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_419), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_404), .B(n_375), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_429), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_415), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_408), .B(n_383), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
OAI211xp5_ASAP7_75t_L g450 ( .A1(n_403), .A2(n_387), .B(n_400), .C(n_371), .Y(n_450) );
NAND5xp2_ASAP7_75t_SL g451 ( .A(n_423), .B(n_371), .C(n_393), .D(n_382), .E(n_386), .Y(n_451) );
OAI33xp33_ASAP7_75t_L g452 ( .A1(n_417), .A2(n_401), .A3(n_379), .B1(n_276), .B2(n_290), .B3(n_195), .Y(n_452) );
OAI221xp5_ASAP7_75t_L g453 ( .A1(n_430), .A2(n_399), .B1(n_383), .B2(n_396), .C(n_338), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_426), .A2(n_399), .B1(n_372), .B2(n_381), .C(n_396), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_412), .B(n_399), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_428), .Y(n_456) );
OAI221xp5_ASAP7_75t_L g457 ( .A1(n_422), .A2(n_399), .B1(n_396), .B2(n_338), .C(n_386), .Y(n_457) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_410), .A2(n_202), .B(n_295), .Y(n_458) );
OAI211xp5_ASAP7_75t_L g459 ( .A1(n_418), .A2(n_393), .B(n_180), .C(n_324), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
BUFx2_ASAP7_75t_L g461 ( .A(n_428), .Y(n_461) );
BUFx2_ASAP7_75t_L g462 ( .A(n_402), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_427), .Y(n_463) );
OAI33xp33_ASAP7_75t_L g464 ( .A1(n_425), .A2(n_295), .A3(n_296), .B1(n_311), .B2(n_309), .B3(n_306), .Y(n_464) );
OAI211xp5_ASAP7_75t_L g465 ( .A1(n_414), .A2(n_393), .B(n_180), .C(n_324), .Y(n_465) );
INVx4_ASAP7_75t_L g466 ( .A(n_402), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_402), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_455), .A2(n_381), .B1(n_372), .B2(n_382), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_467), .B(n_427), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_456), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_467), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_435), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_460), .B(n_138), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_434), .Y(n_474) );
INVxp67_ASAP7_75t_SL g475 ( .A(n_456), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_445), .B(n_393), .Y(n_476) );
BUFx2_ASAP7_75t_L g477 ( .A(n_443), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_435), .Y(n_478) );
OAI31xp33_ASAP7_75t_L g479 ( .A1(n_450), .A2(n_381), .A3(n_372), .B(n_354), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_441), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_441), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_440), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_433), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_434), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_462), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_442), .B(n_381), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_463), .B(n_138), .Y(n_487) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_458), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_445), .B(n_138), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_433), .Y(n_490) );
INVx4_ASAP7_75t_L g491 ( .A(n_443), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_462), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_461), .Y(n_493) );
AOI33xp33_ASAP7_75t_L g494 ( .A1(n_447), .A2(n_372), .A3(n_311), .B1(n_309), .B2(n_306), .B3(n_296), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_442), .B(n_382), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_461), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_448), .B(n_382), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_466), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_466), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_466), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_449), .B(n_382), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_448), .B(n_313), .Y(n_502) );
AND2x4_ASAP7_75t_SL g503 ( .A(n_434), .B(n_313), .Y(n_503) );
OAI221xp5_ASAP7_75t_L g504 ( .A1(n_436), .A2(n_362), .B1(n_331), .B2(n_180), .C(n_359), .Y(n_504) );
AOI221xp5_ASAP7_75t_SL g505 ( .A1(n_455), .A2(n_362), .B1(n_348), .B2(n_333), .C(n_313), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_458), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_458), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_443), .Y(n_508) );
NOR2x1_ASAP7_75t_L g509 ( .A(n_443), .B(n_331), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_439), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_446), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_438), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_432), .B(n_360), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_446), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_432), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_444), .B(n_454), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_444), .B(n_216), .Y(n_517) );
OAI211xp5_ASAP7_75t_L g518 ( .A1(n_459), .A2(n_362), .B(n_360), .C(n_359), .Y(n_518) );
OAI31xp33_ASAP7_75t_L g519 ( .A1(n_465), .A2(n_354), .A3(n_353), .B(n_319), .Y(n_519) );
AOI221x1_ASAP7_75t_L g520 ( .A1(n_431), .A2(n_348), .B1(n_333), .B2(n_313), .C(n_362), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_469), .B(n_21), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_498), .B(n_451), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_469), .B(n_23), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_469), .B(n_25), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_498), .B(n_451), .Y(n_525) );
AND2x2_ASAP7_75t_SL g526 ( .A(n_491), .B(n_431), .Y(n_526) );
INVxp67_ASAP7_75t_L g527 ( .A(n_484), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_483), .B(n_490), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_482), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_482), .B(n_457), .Y(n_530) );
NOR2x1p5_ASAP7_75t_L g531 ( .A(n_510), .B(n_464), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_471), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_500), .B(n_28), .Y(n_533) );
INVxp67_ASAP7_75t_L g534 ( .A(n_484), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_471), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_483), .B(n_453), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_470), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_520), .A2(n_437), .B(n_452), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_472), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_471), .B(n_29), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_472), .B(n_30), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_478), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_491), .Y(n_543) );
AOI32xp33_ASAP7_75t_L g544 ( .A1(n_474), .A2(n_319), .A3(n_353), .B1(n_217), .B2(n_45), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_478), .Y(n_545) );
OAI332xp33_ASAP7_75t_L g546 ( .A1(n_501), .A2(n_271), .A3(n_268), .B1(n_265), .B2(n_262), .B3(n_261), .C1(n_256), .C2(n_246), .Y(n_546) );
AOI31xp33_ASAP7_75t_L g547 ( .A1(n_484), .A2(n_36), .A3(n_37), .B(n_42), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_480), .B(n_47), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_479), .B(n_348), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_480), .Y(n_550) );
INVxp67_ASAP7_75t_L g551 ( .A(n_474), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_481), .B(n_56), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_481), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_485), .B(n_57), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_490), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_485), .B(n_59), .Y(n_556) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_491), .A2(n_360), .B1(n_359), .B2(n_348), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_485), .B(n_60), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_501), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_500), .B(n_61), .Y(n_560) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_470), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_497), .B(n_348), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_497), .B(n_333), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_486), .B(n_313), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_507), .Y(n_565) );
NOR3xp33_ASAP7_75t_SL g566 ( .A(n_479), .B(n_62), .C(n_63), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_486), .B(n_333), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_518), .A2(n_333), .B(n_359), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_516), .B(n_360), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_507), .Y(n_570) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_520), .B(n_238), .C(n_207), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_495), .B(n_68), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_515), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_515), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_492), .B(n_70), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_492), .B(n_71), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_495), .B(n_72), .Y(n_577) );
BUFx2_ASAP7_75t_L g578 ( .A(n_491), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_515), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_477), .B(n_73), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_516), .B(n_217), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_477), .B(n_217), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_555), .B(n_511), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_528), .B(n_508), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_551), .B(n_508), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_559), .A2(n_511), .B1(n_512), .B2(n_514), .C(n_496), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_529), .B(n_512), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_526), .A2(n_514), .B1(n_476), .B2(n_468), .Y(n_588) );
NAND4xp25_ASAP7_75t_L g589 ( .A(n_544), .B(n_505), .C(n_514), .D(n_494), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_547), .A2(n_509), .B(n_504), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_539), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_530), .A2(n_496), .B1(n_493), .B2(n_475), .C(n_473), .Y(n_592) );
OAI321xp33_ASAP7_75t_L g593 ( .A1(n_578), .A2(n_504), .A3(n_476), .B1(n_518), .B2(n_499), .C(n_475), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_526), .A2(n_509), .B1(n_502), .B2(n_473), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_537), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_527), .B(n_502), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_534), .B(n_493), .Y(n_597) );
OR4x1_ASAP7_75t_L g598 ( .A(n_543), .B(n_506), .C(n_505), .D(n_503), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_561), .B(n_492), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_549), .A2(n_503), .B1(n_499), .B2(n_506), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_545), .B(n_499), .Y(n_601) );
NAND2xp33_ASAP7_75t_SL g602 ( .A(n_566), .B(n_488), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_542), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_550), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_553), .Y(n_605) );
INVxp67_ASAP7_75t_L g606 ( .A(n_531), .Y(n_606) );
NAND2xp33_ASAP7_75t_SL g607 ( .A(n_543), .B(n_488), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_545), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_573), .Y(n_609) );
AO22x2_ASAP7_75t_L g610 ( .A1(n_532), .A2(n_507), .B1(n_473), .B2(n_487), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_522), .Y(n_611) );
INVx2_ASAP7_75t_SL g612 ( .A(n_522), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_532), .B(n_487), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_522), .B(n_503), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_535), .B(n_487), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_537), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_525), .B(n_489), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_525), .B(n_489), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_525), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_574), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_535), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_579), .Y(n_622) );
OAI22xp33_ASAP7_75t_L g623 ( .A1(n_549), .A2(n_488), .B1(n_513), .B2(n_517), .Y(n_623) );
AOI32xp33_ASAP7_75t_L g624 ( .A1(n_533), .A2(n_560), .A3(n_524), .B1(n_523), .B2(n_521), .Y(n_624) );
NOR2xp33_ASAP7_75t_R g625 ( .A(n_580), .B(n_517), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_536), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_533), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_546), .B(n_488), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_538), .B(n_519), .C(n_488), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_521), .B(n_488), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_523), .B(n_488), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_571), .A2(n_519), .B(n_261), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_533), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_560), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_SL g635 ( .A1(n_572), .A2(n_256), .B(n_283), .C(n_275), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_560), .B(n_189), .Y(n_636) );
AOI211xp5_ASAP7_75t_L g637 ( .A1(n_524), .A2(n_177), .B(n_207), .C(n_238), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_584), .B(n_565), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g639 ( .A(n_606), .Y(n_639) );
A2O1A1Ixp33_ASAP7_75t_L g640 ( .A1(n_624), .A2(n_557), .B(n_548), .C(n_552), .Y(n_640) );
INVx3_ASAP7_75t_L g641 ( .A(n_612), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_611), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_616), .B(n_565), .Y(n_643) );
CKINVDCx16_ASAP7_75t_R g644 ( .A(n_590), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_626), .B(n_570), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_585), .B(n_570), .Y(n_646) );
INVxp67_ASAP7_75t_SL g647 ( .A(n_595), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_591), .Y(n_648) );
AOI22x1_ASAP7_75t_L g649 ( .A1(n_590), .A2(n_548), .B1(n_541), .B2(n_552), .Y(n_649) );
XNOR2xp5_ASAP7_75t_L g650 ( .A(n_596), .B(n_569), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_603), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_597), .B(n_558), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_583), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_583), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_593), .B(n_600), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_593), .B(n_558), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_617), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_604), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_616), .B(n_564), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_619), .B(n_581), .Y(n_660) );
AND2x4_ASAP7_75t_SL g661 ( .A(n_618), .B(n_540), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_605), .B(n_567), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_587), .B(n_554), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_609), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g665 ( .A1(n_628), .A2(n_541), .B(n_540), .C(n_568), .Y(n_665) );
BUFx2_ASAP7_75t_L g666 ( .A(n_599), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_615), .B(n_563), .Y(n_667) );
XOR2xp5_ASAP7_75t_L g668 ( .A(n_588), .B(n_577), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_586), .B(n_576), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_631), .B(n_554), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_620), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_600), .B(n_576), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_592), .B(n_575), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_621), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_607), .B(n_637), .Y(n_675) );
NAND3xp33_ASAP7_75t_SL g676 ( .A(n_640), .B(n_602), .C(n_614), .Y(n_676) );
NAND4xp75_ASAP7_75t_L g677 ( .A(n_655), .B(n_594), .C(n_636), .D(n_633), .Y(n_677) );
AOI32xp33_ASAP7_75t_L g678 ( .A1(n_655), .A2(n_666), .A3(n_672), .B1(n_656), .B2(n_644), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_653), .B(n_622), .Y(n_679) );
OAI22xp5_ASAP7_75t_SL g680 ( .A1(n_642), .A2(n_598), .B1(n_634), .B2(n_627), .Y(n_680) );
INVx2_ASAP7_75t_SL g681 ( .A(n_638), .Y(n_681) );
INVx3_ASAP7_75t_L g682 ( .A(n_641), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_640), .B(n_623), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_645), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_664), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_672), .A2(n_589), .B1(n_610), .B2(n_629), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_641), .B(n_608), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_671), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_654), .B(n_610), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_643), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_648), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_639), .B(n_613), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_656), .A2(n_610), .B1(n_630), .B2(n_613), .Y(n_693) );
OAI211xp5_ASAP7_75t_L g694 ( .A1(n_649), .A2(n_625), .B(n_635), .C(n_632), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_651), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_658), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_668), .A2(n_562), .B1(n_601), .B2(n_575), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_647), .Y(n_698) );
O2A1O1Ixp33_ASAP7_75t_L g699 ( .A1(n_665), .A2(n_582), .B(n_556), .C(n_265), .Y(n_699) );
AOI221xp5_ASAP7_75t_SL g700 ( .A1(n_683), .A2(n_657), .B1(n_665), .B2(n_642), .C(n_650), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_686), .B(n_669), .Y(n_701) );
OAI22xp33_ASAP7_75t_SL g702 ( .A1(n_686), .A2(n_675), .B1(n_673), .B2(n_662), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_676), .B(n_675), .C(n_660), .Y(n_703) );
NOR2xp67_ASAP7_75t_L g704 ( .A(n_693), .B(n_682), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_678), .B(n_660), .C(n_659), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_684), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_698), .B(n_674), .C(n_663), .Y(n_707) );
NAND5xp2_ASAP7_75t_L g708 ( .A(n_699), .B(n_556), .C(n_652), .D(n_670), .E(n_646), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_685), .Y(n_709) );
INVxp67_ASAP7_75t_L g710 ( .A(n_689), .Y(n_710) );
AOI211xp5_ASAP7_75t_L g711 ( .A1(n_680), .A2(n_667), .B(n_674), .C(n_661), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_679), .A2(n_661), .B1(n_177), .B2(n_207), .C(n_238), .Y(n_712) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_694), .A2(n_177), .B1(n_207), .B2(n_238), .C(n_211), .Y(n_713) );
NAND4xp75_ASAP7_75t_L g714 ( .A(n_692), .B(n_246), .C(n_283), .D(n_275), .Y(n_714) );
OA22x2_ASAP7_75t_L g715 ( .A1(n_682), .A2(n_292), .B1(n_271), .B2(n_268), .Y(n_715) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_697), .A2(n_177), .B1(n_238), .B2(n_207), .C(n_211), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_688), .A2(n_177), .B1(n_189), .B2(n_211), .C(n_229), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_677), .A2(n_189), .B1(n_211), .B2(n_229), .Y(n_718) );
AOI221x1_ASAP7_75t_L g719 ( .A1(n_691), .A2(n_189), .B1(n_229), .B2(n_262), .C(n_292), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_687), .B(n_229), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_687), .B(n_681), .Y(n_721) );
NAND4xp25_ASAP7_75t_L g722 ( .A(n_700), .B(n_703), .C(n_711), .D(n_701), .Y(n_722) );
NOR3xp33_ASAP7_75t_SL g723 ( .A(n_713), .B(n_718), .C(n_705), .Y(n_723) );
OAI222xp33_ASAP7_75t_L g724 ( .A1(n_710), .A2(n_721), .B1(n_702), .B2(n_715), .C1(n_706), .C2(n_709), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_710), .B(n_704), .Y(n_725) );
CKINVDCx5p33_ASAP7_75t_R g726 ( .A(n_695), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_726), .Y(n_727) );
XNOR2xp5_ASAP7_75t_L g728 ( .A(n_722), .B(n_714), .Y(n_728) );
OR2x2_ASAP7_75t_L g729 ( .A(n_725), .B(n_707), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_727), .Y(n_730) );
OR2x2_ASAP7_75t_L g731 ( .A(n_729), .B(n_690), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_730), .A2(n_728), .B1(n_723), .B2(n_724), .Y(n_732) );
INVx3_ASAP7_75t_L g733 ( .A(n_731), .Y(n_733) );
AOI222xp33_ASAP7_75t_L g734 ( .A1(n_733), .A2(n_712), .B1(n_696), .B2(n_720), .C1(n_716), .C2(n_717), .Y(n_734) );
O2A1O1Ixp5_ASAP7_75t_SL g735 ( .A1(n_734), .A2(n_732), .B(n_719), .C(n_708), .Y(n_735) );
endmodule