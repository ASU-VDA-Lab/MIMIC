module fake_jpeg_30818_n_64 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_17),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_14),
.B(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_15),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_28),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_17),
.C(n_20),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_18),
.C(n_11),
.Y(n_38)
);

OR2x2_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_8),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_8),
.B1(n_12),
.B2(n_10),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_34),
.B1(n_9),
.B2(n_19),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_21),
.B1(n_18),
.B2(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_39),
.Y(n_44)
);

OA21x2_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_11),
.B(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_18),
.C(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_45),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_10),
.C(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_37),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_45),
.B(n_2),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_41),
.C(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_55),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_49),
.A2(n_42),
.B1(n_40),
.B2(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_1),
.B(n_3),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_51),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_49),
.C(n_2),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_60),
.B(n_58),
.Y(n_61)
);

AOI322xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_57),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_7),
.C2(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_4),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_7),
.Y(n_64)
);


endmodule