module fake_jpeg_30467_n_226 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_50),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_56),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_58),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_60),
.Y(n_87)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g97 ( 
.A(n_61),
.B(n_66),
.CON(n_97),
.SN(n_97)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_63),
.Y(n_70)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_36),
.B1(n_20),
.B2(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_28),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_26),
.B(n_36),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_41),
.B(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_92),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_34),
.B1(n_24),
.B2(n_37),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_77),
.B1(n_83),
.B2(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_80),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_34),
.B1(n_21),
.B2(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_28),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_33),
.B1(n_40),
.B2(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_30),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_89),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_38),
.B(n_35),
.C(n_22),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_61),
.B(n_64),
.C(n_59),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_22),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_90),
.A2(n_42),
.B1(n_6),
.B2(n_7),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_37),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_48),
.B(n_32),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_0),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_100),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_4),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_88),
.Y(n_103)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_5),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_118),
.Y(n_129)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_114),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_70),
.C(n_76),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_82),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_5),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_125),
.B1(n_128),
.B2(n_9),
.Y(n_138)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_124),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_6),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_81),
.A2(n_96),
.B1(n_98),
.B2(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_8),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_90),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_128)
);

NOR2x1_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_130),
.B(n_117),
.Y(n_165)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_123),
.Y(n_133)
);

NAND2x1_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_113),
.Y(n_162)
);

AOI32xp33_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_86),
.A3(n_87),
.B1(n_77),
.B2(n_73),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_113),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_148),
.B1(n_114),
.B2(n_101),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_91),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_152),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_67),
.B(n_94),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_110),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_96),
.B1(n_74),
.B2(n_93),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_116),
.C(n_112),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_9),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_157),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_107),
.B(n_116),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_158),
.B(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_102),
.B(n_109),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_142),
.B1(n_138),
.B2(n_148),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_165),
.B(n_147),
.C(n_13),
.D(n_15),
.Y(n_187)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_115),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_167),
.C(n_169),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_164),
.B(n_171),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_119),
.B(n_127),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_SL g188 ( 
.A(n_166),
.B(n_147),
.C(n_93),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_103),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_172),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_106),
.C(n_108),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_10),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_146),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_185),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_142),
.A3(n_136),
.B1(n_132),
.B2(n_140),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_182),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_158),
.A2(n_129),
.B(n_132),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_180),
.A2(n_161),
.B(n_131),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_149),
.B1(n_143),
.B2(n_151),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_152),
.A3(n_149),
.B1(n_151),
.B2(n_146),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_146),
.B1(n_118),
.B2(n_122),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_15),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_172),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_167),
.C(n_163),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_193),
.B(n_196),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_170),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_197),
.A2(n_180),
.B(n_174),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_183),
.B(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_200),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_181),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_206),
.Y(n_211)
);

AOI321xp33_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_182),
.A3(n_187),
.B1(n_179),
.B2(n_183),
.C(n_188),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g209 ( 
.A(n_204),
.Y(n_209)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_176),
.C(n_186),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_202),
.C(n_204),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_213),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_210),
.B(n_203),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_208),
.A2(n_191),
.B1(n_186),
.B2(n_199),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_215),
.A2(n_197),
.B1(n_200),
.B2(n_211),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_219),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_209),
.B1(n_12),
.B2(n_13),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_207),
.B(n_208),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_222),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_216),
.B(n_218),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_223),
.B(n_221),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_224),
.Y(n_226)
);


endmodule