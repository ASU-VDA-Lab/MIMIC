module fake_netlist_6_2184_n_1780 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1780);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1780;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx10_ASAP7_75t_L g169 ( 
.A(n_48),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_87),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_93),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_112),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_58),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_166),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_79),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_57),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_139),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_35),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_167),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_45),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_78),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_148),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_102),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_24),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_98),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_46),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_49),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_103),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_156),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_30),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

BUFx2_ASAP7_75t_R g204 ( 
.A(n_97),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_15),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_35),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_92),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_105),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_37),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_73),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_28),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_96),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_154),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_71),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_21),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_56),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_9),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_141),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_2),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_14),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_82),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_130),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_57),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_20),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_26),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_90),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_91),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_116),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_101),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_75),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_12),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_66),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_3),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_70),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_24),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_0),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_53),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_60),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_1),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_89),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_132),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_3),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_6),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_88),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_31),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_77),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_8),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_53),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_21),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_32),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_134),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_25),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_58),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_4),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_14),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_164),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_86),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_2),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_55),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_159),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_63),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_80),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_140),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_52),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_67),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_4),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_104),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_51),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_165),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_32),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_22),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_115),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_107),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_69),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_84),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_52),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_28),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_113),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_29),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_163),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_27),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_16),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_7),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_157),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_145),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_10),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_18),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_11),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_20),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_44),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_99),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_160),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_95),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_40),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_22),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_48),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_72),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_121),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_138),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_56),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_54),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_51),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_129),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_64),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_33),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_74),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_168),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_8),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_9),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_42),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_142),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_152),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_46),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_16),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_55),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_85),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_36),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_131),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_10),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_83),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_59),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_13),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_161),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_27),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_47),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_151),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_143),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_123),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_5),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_18),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_36),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_147),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_81),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_114),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_49),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_171),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_199),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_209),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_174),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_174),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_178),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_183),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_199),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_201),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_212),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_179),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_238),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_199),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_199),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_199),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_237),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_214),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_273),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_196),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_199),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_170),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_199),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_211),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_227),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_211),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_211),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_211),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_211),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_211),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_211),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_251),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_215),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g371 ( 
.A(n_189),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_251),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_251),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_223),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_225),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_251),
.Y(n_376)
);

INVxp33_ASAP7_75t_L g377 ( 
.A(n_297),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_251),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_230),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_227),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_227),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_279),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_279),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_294),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_246),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_232),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_179),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_246),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_181),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_187),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_196),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_216),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_219),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_210),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_236),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_305),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_233),
.Y(n_397)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_189),
.Y(n_398)
);

INVxp33_ASAP7_75t_L g399 ( 
.A(n_250),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_255),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_210),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_258),
.Y(n_402)
);

INVxp33_ASAP7_75t_SL g403 ( 
.A(n_193),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_261),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_193),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_271),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_200),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_243),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_198),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_285),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_298),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_299),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_200),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_169),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_334),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_303),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_312),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_317),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_320),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_322),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_325),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_226),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_169),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_176),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_247),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_425),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_339),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_425),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_344),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_353),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_369),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_369),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_372),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_372),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_345),
.B(n_268),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_R g437 ( 
.A(n_347),
.B(n_287),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_373),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_348),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_424),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_376),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_376),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_355),
.Y(n_445)
);

INVx5_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_378),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_378),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_340),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_391),
.B(n_226),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_370),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_374),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_340),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_342),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_203),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_346),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_346),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_351),
.Y(n_458)
);

AND2x6_ASAP7_75t_L g459 ( 
.A(n_351),
.B(n_176),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_362),
.B(n_203),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_352),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_343),
.A2(n_177),
.B1(n_328),
.B2(n_228),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_396),
.A2(n_228),
.B1(n_328),
.B2(n_177),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_375),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_379),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_352),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_380),
.B(n_173),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_386),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_414),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_358),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_415),
.B(n_204),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_397),
.B(n_173),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_349),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_358),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_357),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_405),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_360),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_380),
.B(n_264),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_387),
.Y(n_479)
);

AND2x2_ASAP7_75t_SL g480 ( 
.A(n_354),
.B(n_264),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_360),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_408),
.B(n_426),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_361),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_361),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_363),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_363),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_364),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_364),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_407),
.B(n_172),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_407),
.B(n_175),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_365),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_365),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_381),
.B(n_180),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_366),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_L g495 ( 
.A(n_409),
.B(n_198),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_405),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_366),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_367),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_367),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_341),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_368),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_368),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_394),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_384),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_475),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_453),
.Y(n_506)
);

INVxp33_ASAP7_75t_L g507 ( 
.A(n_469),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_431),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_453),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_480),
.B(n_371),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_456),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_472),
.B(n_398),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_438),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_475),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_438),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_443),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_482),
.B(n_403),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_L g519 ( 
.A(n_459),
.B(n_176),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_437),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_443),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_440),
.Y(n_522)
);

NAND3xp33_ASAP7_75t_L g523 ( 
.A(n_495),
.B(n_496),
.C(n_460),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_359),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_480),
.B(n_377),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_440),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_500),
.B(n_341),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_457),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_440),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_440),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_494),
.B(n_381),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_457),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_500),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_458),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_431),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_480),
.B(n_428),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_494),
.B(n_188),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_449),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_455),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_504),
.Y(n_540)
);

AND3x2_ASAP7_75t_L g541 ( 
.A(n_471),
.B(n_350),
.C(n_220),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_494),
.B(n_194),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_450),
.B(n_388),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_461),
.Y(n_544)
);

BUFx4f_ASAP7_75t_L g545 ( 
.A(n_449),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_461),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_455),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_458),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_430),
.B(n_287),
.Y(n_549)
);

BUFx4f_ASAP7_75t_L g550 ( 
.A(n_449),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_436),
.B(n_450),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_477),
.B(n_263),
.Y(n_552)
);

AND2x2_ASAP7_75t_SL g553 ( 
.A(n_493),
.B(n_176),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_477),
.B(n_249),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_481),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_466),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_466),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_441),
.B(n_306),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_431),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_431),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_460),
.A2(n_306),
.B1(n_315),
.B2(n_326),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_470),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_445),
.B(n_315),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_431),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_483),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_476),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_470),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_485),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_483),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_485),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_484),
.B(n_259),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_492),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_451),
.B(n_326),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_493),
.B(n_176),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_484),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_492),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_452),
.A2(n_350),
.B1(n_191),
.B2(n_314),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_431),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_464),
.B(n_203),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_486),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_454),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_465),
.B(n_356),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_487),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_487),
.B(n_260),
.Y(n_585)
);

AOI21x1_ASAP7_75t_L g586 ( 
.A1(n_488),
.A2(n_195),
.B(n_182),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_459),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_468),
.B(n_184),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_502),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_476),
.B(n_385),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_442),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_488),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_442),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_498),
.B(n_265),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_493),
.B(n_389),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_489),
.A2(n_192),
.B1(n_191),
.B2(n_190),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_498),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_499),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_499),
.Y(n_599)
);

BUFx10_ASAP7_75t_L g600 ( 
.A(n_493),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_501),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_467),
.A2(n_399),
.B1(n_276),
.B2(n_323),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_446),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_502),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_427),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_446),
.B(n_266),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_467),
.B(n_388),
.Y(n_607)
);

NAND3xp33_ASAP7_75t_L g608 ( 
.A(n_490),
.B(n_205),
.C(n_202),
.Y(n_608)
);

BUFx10_ASAP7_75t_L g609 ( 
.A(n_467),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_427),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_446),
.B(n_275),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_427),
.Y(n_612)
);

CKINVDCx6p67_ASAP7_75t_R g613 ( 
.A(n_473),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_474),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_427),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_446),
.B(n_277),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_474),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_474),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_479),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_432),
.Y(n_620)
);

AND3x1_ASAP7_75t_L g621 ( 
.A(n_463),
.B(n_423),
.C(n_390),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_463),
.A2(n_332),
.B1(n_338),
.B2(n_262),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_427),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_446),
.B(n_281),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_432),
.Y(n_625)
);

NAND3xp33_ASAP7_75t_L g626 ( 
.A(n_467),
.B(n_218),
.C(n_206),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_478),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_503),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_446),
.B(n_283),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_474),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_462),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_449),
.B(n_288),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_449),
.Y(n_633)
);

AND2x6_ASAP7_75t_L g634 ( 
.A(n_478),
.B(n_244),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_478),
.B(n_389),
.Y(n_635)
);

AND3x1_ASAP7_75t_L g636 ( 
.A(n_433),
.B(n_423),
.C(n_392),
.Y(n_636)
);

NAND3xp33_ASAP7_75t_L g637 ( 
.A(n_478),
.B(n_222),
.C(n_221),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_449),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_427),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_491),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_491),
.B(n_401),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_429),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_491),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_433),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_434),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_491),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_434),
.Y(n_647)
);

AO22x2_ASAP7_75t_L g648 ( 
.A1(n_435),
.A2(n_310),
.B1(n_197),
.B2(n_207),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_429),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_491),
.B(n_184),
.Y(n_650)
);

BUFx10_ASAP7_75t_L g651 ( 
.A(n_459),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_429),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_435),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_459),
.A2(n_323),
.B1(n_276),
.B2(n_244),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_551),
.B(n_539),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_522),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_539),
.B(n_491),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_627),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_547),
.B(n_497),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_547),
.B(n_497),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_553),
.B(n_497),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_511),
.B(n_497),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_533),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_553),
.B(n_497),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_607),
.Y(n_665)
);

AND2x4_ASAP7_75t_SL g666 ( 
.A(n_613),
.B(n_169),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_507),
.B(n_257),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_607),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_609),
.B(n_523),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_512),
.B(n_185),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_591),
.B(n_257),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_526),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_609),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_511),
.B(n_497),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_526),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_609),
.B(n_244),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_648),
.A2(n_244),
.B1(n_276),
.B2(n_323),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_529),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_SL g679 ( 
.A1(n_631),
.A2(n_311),
.B1(n_313),
.B2(n_290),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_528),
.Y(n_680)
);

NAND2x1p5_ASAP7_75t_L g681 ( 
.A(n_595),
.B(n_208),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_528),
.B(n_439),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_529),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_532),
.B(n_544),
.Y(n_684)
);

AOI22x1_ASAP7_75t_L g685 ( 
.A1(n_614),
.A2(n_224),
.B1(n_278),
.B2(n_272),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_530),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_600),
.B(n_244),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_632),
.A2(n_550),
.B(n_545),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_593),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_532),
.B(n_444),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_600),
.B(n_276),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_L g692 ( 
.A(n_520),
.B(n_518),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_530),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_544),
.B(n_444),
.Y(n_694)
);

BUFx5_ASAP7_75t_L g695 ( 
.A(n_614),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_591),
.B(n_257),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_600),
.B(n_595),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_546),
.B(n_447),
.Y(n_698)
);

INVx4_ASAP7_75t_SL g699 ( 
.A(n_574),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_546),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_534),
.Y(n_701)
);

OR2x6_ASAP7_75t_L g702 ( 
.A(n_619),
.B(n_392),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_555),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_555),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_510),
.A2(n_324),
.B1(n_295),
.B2(n_300),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_565),
.B(n_575),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_527),
.B(n_393),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_566),
.B(n_533),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_595),
.B(n_276),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_525),
.B(n_185),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_566),
.B(n_393),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_565),
.B(n_447),
.Y(n_712)
);

NAND2x1_ASAP7_75t_L g713 ( 
.A(n_610),
.B(n_459),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_506),
.A2(n_241),
.B(n_213),
.C(n_254),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_602),
.A2(n_235),
.B1(n_319),
.B2(n_231),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_575),
.B(n_448),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_543),
.A2(n_410),
.B(n_395),
.C(n_400),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_543),
.B(n_274),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_534),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_537),
.B(n_542),
.Y(n_720)
);

O2A1O1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_524),
.A2(n_552),
.B(n_531),
.C(n_577),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_581),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_561),
.B(n_395),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_590),
.B(n_400),
.Y(n_724)
);

INVx5_ASAP7_75t_L g725 ( 
.A(n_651),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_648),
.A2(n_584),
.B1(n_597),
.B2(n_581),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_584),
.B(n_323),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_631),
.A2(n_622),
.B1(n_590),
.B2(n_578),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_641),
.A2(n_331),
.B1(n_301),
.B2(n_302),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_548),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_597),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_598),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_590),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_548),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_509),
.B(n_186),
.Y(n_735)
);

INVx6_ASAP7_75t_L g736 ( 
.A(n_540),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_598),
.B(n_459),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_569),
.A2(n_296),
.B(n_229),
.C(n_270),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_556),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_536),
.A2(n_321),
.B1(n_307),
.B2(n_309),
.Y(n_740)
);

A2O1A1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_592),
.A2(n_217),
.B(n_416),
.C(n_422),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_556),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_557),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_599),
.B(n_587),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_601),
.B(n_186),
.Y(n_745)
);

BUFx8_ASAP7_75t_L g746 ( 
.A(n_619),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_599),
.B(n_323),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_635),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_557),
.Y(n_749)
);

NAND2x1_ASAP7_75t_L g750 ( 
.A(n_610),
.B(n_459),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_613),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_635),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_505),
.B(n_429),
.Y(n_753)
);

NOR2xp67_ASAP7_75t_L g754 ( 
.A(n_608),
.B(n_329),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_L g755 ( 
.A(n_514),
.B(n_330),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_514),
.B(n_429),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_562),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_650),
.B(n_429),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_636),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_567),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_554),
.B(n_190),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_628),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_571),
.B(n_314),
.Y(n_763)
);

BUFx5_ASAP7_75t_L g764 ( 
.A(n_617),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_587),
.B(n_335),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_628),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_585),
.B(n_335),
.Y(n_767)
);

BUFx8_ASAP7_75t_L g768 ( 
.A(n_540),
.Y(n_768)
);

BUFx4_ASAP7_75t_L g769 ( 
.A(n_540),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_594),
.B(n_336),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_648),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_648),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_517),
.B(n_402),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_583),
.B(n_517),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_617),
.B(n_337),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_630),
.B(n_337),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_549),
.B(n_274),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_582),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_588),
.B(n_234),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_SL g780 ( 
.A1(n_621),
.A2(n_311),
.B1(n_313),
.B2(n_239),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_620),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_596),
.B(n_240),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_580),
.B(n_242),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_626),
.B(n_637),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_625),
.B(n_402),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_630),
.B(n_404),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_618),
.B(n_404),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_625),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_568),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_568),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_644),
.B(n_406),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_644),
.B(n_406),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_654),
.A2(n_292),
.B1(n_291),
.B2(n_274),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_645),
.B(n_410),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_558),
.Y(n_795)
);

OAI22x1_ASAP7_75t_SL g796 ( 
.A1(n_541),
.A2(n_293),
.B1(n_248),
.B2(n_252),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_653),
.B(n_245),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_570),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_570),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_572),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_647),
.B(n_411),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_563),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_653),
.B(n_411),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_633),
.B(n_638),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_572),
.A2(n_422),
.B(n_421),
.C(n_420),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_633),
.B(n_253),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_638),
.B(n_412),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_573),
.A2(n_643),
.B1(n_640),
.B2(n_574),
.Y(n_808)
);

NOR2xp67_ASAP7_75t_L g809 ( 
.A(n_606),
.B(n_412),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_513),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_701),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_719),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_762),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_655),
.B(n_576),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_673),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_655),
.B(n_651),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_673),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_708),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_670),
.A2(n_640),
.B1(n_643),
.B2(n_574),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_670),
.B(n_538),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_782),
.A2(n_589),
.B1(n_576),
.B2(n_604),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_703),
.B(n_589),
.Y(n_822)
);

AO22x2_ASAP7_75t_L g823 ( 
.A1(n_723),
.A2(n_418),
.B1(n_420),
.B2(n_416),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_781),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_673),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_784),
.A2(n_574),
.B1(n_535),
.B2(n_508),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_766),
.Y(n_827)
);

NOR2xp67_ASAP7_75t_L g828 ( 
.A(n_689),
.B(n_611),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_SL g829 ( 
.A(n_795),
.B(n_733),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_658),
.B(n_417),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_673),
.B(n_651),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_663),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_SL g833 ( 
.A1(n_679),
.A2(n_267),
.B1(n_256),
.B2(n_269),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_703),
.B(n_604),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_751),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_730),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_720),
.B(n_508),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_734),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_R g839 ( 
.A(n_736),
.B(n_586),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_784),
.A2(n_574),
.B1(n_508),
.B2(n_535),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_720),
.B(n_535),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_677),
.A2(n_280),
.B1(n_282),
.B2(n_284),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_R g843 ( 
.A(n_736),
.B(n_586),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_684),
.B(n_706),
.Y(n_844)
);

AOI21x1_ASAP7_75t_L g845 ( 
.A1(n_661),
.A2(n_616),
.B(n_624),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_736),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_711),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_680),
.B(n_560),
.Y(n_848)
);

BUFx4f_ASAP7_75t_L g849 ( 
.A(n_702),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_739),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_689),
.B(n_538),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_692),
.B(n_587),
.Y(n_852)
);

BUFx12f_ASAP7_75t_SL g853 ( 
.A(n_702),
.Y(n_853)
);

AND2x4_ASAP7_75t_SL g854 ( 
.A(n_778),
.B(n_291),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_659),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_707),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_700),
.B(n_704),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_SL g858 ( 
.A1(n_802),
.A2(n_780),
.B1(n_782),
.B2(n_783),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_768),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_802),
.B(n_545),
.Y(n_860)
);

AND2x2_ASAP7_75t_SL g861 ( 
.A(n_793),
.B(n_519),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_722),
.B(n_560),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_731),
.B(n_564),
.Y(n_863)
);

BUFx8_ASAP7_75t_L g864 ( 
.A(n_671),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_732),
.B(n_564),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_721),
.B(n_564),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_788),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_785),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_785),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_718),
.B(n_291),
.Y(n_870)
);

INVx5_ASAP7_75t_L g871 ( 
.A(n_725),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_667),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_726),
.B(n_513),
.Y(n_873)
);

INVx5_ASAP7_75t_L g874 ( 
.A(n_725),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_726),
.B(n_515),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_710),
.A2(n_521),
.B(n_516),
.C(n_515),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_759),
.B(n_538),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_665),
.B(n_516),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_771),
.A2(n_519),
.B(n_521),
.C(n_629),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_748),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_742),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_752),
.Y(n_882)
);

NOR2x1p5_ASAP7_75t_L g883 ( 
.A(n_724),
.B(n_286),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_743),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_669),
.A2(n_668),
.B1(n_697),
.B2(n_710),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_759),
.B(n_646),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_749),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_778),
.B(n_646),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_810),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_L g890 ( 
.A(n_725),
.B(n_574),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_746),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_768),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_695),
.B(n_610),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_757),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_695),
.B(n_612),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_728),
.B(n_646),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_779),
.A2(n_545),
.B(n_550),
.C(n_642),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_774),
.B(n_550),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_760),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_661),
.A2(n_615),
.B(n_642),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_728),
.B(n_779),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_702),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_773),
.B(n_417),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_761),
.B(n_559),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_773),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_696),
.B(n_292),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_725),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_789),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_777),
.B(n_559),
.Y(n_909)
);

OR2x6_ASAP7_75t_L g910 ( 
.A(n_771),
.B(n_418),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_790),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_798),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_697),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_799),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_800),
.Y(n_915)
);

OR2x6_ASAP7_75t_L g916 ( 
.A(n_772),
.B(n_419),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_807),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_791),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_656),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_792),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_763),
.B(n_559),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_699),
.B(n_419),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_794),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_746),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_801),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_713),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_767),
.B(n_559),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_695),
.B(n_764),
.Y(n_928)
);

AND2x6_ASAP7_75t_L g929 ( 
.A(n_808),
.B(n_559),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_695),
.B(n_615),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_796),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_783),
.A2(n_615),
.B(n_623),
.C(n_421),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_695),
.B(n_623),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_770),
.B(n_579),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_735),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_681),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_672),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_750),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_803),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_664),
.A2(n_603),
.B(n_579),
.Y(n_940)
);

BUFx12f_ASAP7_75t_L g941 ( 
.A(n_681),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_695),
.B(n_579),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_675),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_SL g944 ( 
.A1(n_793),
.A2(n_289),
.B1(n_333),
.B2(n_304),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_764),
.B(n_579),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_678),
.Y(n_946)
);

NOR3xp33_ASAP7_75t_L g947 ( 
.A(n_735),
.B(n_308),
.C(n_316),
.Y(n_947)
);

NAND2x1p5_ASAP7_75t_L g948 ( 
.A(n_657),
.B(n_660),
.Y(n_948)
);

NAND2x1p5_ASAP7_75t_L g949 ( 
.A(n_657),
.B(n_652),
.Y(n_949)
);

INVx4_ASAP7_75t_L g950 ( 
.A(n_699),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_683),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_682),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_769),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_775),
.B(n_318),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_764),
.B(n_652),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_690),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_797),
.B(n_740),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_745),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_776),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_694),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_797),
.B(n_652),
.Y(n_961)
);

AND3x1_ASAP7_75t_SL g962 ( 
.A(n_666),
.B(n_383),
.C(n_382),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_699),
.B(n_382),
.Y(n_963)
);

INVx5_ASAP7_75t_L g964 ( 
.A(n_686),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_745),
.B(n_652),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_698),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_712),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_705),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_806),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_787),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_717),
.B(n_383),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_764),
.B(n_652),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_729),
.B(n_649),
.Y(n_973)
);

OR2x6_ASAP7_75t_L g974 ( 
.A(n_717),
.B(n_603),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_693),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_716),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_715),
.A2(n_634),
.B1(n_639),
.B2(n_649),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_809),
.A2(n_634),
.B1(n_639),
.B2(n_649),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_764),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_660),
.B(n_649),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_764),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_804),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_786),
.B(n_649),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_744),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_906),
.B(n_806),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_815),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_901),
.A2(n_664),
.B1(n_709),
.B2(n_676),
.Y(n_987)
);

INVx4_ASAP7_75t_L g988 ( 
.A(n_815),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_844),
.A2(n_676),
.B1(n_687),
.B2(n_691),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_979),
.A2(n_758),
.B(n_688),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_935),
.B(n_687),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_979),
.A2(n_753),
.B(n_756),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_878),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_905),
.B(n_754),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_SL g995 ( 
.A(n_858),
.B(n_292),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_958),
.A2(n_714),
.B(n_738),
.C(n_741),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_957),
.A2(n_755),
.B(n_747),
.C(n_727),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_844),
.B(n_662),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_969),
.B(n_674),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_815),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_813),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_943),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_943),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_975),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_968),
.A2(n_691),
.B1(n_765),
.B2(n_744),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_979),
.A2(n_737),
.B(n_765),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_979),
.A2(n_639),
.B(n_605),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_878),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_872),
.B(n_747),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_952),
.B(n_956),
.Y(n_1010)
);

BUFx2_ASAP7_75t_R g1011 ( 
.A(n_859),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_905),
.B(n_868),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_L g1013 ( 
.A(n_833),
.B(n_805),
.C(n_727),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_975),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_959),
.B(n_639),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_SL g1016 ( 
.A(n_817),
.B(n_685),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_818),
.B(n_639),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_857),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_928),
.A2(n_605),
.B(n_805),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_960),
.B(n_634),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_966),
.B(n_634),
.Y(n_1021)
);

BUFx12f_ASAP7_75t_L g1022 ( 
.A(n_924),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_835),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_825),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_832),
.B(n_605),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_827),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_857),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_880),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_896),
.A2(n_605),
.B1(n_146),
.B2(n_136),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_860),
.A2(n_1),
.B(n_5),
.C(n_6),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_967),
.B(n_135),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_976),
.A2(n_7),
.B(n_11),
.C(n_12),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_856),
.B(n_13),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_882),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_847),
.B(n_15),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_871),
.A2(n_127),
.B(n_125),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_885),
.A2(n_17),
.B(n_19),
.C(n_23),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_SL g1038 ( 
.A(n_891),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_909),
.A2(n_17),
.B(n_19),
.C(n_23),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_919),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_982),
.B(n_25),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_903),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_937),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_905),
.B(n_868),
.Y(n_1044)
);

O2A1O1Ixp5_ASAP7_75t_SL g1045 ( 
.A1(n_961),
.A2(n_26),
.B(n_29),
.C(n_30),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_970),
.B(n_31),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_820),
.A2(n_33),
.B(n_34),
.C(n_37),
.Y(n_1047)
);

AO22x1_ASAP7_75t_L g1048 ( 
.A1(n_864),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_946),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_866),
.A2(n_62),
.B(n_122),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_918),
.B(n_38),
.Y(n_1051)
);

INVx3_ASAP7_75t_SL g1052 ( 
.A(n_892),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_947),
.A2(n_39),
.B(n_40),
.C(n_41),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_870),
.B(n_42),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_824),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_867),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_920),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_917),
.B(n_76),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_846),
.B(n_94),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_871),
.A2(n_68),
.B(n_119),
.Y(n_1060)
);

NOR3xp33_ASAP7_75t_SL g1061 ( 
.A(n_931),
.B(n_43),
.C(n_47),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_923),
.B(n_50),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_950),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_825),
.Y(n_1064)
);

NOR3xp33_ASAP7_75t_SL g1065 ( 
.A(n_944),
.B(n_50),
.C(n_54),
.Y(n_1065)
);

AO32x2_ASAP7_75t_L g1066 ( 
.A1(n_984),
.A2(n_124),
.A3(n_65),
.B1(n_100),
.B2(n_109),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_SL g1067 ( 
.A(n_817),
.B(n_61),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_925),
.B(n_110),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_939),
.A2(n_111),
.B(n_877),
.C(n_886),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_951),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_846),
.B(n_941),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_811),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_814),
.B(n_822),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_965),
.A2(n_869),
.B(n_934),
.C(n_861),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_869),
.B(n_825),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_812),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_814),
.B(n_855),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_888),
.B(n_851),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_913),
.B(n_936),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_903),
.B(n_830),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_910),
.B(n_916),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_950),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_913),
.B(n_849),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_913),
.B(n_849),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_873),
.A2(n_875),
.B1(n_834),
.B2(n_822),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_842),
.A2(n_954),
.B(n_898),
.C(n_932),
.Y(n_1086)
);

BUFx8_ASAP7_75t_SL g1087 ( 
.A(n_910),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_871),
.A2(n_874),
.B(n_981),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_899),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_874),
.A2(n_942),
.B(n_945),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_910),
.A2(n_916),
.B1(n_971),
.B2(n_922),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_874),
.A2(n_942),
.B(n_945),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_916),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_834),
.B(n_889),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_964),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_SL g1096 ( 
.A(n_853),
.B(n_907),
.Y(n_1096)
);

OAI21xp33_ASAP7_75t_L g1097 ( 
.A1(n_854),
.A2(n_823),
.B(n_902),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_828),
.B(n_922),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_873),
.B(n_875),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_955),
.A2(n_972),
.B(n_933),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_955),
.A2(n_972),
.B(n_933),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_893),
.A2(n_930),
.B(n_895),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_971),
.A2(n_963),
.B1(n_894),
.B2(n_908),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_911),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_SL g1105 ( 
.A(n_907),
.B(n_984),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_948),
.B(n_914),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_823),
.B(n_821),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_836),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_953),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_876),
.A2(n_879),
.B(n_897),
.C(n_841),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_839),
.B(n_843),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_893),
.A2(n_930),
.B(n_895),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_883),
.B(n_915),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_837),
.B(n_841),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_964),
.Y(n_1115)
);

CKINVDCx11_ASAP7_75t_R g1116 ( 
.A(n_953),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_963),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_838),
.B(n_881),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_850),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_884),
.B(n_887),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_890),
.A2(n_973),
.B(n_983),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_926),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_912),
.B(n_829),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_900),
.A2(n_819),
.B(n_826),
.C(n_840),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_926),
.Y(n_1125)
);

OR2x6_ASAP7_75t_L g1126 ( 
.A(n_980),
.B(n_974),
.Y(n_1126)
);

AOI222xp33_ASAP7_75t_L g1127 ( 
.A1(n_848),
.A2(n_865),
.B1(n_863),
.B2(n_862),
.C1(n_816),
.C2(n_900),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1074),
.A2(n_1124),
.A3(n_989),
.B(n_1085),
.Y(n_1128)
);

OR2x6_ASAP7_75t_L g1129 ( 
.A(n_1071),
.B(n_980),
.Y(n_1129)
);

O2A1O1Ixp5_ASAP7_75t_SL g1130 ( 
.A1(n_1050),
.A2(n_927),
.B(n_921),
.C(n_904),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1027),
.A2(n_980),
.B1(n_977),
.B2(n_974),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_990),
.A2(n_845),
.B(n_940),
.Y(n_1132)
);

AO32x2_ASAP7_75t_L g1133 ( 
.A1(n_1085),
.A2(n_987),
.A3(n_989),
.B1(n_1045),
.B2(n_1095),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_993),
.B(n_983),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1101),
.A2(n_862),
.B(n_863),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1008),
.B(n_929),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_994),
.B(n_938),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1034),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_987),
.A2(n_929),
.A3(n_949),
.B(n_962),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1073),
.B(n_929),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1110),
.A2(n_929),
.B(n_949),
.Y(n_1141)
);

CKINVDCx14_ASAP7_75t_R g1142 ( 
.A(n_1116),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1102),
.A2(n_1112),
.B(n_1019),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1069),
.A2(n_831),
.B(n_978),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1080),
.B(n_938),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1090),
.A2(n_852),
.B(n_964),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1092),
.A2(n_964),
.B(n_926),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1055),
.Y(n_1148)
);

NAND2x1p5_ASAP7_75t_L g1149 ( 
.A(n_1095),
.B(n_1115),
.Y(n_1149)
);

AO32x2_ASAP7_75t_L g1150 ( 
.A1(n_1115),
.A2(n_1127),
.A3(n_1066),
.B1(n_1037),
.B2(n_988),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1056),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_985),
.B(n_1042),
.Y(n_1152)
);

AOI221x1_ASAP7_75t_L g1153 ( 
.A1(n_1050),
.A2(n_1047),
.B1(n_1078),
.B2(n_1097),
.C(n_1039),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_986),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1127),
.A2(n_1073),
.B(n_998),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_986),
.Y(n_1156)
);

BUFx12f_ASAP7_75t_L g1157 ( 
.A(n_1026),
.Y(n_1157)
);

OA21x2_ASAP7_75t_L g1158 ( 
.A1(n_1114),
.A2(n_992),
.B(n_1077),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1094),
.B(n_998),
.Y(n_1159)
);

INVx6_ASAP7_75t_L g1160 ( 
.A(n_1001),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1042),
.B(n_1096),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_997),
.A2(n_1105),
.B(n_1111),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_1109),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1006),
.A2(n_1007),
.B(n_1088),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1099),
.B(n_991),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1009),
.A2(n_1106),
.B(n_996),
.C(n_1013),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1081),
.B(n_1054),
.Y(n_1167)
);

INVxp67_ASAP7_75t_SL g1168 ( 
.A(n_1122),
.Y(n_1168)
);

BUFx2_ASAP7_75t_SL g1169 ( 
.A(n_1038),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_986),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1068),
.A2(n_1031),
.B(n_1058),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_SL g1172 ( 
.A(n_995),
.B(n_1053),
.C(n_1065),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_999),
.B(n_1107),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1051),
.B(n_1062),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1041),
.B(n_1091),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_994),
.B(n_1083),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1067),
.A2(n_1021),
.B(n_1020),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1005),
.A2(n_1029),
.B(n_1030),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1046),
.A2(n_1032),
.B(n_1123),
.C(n_1113),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1117),
.B(n_1093),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1118),
.A2(n_1120),
.B(n_1075),
.Y(n_1181)
);

INVx5_ASAP7_75t_L g1182 ( 
.A(n_1000),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1036),
.A2(n_1060),
.B(n_1103),
.Y(n_1183)
);

AO21x2_ASAP7_75t_L g1184 ( 
.A1(n_1012),
.A2(n_1044),
.B(n_1098),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1063),
.A2(n_1082),
.B(n_1089),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1093),
.B(n_1015),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1063),
.A2(n_1082),
.B(n_1104),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1119),
.B(n_1079),
.Y(n_1188)
);

AOI221x1_ASAP7_75t_L g1189 ( 
.A1(n_1057),
.A2(n_1035),
.B1(n_1033),
.B2(n_1025),
.C(n_1017),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1040),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1126),
.A2(n_1059),
.B1(n_1084),
.B2(n_1125),
.Y(n_1191)
);

AO21x2_ASAP7_75t_L g1192 ( 
.A1(n_1043),
.A2(n_1108),
.B(n_1049),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1067),
.A2(n_1126),
.B(n_1016),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_SL g1194 ( 
.A1(n_1059),
.A2(n_1122),
.B(n_1125),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1070),
.A2(n_1072),
.B(n_1076),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1002),
.A2(n_1004),
.B(n_1014),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1126),
.A2(n_1016),
.B(n_1122),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1022),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1003),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1066),
.A2(n_1125),
.B(n_988),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1000),
.B(n_1024),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1024),
.B(n_1064),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1064),
.B(n_1071),
.Y(n_1203)
);

AOI21xp33_ASAP7_75t_L g1204 ( 
.A1(n_1071),
.A2(n_1064),
.B(n_1066),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1061),
.B(n_1048),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1052),
.Y(n_1206)
);

INVx5_ASAP7_75t_L g1207 ( 
.A(n_1087),
.Y(n_1207)
);

O2A1O1Ixp5_ASAP7_75t_L g1208 ( 
.A1(n_1038),
.A2(n_957),
.B(n_901),
.C(n_670),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1011),
.A2(n_901),
.B(n_670),
.C(n_1086),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1080),
.B(n_870),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1074),
.A2(n_866),
.B(n_1102),
.Y(n_1211)
);

NOR2x1_ASAP7_75t_R g1212 ( 
.A(n_1023),
.B(n_520),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1086),
.A2(n_901),
.B(n_670),
.C(n_957),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1124),
.A2(n_901),
.B(n_1074),
.Y(n_1214)
);

AOI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1121),
.A2(n_990),
.B(n_866),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1080),
.B(n_870),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_985),
.B(n_795),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1018),
.B(n_1027),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1018),
.B(n_1027),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1018),
.B(n_1027),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_1026),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1048),
.A2(n_901),
.B1(n_670),
.B2(n_177),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1034),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1018),
.B(n_1027),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_985),
.A2(n_901),
.B1(n_858),
.B2(n_670),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1124),
.A2(n_901),
.B(n_1074),
.Y(n_1226)
);

BUFx10_ASAP7_75t_L g1227 ( 
.A(n_1023),
.Y(n_1227)
);

AOI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1121),
.A2(n_990),
.B(n_866),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_SL g1229 ( 
.A1(n_1053),
.A2(n_901),
.B(n_670),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_985),
.A2(n_901),
.B1(n_858),
.B2(n_670),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_990),
.A2(n_1101),
.B(n_1100),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_990),
.A2(n_1101),
.B(n_1100),
.Y(n_1232)
);

O2A1O1Ixp5_ASAP7_75t_L g1233 ( 
.A1(n_1069),
.A2(n_957),
.B(n_901),
.C(n_670),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_990),
.A2(n_1101),
.B(n_1100),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1121),
.A2(n_979),
.B(n_928),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_SL g1236 ( 
.A1(n_1053),
.A2(n_901),
.B(n_670),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_994),
.B(n_1083),
.Y(n_1237)
);

AOI21x1_ASAP7_75t_SL g1238 ( 
.A1(n_1078),
.A2(n_1107),
.B(n_1062),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1018),
.A2(n_901),
.B1(n_1027),
.B2(n_1010),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1018),
.B(n_1027),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_986),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1028),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1121),
.A2(n_979),
.B(n_928),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1018),
.B(n_1027),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_990),
.A2(n_1101),
.B(n_1100),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1124),
.A2(n_901),
.B(n_1074),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1034),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_986),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1074),
.A2(n_1124),
.A3(n_989),
.B(n_1085),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_990),
.A2(n_1101),
.B(n_1100),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1028),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1121),
.A2(n_979),
.B(n_928),
.Y(n_1252)
);

BUFx12f_ASAP7_75t_L g1253 ( 
.A(n_1116),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1018),
.B(n_1027),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1124),
.A2(n_901),
.B(n_1074),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1121),
.A2(n_979),
.B(n_928),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1018),
.B(n_1027),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1086),
.A2(n_901),
.B(n_670),
.C(n_957),
.Y(n_1258)
);

INVx3_ASAP7_75t_SL g1259 ( 
.A(n_1026),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1018),
.B(n_1027),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1074),
.A2(n_1124),
.A3(n_989),
.B(n_1085),
.Y(n_1261)
);

AO31x2_ASAP7_75t_L g1262 ( 
.A1(n_1074),
.A2(n_1124),
.A3(n_989),
.B(n_1085),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1063),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1121),
.A2(n_979),
.B(n_928),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_986),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1167),
.B(n_1210),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1253),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1164),
.A2(n_1132),
.B(n_1215),
.Y(n_1268)
);

NOR3xp33_ASAP7_75t_L g1269 ( 
.A(n_1229),
.B(n_1236),
.C(n_1208),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1228),
.A2(n_1232),
.B(n_1231),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1234),
.A2(n_1250),
.B(n_1245),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1160),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1160),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1138),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1225),
.B(n_1230),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1152),
.B(n_1188),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1135),
.A2(n_1243),
.B(n_1235),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1148),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1151),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1213),
.A2(n_1258),
.B(n_1233),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1252),
.A2(n_1264),
.B(n_1256),
.Y(n_1281)
);

BUFx2_ASAP7_75t_SL g1282 ( 
.A(n_1206),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1165),
.B(n_1224),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1223),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1224),
.B(n_1244),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_SL g1286 ( 
.A1(n_1209),
.A2(n_1166),
.B(n_1229),
.C(n_1236),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1247),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1183),
.A2(n_1146),
.B(n_1147),
.Y(n_1288)
);

CKINVDCx6p67_ASAP7_75t_R g1289 ( 
.A(n_1207),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1192),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1244),
.B(n_1257),
.Y(n_1291)
);

OA21x2_ASAP7_75t_L g1292 ( 
.A1(n_1171),
.A2(n_1155),
.B(n_1141),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1177),
.A2(n_1162),
.B(n_1141),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_SL g1294 ( 
.A1(n_1178),
.A2(n_1204),
.B(n_1172),
.C(n_1136),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1216),
.B(n_1180),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1239),
.B(n_1174),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1159),
.A2(n_1246),
.B(n_1255),
.Y(n_1297)
);

AOI21xp33_ASAP7_75t_L g1298 ( 
.A1(n_1178),
.A2(n_1174),
.B(n_1175),
.Y(n_1298)
);

NAND2x1p5_ASAP7_75t_L g1299 ( 
.A(n_1182),
.B(n_1161),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1130),
.A2(n_1238),
.B(n_1187),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1163),
.Y(n_1301)
);

NOR2xp67_ASAP7_75t_L g1302 ( 
.A(n_1242),
.B(n_1251),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1190),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1185),
.A2(n_1200),
.B(n_1144),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1257),
.B(n_1260),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1217),
.B(n_1173),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1181),
.A2(n_1211),
.B(n_1226),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1211),
.A2(n_1214),
.B(n_1226),
.Y(n_1308)
);

INVx4_ASAP7_75t_L g1309 ( 
.A(n_1182),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1239),
.B(n_1218),
.Y(n_1310)
);

AO21x2_ASAP7_75t_L g1311 ( 
.A1(n_1214),
.A2(n_1246),
.B(n_1204),
.Y(n_1311)
);

CKINVDCx11_ASAP7_75t_R g1312 ( 
.A(n_1259),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1260),
.B(n_1219),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1136),
.A2(n_1140),
.B(n_1196),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1140),
.A2(n_1158),
.B(n_1131),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1175),
.A2(n_1173),
.B1(n_1205),
.B2(n_1240),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1195),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1199),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1220),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1254),
.B(n_1222),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1222),
.A2(n_1131),
.B(n_1179),
.C(n_1134),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1158),
.A2(n_1191),
.B(n_1153),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1128),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1176),
.B(n_1237),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1149),
.A2(n_1189),
.B(n_1186),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1201),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1201),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1149),
.A2(n_1263),
.B(n_1203),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1145),
.B(n_1221),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1137),
.A2(n_1194),
.B(n_1168),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1133),
.A2(n_1128),
.B(n_1249),
.Y(n_1331)
);

CKINVDCx11_ASAP7_75t_R g1332 ( 
.A(n_1227),
.Y(n_1332)
);

NOR2xp67_ASAP7_75t_L g1333 ( 
.A(n_1157),
.B(n_1265),
.Y(n_1333)
);

NAND2xp33_ASAP7_75t_R g1334 ( 
.A(n_1129),
.B(n_1203),
.Y(n_1334)
);

OR2x6_ASAP7_75t_L g1335 ( 
.A(n_1129),
.B(n_1169),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1182),
.A2(n_1202),
.B1(n_1207),
.B2(n_1265),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_SL g1337 ( 
.A(n_1212),
.B(n_1227),
.Y(n_1337)
);

AO32x2_ASAP7_75t_L g1338 ( 
.A1(n_1133),
.A2(n_1262),
.A3(n_1261),
.B1(n_1249),
.B2(n_1150),
.Y(n_1338)
);

NAND3xp33_ASAP7_75t_SL g1339 ( 
.A(n_1202),
.B(n_1142),
.C(n_1156),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1154),
.Y(n_1340)
);

INVx5_ASAP7_75t_L g1341 ( 
.A(n_1154),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1139),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1184),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1133),
.A2(n_1262),
.B(n_1261),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1184),
.A2(n_1207),
.B1(n_1198),
.B2(n_1249),
.Y(n_1345)
);

INVx5_ASAP7_75t_L g1346 ( 
.A(n_1170),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1170),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1241),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1262),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1261),
.B(n_1241),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1248),
.B(n_1156),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1139),
.A2(n_1150),
.B(n_1248),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1160),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1180),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1138),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1138),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1263),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1164),
.A2(n_1132),
.B(n_1215),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1138),
.Y(n_1359)
);

NAND2x1p5_ASAP7_75t_L g1360 ( 
.A(n_1182),
.B(n_817),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1225),
.A2(n_858),
.B1(n_901),
.B2(n_1230),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1167),
.B(n_1210),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1164),
.A2(n_1132),
.B(n_1215),
.Y(n_1363)
);

CKINVDCx6p67_ASAP7_75t_R g1364 ( 
.A(n_1207),
.Y(n_1364)
);

INVxp67_ASAP7_75t_SL g1365 ( 
.A(n_1224),
.Y(n_1365)
);

OR2x6_ASAP7_75t_L g1366 ( 
.A(n_1193),
.B(n_1197),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_SL g1367 ( 
.A1(n_1193),
.A2(n_1197),
.B(n_1178),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1253),
.Y(n_1368)
);

CKINVDCx14_ASAP7_75t_R g1369 ( 
.A(n_1142),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1138),
.Y(n_1370)
);

BUFx12f_ASAP7_75t_L g1371 ( 
.A(n_1253),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1213),
.A2(n_1258),
.B(n_1233),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1172),
.A2(n_901),
.B1(n_1226),
.B2(n_1214),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1164),
.A2(n_1132),
.B(n_1215),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1222),
.A2(n_901),
.B1(n_995),
.B2(n_858),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1225),
.B(n_901),
.Y(n_1376)
);

AOI21xp33_ASAP7_75t_L g1377 ( 
.A1(n_1229),
.A2(n_901),
.B(n_670),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1143),
.A2(n_1232),
.B(n_1231),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1176),
.B(n_1237),
.Y(n_1379)
);

AOI221xp5_ASAP7_75t_L g1380 ( 
.A1(n_1229),
.A2(n_901),
.B1(n_858),
.B2(n_1236),
.C(n_670),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1164),
.A2(n_1132),
.B(n_1215),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1263),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1165),
.B(n_901),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1164),
.A2(n_1132),
.B(n_1215),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1163),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1221),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1383),
.B(n_1283),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_SL g1388 ( 
.A1(n_1365),
.A2(n_1380),
.B(n_1376),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1313),
.B(n_1285),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1321),
.A2(n_1310),
.B(n_1305),
.Y(n_1390)
);

NOR2xp67_ASAP7_75t_L g1391 ( 
.A(n_1339),
.B(n_1385),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1291),
.B(n_1319),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1322),
.A2(n_1281),
.B(n_1280),
.Y(n_1393)
);

A2O1A1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1376),
.A2(n_1275),
.B(n_1297),
.C(n_1377),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1274),
.Y(n_1395)
);

O2A1O1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1286),
.A2(n_1321),
.B(n_1275),
.C(n_1372),
.Y(n_1396)
);

BUFx10_ASAP7_75t_L g1397 ( 
.A(n_1267),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1354),
.B(n_1306),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1310),
.A2(n_1296),
.B(n_1330),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1319),
.B(n_1316),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1366),
.B(n_1328),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1341),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1290),
.Y(n_1403)
);

O2A1O1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1286),
.A2(n_1298),
.B(n_1269),
.C(n_1296),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1375),
.A2(n_1361),
.B1(n_1373),
.B2(n_1320),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1373),
.A2(n_1308),
.B(n_1316),
.C(n_1322),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1295),
.B(n_1266),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1281),
.A2(n_1277),
.B(n_1307),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1276),
.B(n_1326),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1345),
.A2(n_1386),
.B1(n_1299),
.B2(n_1366),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1327),
.B(n_1329),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1335),
.A2(n_1379),
.B1(n_1302),
.B2(n_1301),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1362),
.B(n_1324),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1379),
.B(n_1303),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1318),
.B(n_1340),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1289),
.A2(n_1364),
.B1(n_1359),
.B2(n_1370),
.Y(n_1417)
);

BUFx2_ASAP7_75t_SL g1418 ( 
.A(n_1272),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1289),
.A2(n_1364),
.B1(n_1287),
.B2(n_1355),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_SL g1420 ( 
.A1(n_1360),
.A2(n_1309),
.B(n_1336),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1270),
.A2(n_1293),
.B(n_1300),
.Y(n_1421)
);

AOI21x1_ASAP7_75t_SL g1422 ( 
.A1(n_1351),
.A2(n_1332),
.B(n_1369),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1309),
.A2(n_1360),
.B(n_1311),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1284),
.B(n_1356),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1328),
.B(n_1350),
.Y(n_1425)
);

AOI221x1_ASAP7_75t_SL g1426 ( 
.A1(n_1333),
.A2(n_1348),
.B1(n_1343),
.B2(n_1323),
.C(n_1349),
.Y(n_1426)
);

OAI31xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1325),
.A2(n_1367),
.A3(n_1344),
.B(n_1352),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1357),
.B(n_1382),
.Y(n_1428)
);

NAND4xp25_ASAP7_75t_L g1429 ( 
.A(n_1337),
.B(n_1353),
.C(n_1272),
.D(n_1294),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1268),
.A2(n_1384),
.B(n_1358),
.Y(n_1430)
);

AND2x2_ASAP7_75t_SL g1431 ( 
.A(n_1292),
.B(n_1331),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1282),
.A2(n_1353),
.B1(n_1273),
.B2(n_1309),
.Y(n_1432)
);

NOR2xp67_ASAP7_75t_L g1433 ( 
.A(n_1347),
.B(n_1267),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1292),
.A2(n_1378),
.B(n_1331),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1358),
.A2(n_1381),
.B(n_1374),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1341),
.B(n_1346),
.Y(n_1436)
);

AOI21x1_ASAP7_75t_SL g1437 ( 
.A1(n_1312),
.A2(n_1334),
.B(n_1371),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1341),
.A2(n_1346),
.B1(n_1368),
.B2(n_1292),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1346),
.B(n_1314),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1334),
.A2(n_1312),
.B1(n_1368),
.B2(n_1371),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1315),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1342),
.A2(n_1331),
.B1(n_1317),
.B2(n_1338),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1342),
.A2(n_1338),
.B1(n_1315),
.B2(n_1304),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1344),
.B(n_1304),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1288),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1338),
.B(n_1288),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1338),
.B(n_1363),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_SL g1448 ( 
.A1(n_1271),
.A2(n_1193),
.B(n_1213),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1295),
.B(n_1266),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1272),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1297),
.A2(n_1258),
.B(n_1213),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1354),
.B(n_1306),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1297),
.A2(n_1258),
.B(n_1213),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1295),
.B(n_1266),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1274),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1274),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1375),
.A2(n_1222),
.B1(n_1230),
.B2(n_1225),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1383),
.B(n_1283),
.Y(n_1458)
);

OR2x6_ASAP7_75t_L g1459 ( 
.A(n_1366),
.B(n_1193),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1295),
.B(n_1266),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1354),
.B(n_1306),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1383),
.B(n_1283),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1383),
.B(n_1283),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1295),
.B(n_1266),
.Y(n_1464)
);

AND2x4_ASAP7_75t_SL g1465 ( 
.A(n_1354),
.B(n_1366),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1295),
.B(n_1266),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1365),
.A2(n_1193),
.B(n_1213),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1274),
.Y(n_1468)
);

INVx1_ASAP7_75t_SL g1469 ( 
.A(n_1386),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1375),
.A2(n_1222),
.B1(n_1230),
.B2(n_1225),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1312),
.Y(n_1471)
);

AOI221x1_ASAP7_75t_SL g1472 ( 
.A1(n_1376),
.A2(n_622),
.B1(n_901),
.B2(n_1377),
.C(n_728),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1375),
.A2(n_1222),
.B1(n_1230),
.B2(n_1225),
.Y(n_1473)
);

O2A1O1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1377),
.A2(n_901),
.B(n_1236),
.C(n_1229),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1354),
.B(n_1306),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1441),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1446),
.B(n_1447),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1400),
.B(n_1394),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1405),
.B(n_1396),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1431),
.B(n_1425),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1444),
.B(n_1443),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1457),
.A2(n_1473),
.B1(n_1470),
.B2(n_1451),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1431),
.B(n_1425),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1388),
.B(n_1394),
.Y(n_1484)
);

INVx4_ASAP7_75t_L g1485 ( 
.A(n_1459),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1434),
.A2(n_1406),
.B(n_1453),
.Y(n_1486)
);

INVx4_ASAP7_75t_L g1487 ( 
.A(n_1459),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1459),
.B(n_1448),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1442),
.B(n_1393),
.Y(n_1489)
);

NAND2x1_ASAP7_75t_L g1490 ( 
.A(n_1399),
.B(n_1423),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1403),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1401),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1395),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1408),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1441),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1427),
.B(n_1445),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1445),
.B(n_1421),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1421),
.B(n_1398),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1439),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1421),
.B(n_1455),
.Y(n_1500)
);

OA21x2_ASAP7_75t_L g1501 ( 
.A1(n_1456),
.A2(n_1468),
.B(n_1428),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1416),
.Y(n_1502)
);

AO21x2_ASAP7_75t_L g1503 ( 
.A1(n_1399),
.A2(n_1438),
.B(n_1474),
.Y(n_1503)
);

OAI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1387),
.A2(n_1463),
.B1(n_1462),
.B2(n_1458),
.Y(n_1504)
);

AO21x2_ASAP7_75t_L g1505 ( 
.A1(n_1467),
.A2(n_1423),
.B(n_1404),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1389),
.B(n_1392),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1426),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1424),
.Y(n_1508)
);

AO21x2_ASAP7_75t_L g1509 ( 
.A1(n_1467),
.A2(n_1390),
.B(n_1410),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1390),
.B(n_1409),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1465),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1472),
.B(n_1475),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1452),
.B(n_1461),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1477),
.B(n_1435),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1476),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1500),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1494),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1504),
.B(n_1419),
.Y(n_1518)
);

OAI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1482),
.A2(n_1429),
.B1(n_1440),
.B2(n_1391),
.C(n_1417),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1500),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1482),
.A2(n_1414),
.B1(n_1412),
.B2(n_1413),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1500),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1499),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1495),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1480),
.B(n_1430),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1491),
.Y(n_1526)
);

INVx4_ASAP7_75t_L g1527 ( 
.A(n_1488),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1491),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1480),
.B(n_1430),
.Y(n_1529)
);

INVx5_ASAP7_75t_L g1530 ( 
.A(n_1488),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1501),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1489),
.B(n_1411),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1497),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1504),
.B(n_1432),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1532),
.B(n_1513),
.Y(n_1535)
);

NAND2xp33_ASAP7_75t_R g1536 ( 
.A(n_1518),
.B(n_1484),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1526),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1523),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1526),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1525),
.B(n_1483),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1526),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1532),
.B(n_1516),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1532),
.B(n_1513),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1528),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1519),
.A2(n_1479),
.B1(n_1484),
.B2(n_1478),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1517),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1532),
.B(n_1499),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1516),
.B(n_1498),
.Y(n_1548)
);

NOR2x1_ASAP7_75t_L g1549 ( 
.A(n_1524),
.B(n_1490),
.Y(n_1549)
);

OAI33xp33_ASAP7_75t_L g1550 ( 
.A1(n_1523),
.A2(n_1512),
.A3(n_1478),
.B1(n_1506),
.B2(n_1513),
.B3(n_1510),
.Y(n_1550)
);

OAI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1519),
.A2(n_1479),
.B1(n_1490),
.B2(n_1510),
.Y(n_1551)
);

AOI33xp33_ASAP7_75t_L g1552 ( 
.A1(n_1533),
.A2(n_1469),
.A3(n_1496),
.B1(n_1460),
.B2(n_1407),
.B3(n_1466),
.Y(n_1552)
);

AOI221xp5_ASAP7_75t_L g1553 ( 
.A1(n_1518),
.A2(n_1512),
.B1(n_1507),
.B2(n_1499),
.C(n_1506),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1517),
.Y(n_1554)
);

OR2x6_ASAP7_75t_L g1555 ( 
.A(n_1527),
.B(n_1488),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1524),
.Y(n_1556)
);

INVx4_ASAP7_75t_L g1557 ( 
.A(n_1530),
.Y(n_1557)
);

OAI211xp5_ASAP7_75t_L g1558 ( 
.A1(n_1534),
.A2(n_1507),
.B(n_1496),
.C(n_1489),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1519),
.A2(n_1509),
.B1(n_1503),
.B2(n_1505),
.Y(n_1559)
);

AOI221xp5_ASAP7_75t_L g1560 ( 
.A1(n_1534),
.A2(n_1496),
.B1(n_1486),
.B2(n_1508),
.C(n_1502),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1516),
.B(n_1498),
.Y(n_1561)
);

NOR4xp25_ASAP7_75t_SL g1562 ( 
.A(n_1515),
.B(n_1471),
.C(n_1511),
.D(n_1493),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1524),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1521),
.A2(n_1488),
.B1(n_1487),
.B2(n_1485),
.Y(n_1564)
);

NAND4xp25_ASAP7_75t_L g1565 ( 
.A(n_1521),
.B(n_1481),
.C(n_1449),
.D(n_1464),
.Y(n_1565)
);

OA222x2_ASAP7_75t_L g1566 ( 
.A1(n_1524),
.A2(n_1488),
.B1(n_1489),
.B2(n_1481),
.C1(n_1492),
.C2(n_1509),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1530),
.A2(n_1509),
.B1(n_1505),
.B2(n_1503),
.Y(n_1567)
);

NAND4xp25_ASAP7_75t_L g1568 ( 
.A(n_1521),
.B(n_1481),
.C(n_1454),
.D(n_1415),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1546),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1545),
.B(n_1471),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1537),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1546),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1539),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1541),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1544),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1549),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1556),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1554),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1554),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1540),
.B(n_1525),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1556),
.Y(n_1581)
);

NOR3xp33_ASAP7_75t_L g1582 ( 
.A(n_1551),
.B(n_1433),
.C(n_1487),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1542),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1536),
.Y(n_1584)
);

AOI21xp33_ASAP7_75t_L g1585 ( 
.A1(n_1536),
.A2(n_1509),
.B(n_1486),
.Y(n_1585)
);

BUFx8_ASAP7_75t_L g1586 ( 
.A(n_1558),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1557),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1542),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1538),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1548),
.Y(n_1590)
);

NOR2x1p5_ASAP7_75t_L g1591 ( 
.A(n_1565),
.B(n_1527),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1552),
.B(n_1553),
.Y(n_1592)
);

NOR2x1p5_ASAP7_75t_L g1593 ( 
.A(n_1568),
.B(n_1527),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1547),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1535),
.B(n_1520),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1543),
.B(n_1520),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1548),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1561),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1561),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1584),
.B(n_1560),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1580),
.B(n_1566),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1576),
.B(n_1557),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1583),
.B(n_1533),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1584),
.B(n_1552),
.Y(n_1604)
);

AND2x4_ASAP7_75t_SL g1605 ( 
.A(n_1582),
.B(n_1557),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1571),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1580),
.B(n_1563),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1571),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1574),
.Y(n_1609)
);

OAI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1592),
.A2(n_1559),
.B1(n_1567),
.B2(n_1564),
.C(n_1488),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1574),
.Y(n_1611)
);

CKINVDCx14_ASAP7_75t_R g1612 ( 
.A(n_1570),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1589),
.B(n_1522),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1576),
.B(n_1529),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1594),
.B(n_1529),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1589),
.B(n_1533),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1583),
.B(n_1498),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_1587),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1594),
.B(n_1529),
.Y(n_1619)
);

NAND2xp33_ASAP7_75t_SL g1620 ( 
.A(n_1593),
.B(n_1562),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1569),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1581),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1569),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1581),
.B(n_1529),
.Y(n_1624)
);

NOR3xp33_ASAP7_75t_L g1625 ( 
.A(n_1585),
.B(n_1550),
.C(n_1450),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1573),
.Y(n_1626)
);

BUFx3_ASAP7_75t_L g1627 ( 
.A(n_1577),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1587),
.B(n_1555),
.Y(n_1628)
);

NAND3xp33_ASAP7_75t_L g1629 ( 
.A(n_1586),
.B(n_1559),
.C(n_1531),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1587),
.B(n_1555),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1577),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1573),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1587),
.B(n_1555),
.Y(n_1633)
);

AND2x4_ASAP7_75t_SL g1634 ( 
.A(n_1582),
.B(n_1555),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1569),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1590),
.B(n_1514),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1575),
.Y(n_1637)
);

NOR4xp25_ASAP7_75t_L g1638 ( 
.A(n_1600),
.B(n_1585),
.C(n_1581),
.D(n_1588),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1604),
.B(n_1591),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1604),
.B(n_1599),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1631),
.B(n_1591),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1600),
.B(n_1590),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1631),
.B(n_1593),
.Y(n_1643)
);

INVxp67_ASAP7_75t_SL g1644 ( 
.A(n_1609),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1627),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1627),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1616),
.B(n_1595),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1609),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1625),
.B(n_1627),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1629),
.A2(n_1620),
.B1(n_1625),
.B2(n_1610),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1622),
.B(n_1577),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1618),
.Y(n_1652)
);

NOR2x1_ASAP7_75t_SL g1653 ( 
.A(n_1629),
.B(n_1618),
.Y(n_1653)
);

OAI21xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1601),
.A2(n_1599),
.B(n_1598),
.Y(n_1654)
);

INVx2_ASAP7_75t_SL g1655 ( 
.A(n_1618),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1612),
.A2(n_1486),
.B(n_1505),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1628),
.B(n_1630),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1626),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1622),
.B(n_1597),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1626),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1632),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1610),
.A2(n_1602),
.B(n_1616),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1605),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1628),
.B(n_1597),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1632),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1624),
.B(n_1598),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1624),
.B(n_1595),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1637),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1637),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1605),
.B(n_1397),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1605),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1613),
.B(n_1596),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1606),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1644),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1642),
.B(n_1606),
.Y(n_1675)
);

AND3x1_ASAP7_75t_L g1676 ( 
.A(n_1638),
.B(n_1601),
.C(n_1628),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1653),
.B(n_1634),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1657),
.B(n_1634),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1651),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1650),
.A2(n_1586),
.B1(n_1634),
.B2(n_1486),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1655),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1655),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1652),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1652),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1645),
.B(n_1607),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1644),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1657),
.B(n_1646),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1651),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1658),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1651),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1648),
.Y(n_1691)
);

CKINVDCx16_ASAP7_75t_R g1692 ( 
.A(n_1663),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1660),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1649),
.A2(n_1586),
.B1(n_1488),
.B2(n_1611),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1661),
.Y(n_1695)
);

NOR2x1_ASAP7_75t_L g1696 ( 
.A(n_1673),
.B(n_1608),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1665),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1668),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1639),
.A2(n_1656),
.B1(n_1662),
.B2(n_1642),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1676),
.A2(n_1671),
.B1(n_1670),
.B2(n_1586),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1687),
.Y(n_1701)
);

NAND2xp33_ASAP7_75t_L g1702 ( 
.A(n_1677),
.B(n_1680),
.Y(n_1702)
);

AOI21xp33_ASAP7_75t_L g1703 ( 
.A1(n_1699),
.A2(n_1640),
.B(n_1670),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1692),
.B(n_1664),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1691),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1692),
.B(n_1640),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1676),
.A2(n_1699),
.B1(n_1685),
.B2(n_1694),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1691),
.Y(n_1708)
);

NOR3xp33_ASAP7_75t_L g1709 ( 
.A(n_1679),
.B(n_1643),
.C(n_1641),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1696),
.A2(n_1659),
.B(n_1654),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1687),
.B(n_1664),
.Y(n_1711)
);

NAND4xp25_ASAP7_75t_L g1712 ( 
.A(n_1696),
.B(n_1669),
.C(n_1666),
.D(n_1647),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1674),
.Y(n_1713)
);

OA21x2_ASAP7_75t_L g1714 ( 
.A1(n_1674),
.A2(n_1611),
.B(n_1608),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1686),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1686),
.Y(n_1716)
);

O2A1O1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1694),
.A2(n_1602),
.B(n_1630),
.C(n_1633),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1677),
.A2(n_1602),
.B1(n_1667),
.B2(n_1630),
.C(n_1633),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1690),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1701),
.B(n_1690),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1704),
.B(n_1690),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1719),
.B(n_1688),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1707),
.A2(n_1678),
.B1(n_1586),
.B2(n_1688),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1705),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1708),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1706),
.B(n_1688),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1709),
.B(n_1688),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1711),
.B(n_1678),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1714),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1714),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1713),
.Y(n_1731)
);

OAI21x1_ASAP7_75t_L g1732 ( 
.A1(n_1729),
.A2(n_1710),
.B(n_1682),
.Y(n_1732)
);

NOR3xp33_ASAP7_75t_L g1733 ( 
.A(n_1726),
.B(n_1702),
.C(n_1703),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1723),
.A2(n_1700),
.B(n_1727),
.Y(n_1734)
);

OAI211xp5_ASAP7_75t_L g1735 ( 
.A1(n_1730),
.A2(n_1712),
.B(n_1721),
.C(n_1720),
.Y(n_1735)
);

AND4x1_ASAP7_75t_L g1736 ( 
.A(n_1720),
.B(n_1717),
.C(n_1718),
.D(n_1716),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1728),
.B(n_1712),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1722),
.B(n_1715),
.Y(n_1738)
);

OAI31xp33_ASAP7_75t_L g1739 ( 
.A1(n_1728),
.A2(n_1681),
.A3(n_1675),
.B(n_1682),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1722),
.B(n_1675),
.Y(n_1740)
);

NAND4xp25_ASAP7_75t_L g1741 ( 
.A(n_1724),
.B(n_1698),
.C(n_1697),
.D(n_1695),
.Y(n_1741)
);

AOI221x1_ASAP7_75t_L g1742 ( 
.A1(n_1725),
.A2(n_1682),
.B1(n_1684),
.B2(n_1683),
.C(n_1698),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1733),
.A2(n_1683),
.B1(n_1684),
.B2(n_1731),
.Y(n_1743)
);

AOI221x1_ASAP7_75t_L g1744 ( 
.A1(n_1734),
.A2(n_1731),
.B1(n_1683),
.B2(n_1684),
.C(n_1697),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1732),
.A2(n_1693),
.B(n_1689),
.C(n_1695),
.Y(n_1745)
);

OA22x2_ASAP7_75t_L g1746 ( 
.A1(n_1735),
.A2(n_1693),
.B1(n_1689),
.B2(n_1602),
.Y(n_1746)
);

OAI21xp33_ASAP7_75t_L g1747 ( 
.A1(n_1737),
.A2(n_1633),
.B(n_1614),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1740),
.A2(n_1614),
.B1(n_1607),
.B2(n_1635),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1738),
.A2(n_1614),
.B1(n_1635),
.B2(n_1623),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1742),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1746),
.B(n_1739),
.Y(n_1751)
);

NAND2x1_ASAP7_75t_L g1752 ( 
.A(n_1750),
.B(n_1621),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1743),
.B(n_1736),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1748),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1745),
.Y(n_1755)
);

NAND3xp33_ASAP7_75t_L g1756 ( 
.A(n_1744),
.B(n_1741),
.C(n_1672),
.Y(n_1756)
);

NAND3xp33_ASAP7_75t_L g1757 ( 
.A(n_1747),
.B(n_1623),
.C(n_1621),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1749),
.B(n_1615),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1751),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1752),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1753),
.A2(n_1635),
.B1(n_1623),
.B2(n_1621),
.Y(n_1761)
);

NOR2x1_ASAP7_75t_L g1762 ( 
.A(n_1755),
.B(n_1756),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1754),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1759),
.B(n_1763),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1760),
.B(n_1758),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1761),
.B(n_1757),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1764),
.B(n_1762),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1767),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1765),
.B1(n_1766),
.B2(n_1397),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1768),
.A2(n_1397),
.B1(n_1418),
.B2(n_1450),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1769),
.B(n_1613),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1770),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1771),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1772),
.Y(n_1774)
);

XOR2x2_ASAP7_75t_L g1775 ( 
.A(n_1774),
.B(n_1422),
.Y(n_1775)
);

AO221x2_ASAP7_75t_L g1776 ( 
.A1(n_1775),
.A2(n_1773),
.B1(n_1572),
.B2(n_1578),
.C(n_1579),
.Y(n_1776)
);

OAI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1776),
.A2(n_1603),
.B(n_1617),
.Y(n_1777)
);

XNOR2xp5_ASAP7_75t_L g1778 ( 
.A(n_1777),
.B(n_1437),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1778),
.A2(n_1619),
.B1(n_1615),
.B2(n_1636),
.Y(n_1779)
);

AOI211xp5_ASAP7_75t_L g1780 ( 
.A1(n_1779),
.A2(n_1420),
.B(n_1402),
.C(n_1436),
.Y(n_1780)
);


endmodule