module fake_jpeg_15789_n_215 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_215);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_7),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_1),
.C(n_3),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_43),
.B(n_45),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_15),
.B(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_4),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_55),
.Y(n_67)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_27),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_57),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_32),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_63),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_23),
.B1(n_36),
.B2(n_25),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_64),
.B1(n_70),
.B2(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_35),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_23),
.B1(n_26),
.B2(n_30),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_18),
.B1(n_30),
.B2(n_34),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_66),
.A2(n_87),
.B1(n_10),
.B2(n_11),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_69),
.B(n_74),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_19),
.B1(n_36),
.B2(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_80),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_42),
.B(n_46),
.C(n_39),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_72),
.B1(n_61),
.B2(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_82),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_42),
.A2(n_19),
.B1(n_29),
.B2(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_29),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_37),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_24),
.B1(n_5),
.B2(n_9),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_4),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_69),
.B(n_74),
.C(n_76),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_90),
.B(n_57),
.Y(n_96)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_111),
.B1(n_110),
.B2(n_101),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_98),
.B(n_93),
.Y(n_140)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_63),
.A2(n_86),
.B1(n_91),
.B2(n_64),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_109),
.B1(n_113),
.B2(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_41),
.B1(n_24),
.B2(n_11),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

BUFx2_ASAP7_75t_SL g112 ( 
.A(n_81),
.Y(n_112)
);

CKINVDCx10_ASAP7_75t_R g129 ( 
.A(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_12),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_122),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_115),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_67),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_118),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_75),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_73),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_108),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_72),
.A3(n_73),
.B1(n_75),
.B2(n_79),
.C1(n_68),
.C2(n_61),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_133),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_94),
.B(n_119),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_137),
.B(n_140),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_73),
.B1(n_68),
.B2(n_79),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_130),
.B1(n_145),
.B2(n_146),
.Y(n_155)
);

AO22x2_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_105),
.B1(n_94),
.B2(n_103),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_124),
.B1(n_130),
.B2(n_138),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_111),
.B(n_122),
.Y(n_137)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_93),
.A2(n_122),
.B1(n_97),
.B2(n_95),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_136),
.B(n_150),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_102),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_147),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_164),
.Y(n_179)
);

AO21x1_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_168),
.B(n_162),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_137),
.C(n_138),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_157),
.C(n_160),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_145),
.B1(n_148),
.B2(n_128),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_159),
.B1(n_162),
.B2(n_167),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_149),
.C(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_165),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_130),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_161),
.A2(n_162),
.B(n_167),
.Y(n_184)
);

AND2x4_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_129),
.Y(n_162)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_170),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_126),
.B(n_125),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_182),
.B(n_181),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_143),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_176),
.C(n_168),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_141),
.C(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_158),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_180),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_163),
.C(n_179),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_185),
.A2(n_155),
.B1(n_169),
.B2(n_165),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_177),
.A2(n_159),
.B1(n_156),
.B2(n_155),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_186),
.A2(n_185),
.B1(n_172),
.B2(n_176),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_151),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_190),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_193),
.B1(n_175),
.B2(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_183),
.Y(n_198)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_200),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_184),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_197),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_188),
.B1(n_186),
.B2(n_193),
.Y(n_205)
);

AOI322xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_192),
.A3(n_196),
.B1(n_188),
.B2(n_187),
.C1(n_190),
.C2(n_194),
.Y(n_206)
);

NOR2x1_ASAP7_75t_R g210 ( 
.A(n_206),
.B(n_201),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_205),
.B(n_202),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_211),
.C(n_204),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_207),
.A2(n_201),
.B(n_208),
.Y(n_211)
);

NAND2xp33_ASAP7_75t_R g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_209),
.Y(n_215)
);


endmodule