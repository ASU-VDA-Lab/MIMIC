module fake_jpeg_15182_n_335 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_47),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_19),
.Y(n_55)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_24),
.B1(n_22),
.B2(n_20),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_59),
.B1(n_64),
.B2(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_55),
.B(n_43),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_24),
.B1(n_22),
.B2(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_30),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_62),
.Y(n_73)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_24),
.B1(n_22),
.B2(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_37),
.A2(n_20),
.B1(n_26),
.B2(n_35),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_98),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_49),
.B1(n_47),
.B2(n_46),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_101),
.B1(n_19),
.B2(n_33),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_57),
.A2(n_43),
.B1(n_26),
.B2(n_47),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_69),
.B1(n_23),
.B2(n_32),
.Y(n_112)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_91),
.Y(n_114)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_49),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_95),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_48),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_19),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_39),
.B(n_40),
.C(n_28),
.D(n_34),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_39),
.C(n_40),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_60),
.B(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_23),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_39),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_21),
.B1(n_27),
.B2(n_33),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_39),
.C(n_38),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_39),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_77),
.A2(n_41),
.B1(n_48),
.B2(n_50),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_129),
.B1(n_31),
.B2(n_27),
.Y(n_135)
);

NAND2xp67_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_91),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_111),
.B(n_34),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_118),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_40),
.C(n_78),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_68),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_93),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_41),
.B(n_40),
.C(n_21),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_122),
.Y(n_140)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_78),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_128),
.Y(n_150)
);

INVx5_ASAP7_75t_SL g125 ( 
.A(n_87),
.Y(n_125)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_25),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_50),
.B1(n_31),
.B2(n_33),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_25),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_75),
.A2(n_31),
.B1(n_27),
.B2(n_21),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_136),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_108),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_102),
.B1(n_99),
.B2(n_94),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_146),
.B1(n_148),
.B2(n_119),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_111),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_105),
.A2(n_93),
.B1(n_76),
.B2(n_79),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_108),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_153),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_111),
.B1(n_113),
.B2(n_129),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_155),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_151),
.A2(n_107),
.B(n_124),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_115),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_42),
.C(n_18),
.Y(n_155)
);

AO22x1_ASAP7_75t_SL g156 ( 
.A1(n_110),
.A2(n_90),
.B1(n_85),
.B2(n_100),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_127),
.B1(n_125),
.B2(n_122),
.Y(n_171)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_137),
.A3(n_148),
.B1(n_144),
.B2(n_140),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_158),
.B(n_177),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_28),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_161),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_107),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_162),
.B(n_174),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_141),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_114),
.B(n_132),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_167),
.A2(n_175),
.B(n_180),
.Y(n_204)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_171),
.A2(n_153),
.B1(n_136),
.B2(n_125),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

AO21x1_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_143),
.B(n_117),
.Y(n_191)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_104),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_118),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_138),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_178),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_181),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_177),
.C(n_159),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_207),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_152),
.B1(n_155),
.B2(n_134),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_185),
.B1(n_194),
.B2(n_200),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_175),
.A2(n_134),
.B1(n_156),
.B2(n_147),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_166),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_143),
.A3(n_104),
.B1(n_132),
.B2(n_115),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_190),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_192),
.B(n_210),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_83),
.B1(n_106),
.B2(n_103),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_106),
.B1(n_83),
.B2(n_120),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_202),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_80),
.B1(n_117),
.B2(n_123),
.Y(n_200)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_71),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_168),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_161),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_80),
.B1(n_103),
.B2(n_97),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_163),
.B1(n_172),
.B2(n_170),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_42),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_209),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_157),
.B(n_71),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_167),
.B(n_28),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_207),
.Y(n_233)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_210),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_219),
.B(n_221),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_195),
.B1(n_190),
.B2(n_186),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_229),
.B1(n_222),
.B2(n_230),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_233),
.Y(n_239)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_227),
.A2(n_221),
.B(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_231),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_169),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_163),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_235),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_185),
.A2(n_182),
.B1(n_97),
.B2(n_95),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_SL g252 ( 
.A1(n_234),
.A2(n_194),
.B(n_214),
.C(n_224),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_197),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_42),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_183),
.C(n_187),
.Y(n_244)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_212),
.Y(n_237)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_237),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_253),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_246),
.A2(n_248),
.B1(n_34),
.B2(n_29),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_210),
.B1(n_204),
.B2(n_184),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_250),
.B(n_28),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_191),
.B(n_192),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_206),
.C(n_209),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_254),
.C(n_257),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_252),
.A2(n_219),
.B1(n_234),
.B2(n_232),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_211),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_42),
.C(n_25),
.Y(n_254)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_217),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_225),
.C(n_226),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_259),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_241),
.B(n_220),
.Y(n_260)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_251),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_257),
.C(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_258),
.A2(n_234),
.B1(n_216),
.B2(n_29),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_263),
.A2(n_272),
.B1(n_274),
.B2(n_247),
.Y(n_278)
);

BUFx12_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_242),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_240),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_266),
.B(n_269),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_234),
.Y(n_267)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_275),
.B(n_14),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_255),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_272),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_252),
.A2(n_29),
.B1(n_34),
.B2(n_2),
.Y(n_272)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_11),
.C(n_16),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_9),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_252),
.A2(n_42),
.B1(n_29),
.B2(n_3),
.Y(n_274)
);

OAI321xp33_ASAP7_75t_L g275 ( 
.A1(n_252),
.A2(n_9),
.A3(n_16),
.B1(n_3),
.B2(n_4),
.C(n_6),
.Y(n_275)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_278),
.B(n_288),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_284),
.C(n_285),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_283),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_239),
.C(n_254),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_239),
.C(n_25),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_274),
.B(n_268),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_290),
.B(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_25),
.C(n_2),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_289),
.B(n_290),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_7),
.C(n_8),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_264),
.B1(n_276),
.B2(n_263),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_298),
.B1(n_300),
.B2(n_303),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_279),
.B(n_265),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_305),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_265),
.B1(n_1),
.B2(n_4),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_25),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_302),
.B(n_6),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_8),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_286),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_288),
.B(n_278),
.Y(n_305)
);

AO21x2_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_284),
.B(n_281),
.Y(n_306)
);

AOI21x1_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_313),
.B(n_304),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_295),
.B(n_292),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_307),
.A2(n_13),
.B(n_14),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_15),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_315),
.Y(n_321)
);

AOI211xp5_ASAP7_75t_L g313 ( 
.A1(n_293),
.A2(n_7),
.B(n_8),
.C(n_11),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_11),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_314),
.B(n_316),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_296),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_300),
.Y(n_316)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

AOI21x1_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_309),
.B(n_311),
.Y(n_318)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_318),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_296),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_319),
.B(n_320),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_306),
.B(n_13),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_324),
.B(n_15),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_15),
.B(n_16),
.Y(n_326)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_326),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_328),
.B(n_322),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_322),
.C(n_325),
.Y(n_332)
);

OAI21x1_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_327),
.B(n_329),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_333),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_331),
.Y(n_335)
);


endmodule