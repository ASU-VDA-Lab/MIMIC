module fake_aes_9286_n_569 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_569);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_569;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_73;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g71 ( .A(n_69), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_58), .Y(n_72) );
INVxp67_ASAP7_75t_SL g73 ( .A(n_50), .Y(n_73) );
CKINVDCx5p33_ASAP7_75t_R g74 ( .A(n_33), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_4), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_35), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_20), .Y(n_77) );
BUFx6f_ASAP7_75t_L g78 ( .A(n_22), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_60), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_30), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_41), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_64), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_19), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_62), .Y(n_84) );
INVxp67_ASAP7_75t_L g85 ( .A(n_52), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_18), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_66), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_36), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_24), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_17), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_0), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_8), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_43), .Y(n_93) );
INVxp33_ASAP7_75t_L g94 ( .A(n_25), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_68), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_13), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_21), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_13), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_32), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_3), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_15), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_29), .Y(n_102) );
BUFx5_ASAP7_75t_L g103 ( .A(n_2), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_34), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_6), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_46), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_55), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_38), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_17), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_45), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_15), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_48), .Y(n_112) );
NOR2xp67_ASAP7_75t_L g113 ( .A(n_11), .B(n_23), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_27), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_11), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_47), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_103), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_78), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_83), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_78), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_98), .B(n_0), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_98), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_103), .B(n_1), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_103), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_90), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_103), .Y(n_126) );
AND2x4_ASAP7_75t_L g127 ( .A(n_90), .B(n_1), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_94), .B(n_2), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_103), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_103), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_103), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_78), .Y(n_132) );
CKINVDCx8_ASAP7_75t_R g133 ( .A(n_114), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_78), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_103), .B(n_3), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_101), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_78), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_101), .B(n_4), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_107), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_107), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_72), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_75), .B(n_5), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
XOR2x2_ASAP7_75t_L g144 ( .A(n_91), .B(n_5), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_76), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_92), .B(n_6), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_79), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_81), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_86), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_96), .B(n_7), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_87), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_93), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_100), .B(n_7), .Y(n_155) );
NAND2xp33_ASAP7_75t_SL g156 ( .A(n_71), .B(n_8), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_128), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_146), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_146), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_128), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_127), .B(n_111), .Y(n_161) );
NAND2x1p5_ASAP7_75t_L g162 ( .A(n_135), .B(n_116), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_117), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_135), .B(n_106), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_117), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_127), .B(n_105), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_119), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_124), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_124), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_122), .B(n_85), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_125), .B(n_108), .Y(n_171) );
OR2x2_ASAP7_75t_L g172 ( .A(n_121), .B(n_115), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_118), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_126), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_141), .B(n_97), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_126), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_118), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_129), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_129), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_130), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_127), .B(n_113), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_141), .B(n_97), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_118), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_130), .Y(n_184) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_146), .B(n_102), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_118), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_131), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_131), .Y(n_188) );
NAND3xp33_ASAP7_75t_L g189 ( .A(n_123), .B(n_104), .C(n_110), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_147), .B(n_88), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_119), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_145), .Y(n_193) );
INVxp33_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_145), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_145), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_147), .B(n_88), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_133), .A2(n_109), .B1(n_71), .B2(n_89), .Y(n_198) );
AND2x6_ASAP7_75t_L g199 ( .A(n_151), .B(n_112), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_145), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_149), .B(n_108), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_145), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_145), .Y(n_203) );
INVx2_ASAP7_75t_SL g204 ( .A(n_119), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_151), .A2(n_106), .B1(n_74), .B2(n_77), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_120), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_120), .Y(n_207) );
NAND2xp33_ASAP7_75t_L g208 ( .A(n_149), .B(n_82), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_150), .B(n_82), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_140), .Y(n_210) );
NAND2x1p5_ASAP7_75t_L g211 ( .A(n_127), .B(n_80), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_143), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_164), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_190), .B(n_150), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_185), .A2(n_151), .B1(n_154), .B2(n_152), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_158), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_157), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_185), .B(n_151), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_175), .B(n_154), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_158), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_164), .B(n_182), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_171), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_185), .A2(n_156), .B1(n_155), .B2(n_138), .Y(n_224) );
INVx8_ASAP7_75t_L g225 ( .A(n_199), .Y(n_225) );
INVxp67_ASAP7_75t_SL g226 ( .A(n_162), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_212), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_182), .B(n_152), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_201), .B(n_138), .Y(n_229) );
NOR2xp67_ASAP7_75t_L g230 ( .A(n_189), .B(n_153), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_161), .A2(n_153), .B1(n_148), .B2(n_140), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_158), .B(n_143), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_212), .Y(n_233) );
BUFx2_ASAP7_75t_L g234 ( .A(n_171), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_201), .B(n_148), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_167), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_195), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_209), .B(n_142), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_158), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_167), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_195), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_192), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_157), .A2(n_89), .B1(n_144), .B2(n_74), .Y(n_243) );
OR2x6_ASAP7_75t_L g244 ( .A(n_211), .B(n_133), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_209), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_162), .Y(n_246) );
OAI22xp5_ASAP7_75t_SL g247 ( .A1(n_160), .A2(n_144), .B1(n_77), .B2(n_80), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_181), .B(n_136), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_192), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_172), .A2(n_136), .B(n_139), .C(n_143), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_162), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_159), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_181), .B(n_139), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_160), .B(n_139), .Y(n_254) );
OR2x2_ASAP7_75t_SL g255 ( .A(n_198), .B(n_9), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_197), .B(n_139), .Y(n_256) );
BUFx4f_ASAP7_75t_L g257 ( .A(n_211), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_211), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_205), .Y(n_259) );
OR2x2_ASAP7_75t_SL g260 ( .A(n_172), .B(n_9), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_181), .B(n_99), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_206), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_159), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_199), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_210), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_210), .Y(n_266) );
AND2x6_ASAP7_75t_SL g267 ( .A(n_181), .B(n_10), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_213), .A2(n_73), .B(n_132), .C(n_120), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_213), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_161), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_161), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_159), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_159), .B(n_137), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_226), .B(n_194), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_265), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_263), .Y(n_276) );
NOR2xp67_ASAP7_75t_L g277 ( .A(n_221), .B(n_191), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_262), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_218), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_247), .Y(n_280) );
INVx5_ASAP7_75t_L g281 ( .A(n_263), .Y(n_281) );
INVxp67_ASAP7_75t_L g282 ( .A(n_234), .Y(n_282) );
INVx4_ASAP7_75t_L g283 ( .A(n_263), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_263), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_262), .Y(n_285) );
INVx3_ASAP7_75t_SL g286 ( .A(n_244), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_266), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_221), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_257), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_220), .A2(n_189), .B(n_161), .C(n_166), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_269), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_240), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_219), .A2(n_199), .B1(n_191), .B2(n_166), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_223), .B(n_170), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_219), .A2(n_199), .B1(n_191), .B2(n_166), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_238), .B(n_166), .Y(n_296) );
AOI22xp33_ASAP7_75t_SL g297 ( .A1(n_257), .A2(n_199), .B1(n_208), .B2(n_191), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_221), .Y(n_298) );
BUFx8_ASAP7_75t_L g299 ( .A(n_246), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_239), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_218), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_229), .B(n_199), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_SL g303 ( .A1(n_268), .A2(n_204), .B(n_165), .C(n_163), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_240), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_233), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_216), .A2(n_199), .B1(n_204), .B2(n_163), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_251), .B(n_180), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_239), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_243), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_227), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_239), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_272), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_272), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_227), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_222), .B(n_165), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_233), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_258), .B(n_180), .Y(n_317) );
INVx2_ASAP7_75t_SL g318 ( .A(n_272), .Y(n_318) );
BUFx12f_ASAP7_75t_L g319 ( .A(n_267), .Y(n_319) );
OAI22xp33_ASAP7_75t_L g320 ( .A1(n_286), .A2(n_244), .B1(n_306), .B2(n_295), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_279), .A2(n_259), .B1(n_244), .B2(n_216), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_301), .A2(n_259), .B1(n_224), .B2(n_238), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_301), .A2(n_214), .B1(n_245), .B2(n_238), .Y(n_323) );
INVx4_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_299), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_274), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_274), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_299), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_276), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_290), .A2(n_228), .B(n_250), .C(n_256), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g331 ( .A1(n_286), .A2(n_225), .B1(n_271), .B2(n_255), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_275), .Y(n_332) );
OAI22xp33_ASAP7_75t_L g333 ( .A1(n_286), .A2(n_225), .B1(n_260), .B2(n_235), .Y(n_333) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_306), .A2(n_225), .B1(n_235), .B2(n_264), .Y(n_334) );
AOI222xp33_ASAP7_75t_L g335 ( .A1(n_319), .A2(n_294), .B1(n_282), .B2(n_309), .C1(n_299), .C2(n_229), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_307), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_296), .A2(n_268), .B(n_261), .C(n_220), .Y(n_337) );
OR2x6_ASAP7_75t_L g338 ( .A(n_289), .B(n_229), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_281), .B(n_233), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_295), .A2(n_270), .B1(n_230), .B2(n_248), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_281), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_289), .B(n_254), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_307), .B(n_248), .Y(n_343) );
NAND2x1p5_ASAP7_75t_L g344 ( .A(n_281), .B(n_217), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_302), .A2(n_248), .B1(n_253), .B2(n_215), .Y(n_345) );
AOI222xp33_ASAP7_75t_L g346 ( .A1(n_319), .A2(n_253), .B1(n_215), .B2(n_231), .C1(n_232), .C2(n_252), .Y(n_346) );
INVx6_ASAP7_75t_L g347 ( .A(n_281), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_276), .Y(n_348) );
BUFx12f_ASAP7_75t_L g349 ( .A(n_328), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_331), .A2(n_302), .B1(n_280), .B2(n_315), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_347), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_330), .A2(n_334), .B(n_303), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_333), .B(n_307), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_334), .A2(n_285), .B(n_278), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_332), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_348), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_329), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_326), .B(n_275), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_325), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_336), .B(n_287), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_327), .B(n_291), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_337), .A2(n_278), .B(n_285), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_331), .B(n_291), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_324), .Y(n_364) );
AO31x2_ASAP7_75t_L g365 ( .A1(n_324), .A2(n_287), .A3(n_132), .B(n_314), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_333), .A2(n_253), .B1(n_297), .B2(n_293), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_320), .A2(n_231), .B1(n_316), .B2(n_305), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_320), .A2(n_313), .B1(n_311), .B2(n_288), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_346), .A2(n_313), .B1(n_311), .B2(n_288), .Y(n_369) );
AOI222xp33_ASAP7_75t_L g370 ( .A1(n_323), .A2(n_312), .B1(n_308), .B2(n_298), .C1(n_300), .C2(n_317), .Y(n_370) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_340), .A2(n_310), .B(n_314), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_322), .B(n_298), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_335), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_321), .A2(n_288), .B1(n_313), .B2(n_311), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_355), .B(n_341), .Y(n_375) );
INVx4_ASAP7_75t_L g376 ( .A(n_349), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_373), .A2(n_340), .B1(n_345), .B2(n_343), .C(n_342), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_360), .Y(n_378) );
OAI31xp33_ASAP7_75t_L g379 ( .A1(n_353), .A2(n_344), .A3(n_341), .B(n_308), .Y(n_379) );
NAND3xp33_ASAP7_75t_L g380 ( .A(n_350), .B(n_339), .C(n_134), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_366), .A2(n_338), .B1(n_347), .B2(n_283), .Y(n_381) );
NAND3xp33_ASAP7_75t_L g382 ( .A(n_370), .B(n_137), .C(n_134), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_355), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_360), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_365), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_363), .B(n_338), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g387 ( .A(n_370), .B(n_137), .C(n_134), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_358), .B(n_338), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_356), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_364), .B(n_347), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g391 ( .A1(n_352), .A2(n_232), .B(n_277), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_363), .A2(n_312), .B1(n_283), .B2(n_273), .C(n_318), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_372), .B(n_344), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_372), .A2(n_283), .B1(n_273), .B2(n_318), .C(n_200), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_359), .B(n_281), .Y(n_395) );
AOI33xp33_ASAP7_75t_L g396 ( .A1(n_374), .A2(n_132), .A3(n_202), .B1(n_200), .B2(n_193), .B3(n_196), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_349), .B(n_361), .Y(n_397) );
AOI211xp5_ASAP7_75t_SL g398 ( .A1(n_367), .A2(n_277), .B(n_310), .C(n_203), .Y(n_398) );
AOI322xp5_ASAP7_75t_L g399 ( .A1(n_349), .A2(n_10), .A3(n_12), .B1(n_14), .B2(n_16), .C1(n_196), .C2(n_203), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_356), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_356), .Y(n_401) );
OAI211xp5_ASAP7_75t_L g402 ( .A1(n_369), .A2(n_193), .B(n_202), .C(n_137), .Y(n_402) );
AOI21x1_ASAP7_75t_L g403 ( .A1(n_367), .A2(n_241), .B(n_237), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_368), .A2(n_316), .B1(n_305), .B2(n_304), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_371), .A2(n_284), .B1(n_276), .B2(n_249), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_361), .B(n_276), .Y(n_406) );
AOI33xp33_ASAP7_75t_L g407 ( .A1(n_377), .A2(n_207), .A3(n_206), .B1(n_364), .B2(n_16), .B3(n_14), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_397), .B(n_364), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_378), .B(n_351), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_383), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_385), .B(n_371), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_388), .A2(n_362), .B1(n_371), .B2(n_354), .C(n_351), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_385), .B(n_371), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_389), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_384), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_375), .B(n_365), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_375), .B(n_365), .Y(n_417) );
NAND3xp33_ASAP7_75t_L g418 ( .A(n_399), .B(n_118), .C(n_134), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_389), .Y(n_419) );
OAI33xp33_ASAP7_75t_L g420 ( .A1(n_386), .A2(n_12), .A3(n_357), .B1(n_207), .B2(n_137), .B3(n_134), .Y(n_420) );
AO21x2_ASAP7_75t_L g421 ( .A1(n_382), .A2(n_357), .B(n_365), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_400), .B(n_365), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_380), .A2(n_351), .B1(n_357), .B2(n_284), .Y(n_423) );
NOR3xp33_ASAP7_75t_SL g424 ( .A(n_395), .B(n_365), .C(n_169), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_401), .B(n_118), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_401), .B(n_134), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_376), .Y(n_427) );
AOI211xp5_ASAP7_75t_L g428 ( .A1(n_387), .A2(n_284), .B(n_276), .C(n_304), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_403), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_393), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_393), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_403), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_386), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_380), .A2(n_292), .B1(n_305), .B2(n_316), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_390), .B(n_316), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_406), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_390), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_399), .B(n_284), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_404), .Y(n_439) );
NOR2xp67_ASAP7_75t_L g440 ( .A(n_405), .B(n_26), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_391), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_379), .B(n_316), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_376), .Y(n_444) );
AOI33xp33_ASAP7_75t_L g445 ( .A1(n_381), .A2(n_184), .A3(n_179), .B1(n_168), .B2(n_188), .B3(n_237), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_376), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_379), .B(n_305), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_398), .B(n_305), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_415), .B(n_402), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_418), .A2(n_392), .B1(n_394), .B2(n_284), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_437), .B(n_28), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_416), .B(n_31), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_410), .Y(n_453) );
NAND2x1_ASAP7_75t_L g454 ( .A(n_444), .B(n_233), .Y(n_454) );
NAND4xp25_ASAP7_75t_L g455 ( .A(n_418), .B(n_249), .C(n_236), .D(n_252), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_416), .B(n_37), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_410), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_419), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_424), .B(n_186), .C(n_177), .Y(n_459) );
NAND4xp25_ASAP7_75t_L g460 ( .A(n_408), .B(n_236), .C(n_217), .D(n_241), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_430), .B(n_242), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_431), .B(n_242), .Y(n_462) );
NAND4xp25_ASAP7_75t_L g463 ( .A(n_407), .B(n_188), .C(n_179), .D(n_187), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_417), .B(n_39), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_444), .B(n_40), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_444), .B(n_446), .Y(n_466) );
NOR3xp33_ASAP7_75t_SL g467 ( .A(n_420), .B(n_42), .C(n_44), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_431), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_436), .B(n_242), .Y(n_469) );
OAI311xp33_ASAP7_75t_L g470 ( .A1(n_438), .A2(n_49), .A3(n_51), .B1(n_53), .C1(n_54), .Y(n_470) );
OAI211xp5_ASAP7_75t_L g471 ( .A1(n_427), .A2(n_240), .B(n_173), .C(n_186), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_436), .B(n_56), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_417), .B(n_57), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_409), .B(n_59), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_433), .B(n_61), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_433), .B(n_63), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_414), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_433), .B(n_65), .Y(n_478) );
NAND4xp25_ASAP7_75t_L g479 ( .A(n_446), .B(n_187), .C(n_178), .D(n_176), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_419), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_433), .B(n_67), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g482 ( .A1(n_446), .A2(n_177), .B1(n_173), .B2(n_183), .C(n_186), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_435), .B(n_70), .Y(n_483) );
AOI32xp33_ASAP7_75t_L g484 ( .A1(n_428), .A2(n_174), .A3(n_176), .B1(n_178), .B2(n_177), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_422), .B(n_173), .Y(n_485) );
INVx4_ASAP7_75t_L g486 ( .A(n_442), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_422), .Y(n_487) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_441), .A2(n_443), .B1(n_413), .B2(n_411), .C(n_412), .Y(n_488) );
AND2x4_ASAP7_75t_SL g489 ( .A(n_447), .B(n_183), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_468), .B(n_413), .Y(n_490) );
OAI31xp33_ASAP7_75t_L g491 ( .A1(n_455), .A2(n_443), .A3(n_447), .B(n_448), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_484), .B(n_428), .Y(n_492) );
INVxp67_ASAP7_75t_SL g493 ( .A(n_466), .Y(n_493) );
AO211x2_ASAP7_75t_L g494 ( .A1(n_460), .A2(n_432), .B(n_440), .C(n_445), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_487), .B(n_411), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_466), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_487), .B(n_411), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_477), .B(n_421), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_453), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_449), .Y(n_500) );
AO211x2_ASAP7_75t_L g501 ( .A1(n_459), .A2(n_432), .B(n_440), .C(n_423), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_486), .B(n_439), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_452), .B(n_426), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_457), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_457), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_486), .B(n_448), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_486), .B(n_439), .Y(n_507) );
NAND3xp33_ASAP7_75t_SL g508 ( .A(n_467), .B(n_434), .C(n_426), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_458), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_474), .B(n_425), .C(n_429), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_473), .B(n_183), .Y(n_511) );
XNOR2xp5_ASAP7_75t_L g512 ( .A(n_473), .B(n_183), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_454), .Y(n_513) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_472), .B(n_183), .C(n_186), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_489), .B(n_480), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_480), .B(n_485), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_488), .B(n_465), .C(n_463), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_456), .A2(n_464), .B1(n_479), .B2(n_465), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_450), .A2(n_489), .B1(n_451), .B2(n_483), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_469), .B(n_461), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_462), .B(n_475), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_517), .A2(n_467), .B(n_450), .C(n_471), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_500), .B(n_481), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_515), .B(n_478), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_496), .B(n_476), .Y(n_525) );
INVxp67_ASAP7_75t_SL g526 ( .A(n_493), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_518), .A2(n_470), .B1(n_482), .B2(n_492), .Y(n_527) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_512), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_492), .A2(n_501), .B(n_494), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_506), .Y(n_530) );
XNOR2xp5_ASAP7_75t_L g531 ( .A(n_494), .B(n_519), .Y(n_531) );
AOI31xp33_ASAP7_75t_SL g532 ( .A1(n_495), .A2(n_497), .A3(n_507), .B(n_502), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_490), .B(n_520), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_504), .Y(n_534) );
NAND2xp33_ASAP7_75t_SL g535 ( .A(n_515), .B(n_503), .Y(n_535) );
XNOR2x1_ASAP7_75t_L g536 ( .A(n_501), .B(n_516), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_510), .A2(n_508), .B1(n_521), .B2(n_515), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g538 ( .A1(n_498), .A2(n_499), .B1(n_505), .B2(n_509), .C(n_511), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_514), .A2(n_492), .B(n_501), .Y(n_539) );
XNOR2xp5_ASAP7_75t_L g540 ( .A(n_500), .B(n_359), .Y(n_540) );
XNOR2x1_ASAP7_75t_L g541 ( .A(n_500), .B(n_144), .Y(n_541) );
OAI221xp5_ASAP7_75t_L g542 ( .A1(n_517), .A2(n_373), .B1(n_491), .B2(n_519), .C(n_518), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_513), .B(n_515), .Y(n_543) );
NOR3xp33_ASAP7_75t_L g544 ( .A(n_517), .B(n_333), .C(n_373), .Y(n_544) );
AOI31xp33_ASAP7_75t_L g545 ( .A1(n_519), .A2(n_492), .A3(n_506), .B(n_427), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_515), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_526), .Y(n_547) );
INVxp67_ASAP7_75t_L g548 ( .A(n_540), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g549 ( .A(n_529), .B(n_539), .C(n_531), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_545), .A2(n_531), .B1(n_528), .B2(n_536), .Y(n_550) );
AOI211x1_ASAP7_75t_SL g551 ( .A1(n_522), .A2(n_543), .B(n_536), .C(n_524), .Y(n_551) );
AOI211xp5_ASAP7_75t_L g552 ( .A1(n_542), .A2(n_532), .B(n_544), .C(n_522), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_533), .B(n_538), .Y(n_553) );
OAI221xp5_ASAP7_75t_L g554 ( .A1(n_550), .A2(n_527), .B1(n_537), .B2(n_544), .C(n_530), .Y(n_554) );
AO22x2_ASAP7_75t_L g555 ( .A1(n_549), .A2(n_541), .B1(n_543), .B2(n_546), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_SL g556 ( .A1(n_552), .A2(n_525), .B(n_523), .C(n_534), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_547), .Y(n_557) );
XNOR2x2_ASAP7_75t_L g558 ( .A(n_551), .B(n_524), .Y(n_558) );
AOI211xp5_ASAP7_75t_L g559 ( .A1(n_554), .A2(n_548), .B(n_553), .C(n_535), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_557), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_555), .Y(n_561) );
AO22x2_ASAP7_75t_L g562 ( .A1(n_561), .A2(n_555), .B1(n_558), .B2(n_556), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_560), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_563), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_562), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_564), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_566), .Y(n_567) );
BUFx2_ASAP7_75t_L g568 ( .A(n_567), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_568), .A2(n_565), .B(n_559), .Y(n_569) );
endmodule