module fake_ibex_481_n_4501 (n_151, n_85, n_599, n_778, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_785, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_810, n_768, n_338, n_173, n_696, n_796, n_797, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_799, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_217, n_324, n_391, n_537, n_728, n_78, n_805, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_232, n_380, n_749, n_281, n_559, n_425, n_4501);

input n_151;
input n_85;
input n_599;
input n_778;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_785;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_810;
input n_768;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4501;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4449;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_845;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_4343;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4353;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4421;
wire n_4179;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_4360;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_4378;
wire n_850;
wire n_4169;
wire n_3175;
wire n_3729;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_4477;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_4418;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_875;
wire n_1307;
wire n_4431;
wire n_1327;
wire n_2644;
wire n_4445;
wire n_876;
wire n_3211;
wire n_3479;
wire n_1840;
wire n_2837;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_4470;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3896;
wire n_3753;
wire n_2192;
wire n_4423;
wire n_1766;
wire n_3566;
wire n_3184;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_824;
wire n_4304;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_4382;
wire n_2860;
wire n_2448;
wire n_4002;
wire n_3631;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_4450;
wire n_3969;
wire n_4467;
wire n_1081;
wire n_4437;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_4447;
wire n_4491;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3884;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_4389;
wire n_2846;
wire n_2685;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_4312;
wire n_917;
wire n_2249;
wire n_3022;
wire n_2362;
wire n_968;
wire n_2413;
wire n_3148;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_3973;
wire n_1313;
wire n_4214;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_4430;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_4433;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_4428;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3097;
wire n_3030;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_4479;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_4422;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_4481;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_971;
wire n_1326;
wire n_4444;
wire n_1350;
wire n_3627;
wire n_906;
wire n_4499;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_3199;
wire n_1616;
wire n_2723;
wire n_3808;
wire n_4455;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_4480;
wire n_1613;
wire n_820;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_4290;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_4252;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_4476;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_3317;
wire n_3887;
wire n_3800;
wire n_3963;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4126;
wire n_3583;
wire n_2019;
wire n_4103;
wire n_1407;
wire n_3282;
wire n_4435;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_819;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4156;
wire n_1964;
wire n_4411;
wire n_4408;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_4489;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_4419;
wire n_1583;
wire n_3520;
wire n_4404;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3733;
wire n_3626;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_4494;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4122;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_4374;
wire n_1140;
wire n_1985;
wire n_4375;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_4403;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_2573;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2423;
wire n_4230;
wire n_859;
wire n_3849;
wire n_965;
wire n_1109;
wire n_4402;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4469;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_4460;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_4485;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_1236;
wire n_3364;
wire n_4384;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4323;
wire n_4407;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_907;
wire n_1990;
wire n_3680;
wire n_4462;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_4490;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_3503;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1566;
wire n_1464;
wire n_4362;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_3331;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2590;
wire n_3119;
wire n_4414;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_4409;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_4443;
wire n_1682;
wire n_4151;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2991;
wire n_2234;
wire n_847;
wire n_2699;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_4424;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_4415;
wire n_1345;
wire n_4215;
wire n_4456;
wire n_4315;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_4492;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_3470;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_4500;
wire n_1395;
wire n_998;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_4427;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_882;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_3829;
wire n_1864;
wire n_943;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_3460;
wire n_2905;
wire n_3978;
wire n_3954;
wire n_2570;
wire n_4051;
wire n_4321;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4416;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_817;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_863;
wire n_2185;
wire n_4141;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_4117;
wire n_3999;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_4496;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4195;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1185;
wire n_1683;
wire n_4256;
wire n_3575;
wire n_4454;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_4278;
wire n_874;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_4458;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_3158;
wire n_1535;
wire n_2985;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_4276;
wire n_831;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_2875;
wire n_3284;
wire n_2524;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1941;
wire n_1707;
wire n_3927;
wire n_3902;
wire n_2422;
wire n_4185;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_920;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_4441;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_961;
wire n_1331;
wire n_991;
wire n_1223;
wire n_2127;
wire n_3891;
wire n_3735;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3228;
wire n_3028;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_4497;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_4483;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4488;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4142;
wire n_4118;
wire n_2138;
wire n_1380;
wire n_4302;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1458;
wire n_1694;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_4066;
wire n_3990;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3269;
wire n_3029;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4123;
wire n_3154;
wire n_4000;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2683;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3696;
wire n_3113;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_4007;
wire n_3960;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_4286;
wire n_4429;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_4438;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_4498;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1348;
wire n_838;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_3930;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_4149;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_4319;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_3773;
wire n_2528;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_4466;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_4417;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1946;
wire n_1726;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2984;
wire n_3162;
wire n_2732;
wire n_4436;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_3333;
wire n_3096;
wire n_839;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_4434;
wire n_2737;
wire n_2251;
wire n_2012;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2447;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_4367;
wire n_950;
wire n_3139;
wire n_2700;
wire n_1222;
wire n_4282;
wire n_1630;
wire n_3408;
wire n_4475;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3647;
wire n_3623;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_4410;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_3229;
wire n_2225;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_4440;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2576;
wire n_2675;
wire n_2417;
wire n_2348;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4111;
wire n_4162;
wire n_4200;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_4439;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_4058;
wire n_4487;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4148;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_2803;
wire n_2816;
wire n_2433;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4017;
wire n_1542;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1547;
wire n_3497;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_3561;
wire n_2313;
wire n_2381;
wire n_3586;
wire n_956;
wire n_4125;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_2574;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_2911;
wire n_1623;
wire n_861;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_4453;
wire n_1098;
wire n_4474;
wire n_1366;
wire n_1518;
wire n_4350;
wire n_4380;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_4281;
wire n_4345;
wire n_4478;
wire n_2411;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_4473;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_4464;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2929;
wire n_2701;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_854;
wire n_4432;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_4405;
wire n_3118;
wire n_1369;
wire n_1912;
wire n_1297;
wire n_3143;
wire n_3543;
wire n_1734;
wire n_3655;
wire n_3791;
wire n_3742;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4461;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_914;
wire n_3992;
wire n_4147;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_4471;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3547;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_4386;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_4482;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_4406;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_4493;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1488;
wire n_849;
wire n_1193;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3380;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1904;
wire n_1262;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_4412;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3483;
wire n_3160;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3124;
wire n_999;
wire n_2634;
wire n_2982;
wire n_3286;
wire n_1092;
wire n_4038;
wire n_4472;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_1230;
wire n_4459;
wire n_1027;
wire n_1516;
wire n_3893;
wire n_4484;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_3938;
wire n_4354;
wire n_924;
wire n_4448;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_4401;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_4413;
wire n_1757;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2560;
wire n_2302;
wire n_3056;
wire n_2453;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3189;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_2066;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_4275;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_3283;
wire n_4468;
wire n_1736;
wire n_4442;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_3613;
wire n_1383;
wire n_990;
wire n_4108;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2749;
wire n_888;
wire n_2378;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2738;
wire n_2324;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_4486;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_4327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_4465;
wire n_1355;
wire n_3691;
wire n_4452;
wire n_2544;
wire n_856;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_4183;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_4425;
wire n_3980;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_2970;
wire n_1393;
wire n_2497;
wire n_984;
wire n_1655;
wire n_3494;
wire n_3040;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_642),
.Y(n_816)
);

BUFx10_ASAP7_75t_L g817 ( 
.A(n_721),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_208),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_191),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_700),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_589),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_559),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_720),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_454),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_510),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_690),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_586),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_667),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_380),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_416),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_401),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_704),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_43),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_728),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_708),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_679),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_469),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_650),
.Y(n_838)
);

BUFx10_ASAP7_75t_L g839 ( 
.A(n_247),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_654),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_599),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_306),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_333),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_253),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_802),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_139),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_468),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_493),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_81),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_613),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_614),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_165),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_650),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_752),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_749),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_52),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_686),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_730),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_310),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_669),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_748),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_651),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_778),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_6),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_392),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_529),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_662),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_733),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_736),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_28),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_331),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_537),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_715),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_528),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_46),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_358),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_527),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_788),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_646),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_16),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_616),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_352),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_339),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_603),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_562),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_737),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_161),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_376),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_804),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_786),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_305),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_580),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_98),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_103),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_67),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_717),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_741),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_490),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_351),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_161),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_611),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_735),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_363),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_101),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_380),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_747),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_467),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_620),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_553),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_776),
.Y(n_910)
);

CKINVDCx20_ASAP7_75t_R g911 ( 
.A(n_725),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_764),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_680),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_501),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_132),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_75),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_285),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_121),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_149),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_357),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_543),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_12),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_444),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_803),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_610),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_435),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_748),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_437),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_534),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_556),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_178),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_664),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_719),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_469),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_128),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_31),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_272),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_110),
.Y(n_938)
);

BUFx10_ASAP7_75t_L g939 ( 
.A(n_570),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_646),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_544),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_254),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_815),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_224),
.Y(n_944)
);

CKINVDCx16_ASAP7_75t_R g945 ( 
.A(n_698),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_289),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_69),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_309),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_271),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_21),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_680),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_257),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_172),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_562),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_557),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_701),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_24),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_258),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_258),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_740),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_505),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_276),
.Y(n_962)
);

INVx4_ASAP7_75t_R g963 ( 
.A(n_738),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_294),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_509),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_491),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_811),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_223),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_397),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_421),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_713),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_136),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_271),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_278),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_478),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_470),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_105),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_51),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_81),
.Y(n_979)
);

CKINVDCx14_ASAP7_75t_R g980 ( 
.A(n_421),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_44),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_737),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_198),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_762),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_447),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_535),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_457),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_577),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_653),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_529),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_563),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_653),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_694),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_32),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_743),
.Y(n_995)
);

CKINVDCx16_ASAP7_75t_R g996 ( 
.A(n_124),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_245),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_514),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_703),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_579),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_195),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_19),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_586),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_39),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_8),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_363),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_229),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_347),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_725),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_35),
.Y(n_1010)
);

CKINVDCx14_ASAP7_75t_R g1011 ( 
.A(n_579),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_225),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_643),
.Y(n_1013)
);

CKINVDCx11_ASAP7_75t_R g1014 ( 
.A(n_798),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_721),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_440),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_641),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_408),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_591),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_158),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_381),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_688),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_116),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_449),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_691),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_197),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_666),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_807),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_541),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_365),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_109),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_132),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_808),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_405),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_427),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_407),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_220),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_101),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_316),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_711),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_602),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_316),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_256),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_326),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_681),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_403),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_768),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_108),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_536),
.Y(n_1049)
);

INVxp33_ASAP7_75t_L g1050 ( 
.A(n_681),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_457),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_568),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_657),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_131),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_236),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_279),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_458),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_52),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_777),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_542),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_402),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_538),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_257),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_154),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_746),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_547),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_720),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_706),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_234),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_750),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_727),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_238),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_454),
.Y(n_1073)
);

BUFx10_ASAP7_75t_L g1074 ( 
.A(n_729),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_3),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_173),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_709),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_345),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_188),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_734),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_396),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_565),
.Y(n_1082)
);

BUFx5_ASAP7_75t_L g1083 ( 
.A(n_672),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_424),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_793),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_691),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_83),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_633),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_105),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_301),
.Y(n_1090)
);

CKINVDCx16_ASAP7_75t_R g1091 ( 
.A(n_371),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_665),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_250),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_714),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_494),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_104),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_248),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_83),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_387),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_410),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_515),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_710),
.Y(n_1102)
);

BUFx10_ASAP7_75t_L g1103 ( 
.A(n_17),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_500),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_84),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_558),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_305),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_372),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_85),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_278),
.Y(n_1110)
);

BUFx10_ASAP7_75t_L g1111 ( 
.A(n_629),
.Y(n_1111)
);

CKINVDCx14_ASAP7_75t_R g1112 ( 
.A(n_118),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_207),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_215),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_706),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_289),
.Y(n_1116)
);

BUFx10_ASAP7_75t_L g1117 ( 
.A(n_571),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_456),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_747),
.Y(n_1119)
);

BUFx10_ASAP7_75t_L g1120 ( 
.A(n_455),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_133),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_40),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_533),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_712),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_502),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_210),
.Y(n_1126)
);

CKINVDCx16_ASAP7_75t_R g1127 ( 
.A(n_741),
.Y(n_1127)
);

BUFx10_ASAP7_75t_L g1128 ( 
.A(n_814),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_361),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_393),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_722),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_754),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_673),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_731),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_765),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_118),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_125),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_48),
.Y(n_1138)
);

CKINVDCx14_ASAP7_75t_R g1139 ( 
.A(n_489),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_125),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_534),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_809),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_284),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_466),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_476),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_183),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_286),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_447),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_73),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_724),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_698),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_607),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_114),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_220),
.Y(n_1154)
);

INVxp67_ASAP7_75t_SL g1155 ( 
.A(n_61),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_6),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_612),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_770),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_39),
.Y(n_1159)
);

CKINVDCx20_ASAP7_75t_R g1160 ( 
.A(n_424),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_119),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_136),
.Y(n_1162)
);

BUFx3_ASAP7_75t_L g1163 ( 
.A(n_282),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_746),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_144),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_717),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_335),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_219),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_313),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_708),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_488),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_210),
.Y(n_1172)
);

CKINVDCx14_ASAP7_75t_R g1173 ( 
.A(n_563),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_328),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_658),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_407),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_742),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_226),
.Y(n_1178)
);

CKINVDCx16_ASAP7_75t_R g1179 ( 
.A(n_71),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_508),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_2),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_234),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_568),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_429),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_644),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_805),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_616),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_648),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_392),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_726),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_86),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_190),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_89),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_640),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_569),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_353),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_609),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_134),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_584),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_701),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_222),
.Y(n_1201)
);

BUFx10_ASAP7_75t_L g1202 ( 
.A(n_154),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_435),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_311),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_775),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_718),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_707),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_578),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_810),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_473),
.Y(n_1210)
);

BUFx10_ASAP7_75t_L g1211 ( 
.A(n_394),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_261),
.Y(n_1212)
);

BUFx10_ASAP7_75t_L g1213 ( 
.A(n_611),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_139),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_527),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_335),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_742),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_25),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_281),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_723),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_152),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_144),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_241),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_245),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_207),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_302),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_702),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_697),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_95),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_812),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_618),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_331),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_193),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_397),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_772),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_313),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_170),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_657),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_151),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_656),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_705),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_745),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_231),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_445),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_626),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_82),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_17),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_249),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_255),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_669),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_604),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_281),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_354),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_34),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_196),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_673),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_111),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_337),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_405),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_704),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_56),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_464),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_495),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_423),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_743),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_99),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_322),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_744),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_384),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_165),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_716),
.Y(n_1272)
);

CKINVDCx16_ASAP7_75t_R g1273 ( 
.A(n_476),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_152),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_344),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_108),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_702),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_490),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_759),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_440),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_739),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_138),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_175),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_473),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_630),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_127),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_332),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_224),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_662),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_254),
.Y(n_1290)
);

BUFx5_ASAP7_75t_L g1291 ( 
.A(n_714),
.Y(n_1291)
);

BUFx8_ASAP7_75t_SL g1292 ( 
.A(n_87),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_732),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_67),
.Y(n_1294)
);

BUFx2_ASAP7_75t_SL g1295 ( 
.A(n_11),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_536),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_658),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_282),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_121),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_93),
.Y(n_1300)
);

INVx1_ASAP7_75t_SL g1301 ( 
.A(n_349),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_138),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_437),
.Y(n_1303)
);

INVxp33_ASAP7_75t_SL g1304 ( 
.A(n_295),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_467),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_8),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_622),
.Y(n_1307)
);

BUFx5_ASAP7_75t_L g1308 ( 
.A(n_48),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_730),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_607),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_609),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_415),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_141),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_205),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_500),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_732),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_574),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_250),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_361),
.Y(n_1319)
);

INVx5_ASAP7_75t_L g1320 ( 
.A(n_1142),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1142),
.B(n_0),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_958),
.Y(n_1322)
);

CKINVDCx6p67_ASAP7_75t_R g1323 ( 
.A(n_1014),
.Y(n_1323)
);

AND2x2_ASAP7_75t_SL g1324 ( 
.A(n_889),
.B(n_0),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_830),
.B(n_2),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1142),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_861),
.Y(n_1327)
);

NAND2xp33_ASAP7_75t_L g1328 ( 
.A(n_1083),
.B(n_751),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_901),
.B(n_3),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_861),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_861),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_SL g1332 ( 
.A(n_845),
.B(n_801),
.Y(n_1332)
);

INVx4_ASAP7_75t_L g1333 ( 
.A(n_1128),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_943),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_827),
.B(n_1),
.Y(n_1335)
);

BUFx8_ASAP7_75t_SL g1336 ( 
.A(n_1292),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_943),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_943),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_943),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1128),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1083),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_868),
.Y(n_1342)
);

INVx5_ASAP7_75t_L g1343 ( 
.A(n_1128),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1056),
.Y(n_1344)
);

BUFx8_ASAP7_75t_SL g1345 ( 
.A(n_1292),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_931),
.B(n_5),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1083),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_868),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1079),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1158),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1050),
.B(n_1146),
.Y(n_1351)
);

BUFx8_ASAP7_75t_L g1352 ( 
.A(n_1159),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1158),
.B(n_4),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1226),
.B(n_5),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_868),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1083),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1050),
.B(n_4),
.Y(n_1357)
);

INVx5_ASAP7_75t_L g1358 ( 
.A(n_868),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_877),
.Y(n_1359)
);

INVx5_ASAP7_75t_L g1360 ( 
.A(n_877),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1083),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_877),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_877),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1083),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_827),
.B(n_7),
.Y(n_1365)
);

INVx5_ASAP7_75t_L g1366 ( 
.A(n_893),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1083),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_843),
.B(n_9),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_945),
.B(n_7),
.Y(n_1369)
);

INVx4_ASAP7_75t_L g1370 ( 
.A(n_912),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1014),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_843),
.B(n_10),
.Y(n_1372)
);

NOR2x1_ASAP7_75t_L g1373 ( 
.A(n_1009),
.B(n_753),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_924),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_893),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_980),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1009),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_921),
.B(n_9),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_893),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_817),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1291),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_921),
.B(n_10),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_996),
.B(n_11),
.Y(n_1383)
);

INVx5_ASAP7_75t_L g1384 ( 
.A(n_893),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1091),
.B(n_12),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1021),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1021),
.B(n_14),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_SL g1388 ( 
.A(n_984),
.B(n_813),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_959),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_959),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1043),
.B(n_14),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1127),
.B(n_13),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1043),
.B(n_13),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1011),
.Y(n_1394)
);

BUFx12f_ASAP7_75t_L g1395 ( 
.A(n_817),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_959),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_967),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1179),
.B(n_1273),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_SL g1399 ( 
.A(n_1033),
.B(n_1047),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1112),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1219),
.B(n_16),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_854),
.B(n_15),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1219),
.B(n_18),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1291),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_959),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1229),
.B(n_15),
.Y(n_1406)
);

INVx5_ASAP7_75t_L g1407 ( 
.A(n_1002),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1291),
.Y(n_1408)
);

INVx4_ASAP7_75t_L g1409 ( 
.A(n_1059),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1229),
.B(n_19),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1291),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1306),
.Y(n_1412)
);

BUFx8_ASAP7_75t_L g1413 ( 
.A(n_1291),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1306),
.B(n_18),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_865),
.B(n_21),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1291),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1078),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1087),
.B(n_22),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1139),
.B(n_20),
.Y(n_1419)
);

INVx5_ASAP7_75t_L g1420 ( 
.A(n_1002),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1002),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1002),
.Y(n_1422)
);

BUFx12f_ASAP7_75t_L g1423 ( 
.A(n_817),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1078),
.B(n_20),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1173),
.B(n_22),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1102),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1080),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_856),
.B(n_24),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1291),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1080),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_839),
.B(n_23),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1131),
.B(n_23),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_839),
.B(n_25),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_839),
.B(n_26),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_939),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1308),
.Y(n_1436)
);

BUFx12f_ASAP7_75t_L g1437 ( 
.A(n_939),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_878),
.B(n_26),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_939),
.B(n_27),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1308),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1074),
.B(n_1103),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1074),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_856),
.B(n_28),
.Y(n_1443)
);

INVx5_ASAP7_75t_L g1444 ( 
.A(n_1102),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1308),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1351),
.A2(n_1323),
.B1(n_1344),
.B2(n_1322),
.Y(n_1446)
);

BUFx10_ASAP7_75t_L g1447 ( 
.A(n_1371),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1335),
.Y(n_1448)
);

OAI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1428),
.A2(n_1304),
.B1(n_860),
.B2(n_862),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1398),
.A2(n_1304),
.B1(n_860),
.B2(n_862),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1335),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1394),
.B(n_1400),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1349),
.B(n_1074),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1333),
.B(n_890),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1357),
.A2(n_1088),
.B1(n_1314),
.B2(n_859),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1376),
.B(n_1333),
.Y(n_1456)
);

BUFx10_ASAP7_75t_L g1457 ( 
.A(n_1365),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1365),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1324),
.A2(n_1088),
.B1(n_1314),
.B2(n_859),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1325),
.A2(n_1318),
.B1(n_1316),
.B2(n_844),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1343),
.B(n_1442),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1441),
.A2(n_1316),
.B1(n_1318),
.B2(n_967),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1380),
.A2(n_1442),
.B1(n_1346),
.B2(n_1329),
.Y(n_1463)
);

OAI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1354),
.A2(n_844),
.B1(n_846),
.B2(n_842),
.Y(n_1464)
);

OAI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1443),
.A2(n_846),
.B1(n_871),
.B2(n_842),
.Y(n_1465)
);

OAI22xp33_ASAP7_75t_SL g1466 ( 
.A1(n_1415),
.A2(n_818),
.B1(n_821),
.B2(n_816),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1340),
.B(n_1103),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1377),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1395),
.A2(n_1309),
.B1(n_873),
.B2(n_883),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1423),
.A2(n_1437),
.B1(n_1435),
.B2(n_1418),
.Y(n_1470)
);

AO22x2_ASAP7_75t_L g1471 ( 
.A1(n_1369),
.A2(n_1295),
.B1(n_1155),
.B2(n_850),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1343),
.B(n_1103),
.Y(n_1472)
);

OA22x2_ASAP7_75t_L g1473 ( 
.A1(n_1397),
.A2(n_824),
.B1(n_894),
.B2(n_834),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1368),
.A2(n_873),
.B1(n_883),
.B2(n_871),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1343),
.B(n_1111),
.Y(n_1475)
);

AO22x2_ASAP7_75t_L g1476 ( 
.A1(n_1383),
.A2(n_923),
.B1(n_929),
.B2(n_848),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1378),
.Y(n_1477)
);

AO22x2_ASAP7_75t_L g1478 ( 
.A1(n_1385),
.A2(n_1064),
.B1(n_1066),
.B2(n_982),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1413),
.Y(n_1479)
);

AOI22x1_ASAP7_75t_L g1480 ( 
.A1(n_1347),
.A2(n_1132),
.B1(n_1028),
.B2(n_1070),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1372),
.A2(n_1309),
.B1(n_911),
.B2(n_913),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1330),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1330),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1327),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1378),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1370),
.B(n_1305),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1413),
.Y(n_1487)
);

OA22x2_ASAP7_75t_L g1488 ( 
.A1(n_1386),
.A2(n_825),
.B1(n_867),
.B2(n_852),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1382),
.Y(n_1489)
);

AO22x2_ASAP7_75t_L g1490 ( 
.A1(n_1392),
.A2(n_1075),
.B1(n_1077),
.B2(n_1067),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1412),
.A2(n_911),
.B1(n_913),
.B2(n_887),
.Y(n_1491)
);

AO22x2_ASAP7_75t_L g1492 ( 
.A1(n_1382),
.A2(n_1161),
.B1(n_1201),
.B2(n_1096),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1387),
.A2(n_927),
.B1(n_957),
.B2(n_887),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1391),
.A2(n_957),
.B1(n_983),
.B2(n_927),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1336),
.A2(n_993),
.B1(n_1030),
.B2(n_983),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1327),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1393),
.Y(n_1497)
);

NOR2x1p5_ASAP7_75t_L g1498 ( 
.A(n_1345),
.B(n_1131),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1393),
.A2(n_826),
.B1(n_829),
.B2(n_822),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1331),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1401),
.A2(n_1030),
.B1(n_1041),
.B2(n_993),
.Y(n_1501)
);

INVxp67_ASAP7_75t_SL g1502 ( 
.A(n_1419),
.Y(n_1502)
);

OR2x6_ASAP7_75t_L g1503 ( 
.A(n_1431),
.B(n_1433),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1406),
.A2(n_833),
.B1(n_835),
.B2(n_831),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_R g1505 ( 
.A(n_1352),
.B(n_1085),
.Y(n_1505)
);

AO22x2_ASAP7_75t_L g1506 ( 
.A1(n_1406),
.A2(n_1228),
.B1(n_1244),
.B2(n_1207),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1358),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1358),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1350),
.B(n_1163),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1414),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1425),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1414),
.A2(n_841),
.B1(n_847),
.B2(n_838),
.Y(n_1512)
);

AO22x2_ASAP7_75t_L g1513 ( 
.A1(n_1424),
.A2(n_1301),
.B1(n_1310),
.B2(n_1300),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1358),
.Y(n_1514)
);

INVx8_ASAP7_75t_L g1515 ( 
.A(n_1424),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1370),
.Y(n_1516)
);

AO22x2_ASAP7_75t_L g1517 ( 
.A1(n_1432),
.A2(n_1319),
.B1(n_1313),
.B2(n_1315),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1432),
.A2(n_851),
.B1(n_855),
.B2(n_849),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1326),
.B(n_1111),
.Y(n_1519)
);

AND2x2_ASAP7_75t_SL g1520 ( 
.A(n_1434),
.B(n_836),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1360),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1360),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1360),
.Y(n_1523)
);

INVx1_ASAP7_75t_SL g1524 ( 
.A(n_1439),
.Y(n_1524)
);

OAI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1403),
.A2(n_870),
.B1(n_872),
.B2(n_866),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1366),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1326),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1410),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1417),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1374),
.B(n_1111),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1374),
.B(n_1117),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1366),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1409),
.B(n_1117),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1320),
.Y(n_1534)
);

AO22x2_ASAP7_75t_L g1535 ( 
.A1(n_1427),
.A2(n_1311),
.B1(n_1317),
.B2(n_1298),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1366),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1430),
.A2(n_1084),
.B1(n_1119),
.B2(n_1041),
.Y(n_1537)
);

OAI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1320),
.A2(n_1119),
.B1(n_1160),
.B2(n_1084),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1353),
.A2(n_875),
.B1(n_876),
.B2(n_874),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1409),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1320),
.A2(n_880),
.B1(n_881),
.B2(n_879),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1399),
.B(n_910),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1356),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1341),
.B(n_1117),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_SL g1545 ( 
.A1(n_1332),
.A2(n_884),
.B1(n_885),
.B2(n_882),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1341),
.B(n_1120),
.Y(n_1546)
);

OAI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1388),
.A2(n_1188),
.B1(n_1196),
.B2(n_1160),
.Y(n_1547)
);

OAI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1321),
.A2(n_888),
.B1(n_891),
.B2(n_886),
.Y(n_1548)
);

AND2x2_ASAP7_75t_SL g1549 ( 
.A(n_1328),
.B(n_836),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1381),
.B(n_1120),
.Y(n_1550)
);

OR2x6_ASAP7_75t_L g1551 ( 
.A(n_1352),
.B(n_936),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1384),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1381),
.B(n_1120),
.Y(n_1553)
);

OAI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1402),
.A2(n_1196),
.B1(n_1218),
.B2(n_1188),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1404),
.B(n_1202),
.Y(n_1555)
);

OAI22xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1438),
.A2(n_898),
.B1(n_900),
.B2(n_896),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1373),
.B(n_1000),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1384),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1384),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1361),
.Y(n_1560)
);

OAI22xp33_ASAP7_75t_R g1561 ( 
.A1(n_1404),
.A2(n_820),
.B1(n_823),
.B2(n_819),
.Y(n_1561)
);

OR2x6_ASAP7_75t_L g1562 ( 
.A(n_1440),
.B(n_1287),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1440),
.A2(n_903),
.B1(n_905),
.B2(n_902),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1364),
.A2(n_908),
.B1(n_909),
.B2(n_906),
.Y(n_1564)
);

OAI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1367),
.A2(n_1220),
.B1(n_1232),
.B2(n_1218),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_SL g1566 ( 
.A1(n_1408),
.A2(n_1232),
.B1(n_1252),
.B2(n_1220),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1445),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1411),
.A2(n_915),
.B1(n_918),
.B2(n_914),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1416),
.Y(n_1569)
);

OA22x2_ASAP7_75t_L g1570 ( 
.A1(n_1429),
.A2(n_922),
.B1(n_965),
.B2(n_935),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1436),
.B(n_828),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1407),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1407),
.Y(n_1573)
);

OAI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1407),
.A2(n_925),
.B1(n_926),
.B2(n_920),
.Y(n_1574)
);

OR2x6_ASAP7_75t_L g1575 ( 
.A(n_1342),
.B(n_1190),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1420),
.A2(n_930),
.B1(n_937),
.B2(n_928),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1444),
.B(n_1202),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1420),
.Y(n_1578)
);

OAI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1420),
.A2(n_940),
.B1(n_947),
.B2(n_938),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1444),
.A2(n_950),
.B1(n_951),
.B2(n_948),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1444),
.B(n_1202),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1342),
.Y(n_1582)
);

OAI22xp33_ASAP7_75t_R g1583 ( 
.A1(n_1342),
.A2(n_837),
.B1(n_853),
.B2(n_832),
.Y(n_1583)
);

OAI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1348),
.A2(n_1258),
.B1(n_1252),
.B2(n_857),
.Y(n_1584)
);

OAI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1348),
.A2(n_1258),
.B1(n_858),
.B2(n_869),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1348),
.B(n_1294),
.Y(n_1586)
);

OR2x6_ASAP7_75t_L g1587 ( 
.A(n_1355),
.B(n_840),
.Y(n_1587)
);

OAI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1355),
.A2(n_953),
.B1(n_955),
.B2(n_952),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1355),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1359),
.A2(n_964),
.B1(n_968),
.B2(n_961),
.Y(n_1590)
);

INVx8_ASAP7_75t_L g1591 ( 
.A(n_1359),
.Y(n_1591)
);

OAI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1359),
.A2(n_864),
.B1(n_895),
.B2(n_892),
.Y(n_1592)
);

OAI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1362),
.A2(n_897),
.B1(n_904),
.B2(n_899),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1334),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1362),
.B(n_1163),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1362),
.A2(n_907),
.B1(n_917),
.B2(n_916),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1363),
.B(n_1186),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1363),
.B(n_1211),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1363),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1375),
.Y(n_1600)
);

OAI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1375),
.A2(n_919),
.B1(n_933),
.B2(n_932),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1375),
.B(n_1211),
.Y(n_1602)
);

OA22x2_ASAP7_75t_L g1603 ( 
.A1(n_1379),
.A2(n_986),
.B1(n_995),
.B2(n_974),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1379),
.A2(n_971),
.B1(n_972),
.B2(n_970),
.Y(n_1604)
);

INVxp33_ASAP7_75t_L g1605 ( 
.A(n_1379),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1389),
.A2(n_975),
.B1(n_976),
.B2(n_973),
.Y(n_1606)
);

XOR2xp5_ASAP7_75t_L g1607 ( 
.A(n_1389),
.B(n_1289),
.Y(n_1607)
);

OR2x6_ASAP7_75t_L g1608 ( 
.A(n_1389),
.B(n_997),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1390),
.Y(n_1609)
);

OAI22xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1390),
.A2(n_978),
.B1(n_988),
.B2(n_977),
.Y(n_1610)
);

OAI22xp33_ASAP7_75t_R g1611 ( 
.A1(n_1390),
.A2(n_942),
.B1(n_944),
.B2(n_941),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1396),
.Y(n_1612)
);

AO22x2_ASAP7_75t_L g1613 ( 
.A1(n_1396),
.A2(n_949),
.B1(n_954),
.B2(n_946),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1396),
.B(n_1312),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1405),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1405),
.Y(n_1616)
);

OAI22xp33_ASAP7_75t_SL g1617 ( 
.A1(n_1405),
.A2(n_991),
.B1(n_992),
.B2(n_989),
.Y(n_1617)
);

OAI22xp33_ASAP7_75t_R g1618 ( 
.A1(n_1421),
.A2(n_962),
.B1(n_966),
.B2(n_960),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1421),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1421),
.A2(n_1003),
.B1(n_1004),
.B2(n_994),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1422),
.A2(n_1006),
.B1(n_1010),
.B2(n_1005),
.Y(n_1621)
);

AO22x2_ASAP7_75t_L g1622 ( 
.A1(n_1422),
.A2(n_979),
.B1(n_981),
.B2(n_969),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1422),
.A2(n_1013),
.B1(n_1016),
.B2(n_1012),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1426),
.B(n_1211),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1426),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1426),
.A2(n_1018),
.B1(n_1022),
.B2(n_1017),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1334),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1334),
.B(n_1288),
.Y(n_1628)
);

OAI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1337),
.A2(n_987),
.B1(n_990),
.B2(n_985),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_SL g1630 ( 
.A1(n_1337),
.A2(n_1025),
.B1(n_1026),
.B2(n_1023),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1337),
.A2(n_1029),
.B1(n_1031),
.B2(n_1027),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_SL g1632 ( 
.A1(n_1338),
.A2(n_1035),
.B1(n_1042),
.B2(n_1034),
.Y(n_1632)
);

AOI22x1_ASAP7_75t_SL g1633 ( 
.A1(n_1338),
.A2(n_1051),
.B1(n_1052),
.B2(n_1049),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1338),
.B(n_1213),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1339),
.B(n_1209),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1339),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1339),
.A2(n_1054),
.B1(n_1055),
.B2(n_1053),
.Y(n_1637)
);

AND2x2_ASAP7_75t_SL g1638 ( 
.A(n_1324),
.B(n_840),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1377),
.Y(n_1639)
);

OAI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1323),
.A2(n_999),
.B1(n_1007),
.B2(n_998),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1351),
.B(n_1213),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1333),
.B(n_1132),
.Y(n_1642)
);

NAND3x1_ASAP7_75t_L g1643 ( 
.A(n_1398),
.B(n_1015),
.C(n_1008),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1377),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1351),
.B(n_1213),
.Y(n_1645)
);

AO22x2_ASAP7_75t_L g1646 ( 
.A1(n_1351),
.A2(n_1285),
.B1(n_1284),
.B2(n_1020),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1351),
.A2(n_1062),
.B1(n_1063),
.B2(n_1058),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1335),
.Y(n_1648)
);

BUFx10_ASAP7_75t_L g1649 ( 
.A(n_1371),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1377),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1351),
.B(n_1308),
.Y(n_1651)
);

OA22x2_ASAP7_75t_L g1652 ( 
.A1(n_1322),
.A2(n_1124),
.B1(n_1136),
.B2(n_1073),
.Y(n_1652)
);

AOI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1351),
.A2(n_1068),
.B1(n_1076),
.B2(n_1065),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1351),
.A2(n_1082),
.B1(n_1086),
.B2(n_1081),
.Y(n_1654)
);

OA22x2_ASAP7_75t_L g1655 ( 
.A1(n_1322),
.A2(n_1110),
.B1(n_1123),
.B2(n_1101),
.Y(n_1655)
);

OAI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1323),
.A2(n_1024),
.B1(n_1032),
.B2(n_1019),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1442),
.B(n_934),
.Y(n_1657)
);

CKINVDCx6p67_ASAP7_75t_R g1658 ( 
.A(n_1323),
.Y(n_1658)
);

OAI22xp33_ASAP7_75t_SL g1659 ( 
.A1(n_1428),
.A2(n_1095),
.B1(n_1097),
.B2(n_1090),
.Y(n_1659)
);

AO22x2_ASAP7_75t_L g1660 ( 
.A1(n_1351),
.A2(n_1037),
.B1(n_1038),
.B2(n_1036),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1335),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1657),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1657),
.Y(n_1663)
);

BUFx2_ASAP7_75t_L g1664 ( 
.A(n_1479),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1489),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1641),
.B(n_1098),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1485),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_1495),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1497),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1528),
.B(n_1205),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1595),
.Y(n_1671)
);

INVx2_ASAP7_75t_SL g1672 ( 
.A(n_1515),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1482),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1483),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1524),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1527),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1484),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1453),
.B(n_1099),
.Y(n_1678)
);

NAND2xp33_ASAP7_75t_SL g1679 ( 
.A(n_1505),
.B(n_1100),
.Y(n_1679)
);

BUFx5_ASAP7_75t_L g1680 ( 
.A(n_1543),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1496),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1500),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1634),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1598),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1602),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1544),
.B(n_1230),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1624),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1448),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1451),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1457),
.B(n_1235),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1458),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1477),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1546),
.B(n_1279),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1510),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1648),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1516),
.B(n_863),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1487),
.B(n_1530),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1661),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1645),
.B(n_1105),
.Y(n_1699)
);

XOR2xp5_ASAP7_75t_L g1700 ( 
.A(n_1446),
.B(n_1290),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1529),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_SL g1702 ( 
.A(n_1551),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_SL g1703 ( 
.A(n_1551),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1468),
.Y(n_1704)
);

NAND2xp33_ASAP7_75t_SL g1705 ( 
.A(n_1516),
.B(n_1293),
.Y(n_1705)
);

OR2x6_ASAP7_75t_L g1706 ( 
.A(n_1515),
.B(n_934),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1535),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1535),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1613),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1613),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1639),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1622),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1622),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1550),
.A2(n_1135),
.B(n_956),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1586),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1614),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1571),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1509),
.Y(n_1718)
);

INVxp33_ASAP7_75t_L g1719 ( 
.A(n_1607),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1509),
.Y(n_1720)
);

AND2x6_ASAP7_75t_L g1721 ( 
.A(n_1553),
.B(n_936),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1658),
.Y(n_1722)
);

CKINVDCx20_ASAP7_75t_R g1723 ( 
.A(n_1491),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1531),
.B(n_1039),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1486),
.B(n_1106),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1628),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1651),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1555),
.B(n_1308),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1447),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1644),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1452),
.B(n_1107),
.Y(n_1731)
);

OR2x2_ASAP7_75t_SL g1732 ( 
.A(n_1469),
.B(n_1044),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1463),
.B(n_1102),
.Y(n_1733)
);

XNOR2xp5_ASAP7_75t_L g1734 ( 
.A(n_1462),
.B(n_1108),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1456),
.B(n_1109),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1650),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1519),
.Y(n_1737)
);

OAI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1549),
.A2(n_1046),
.B(n_1045),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1502),
.B(n_1114),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1517),
.Y(n_1740)
);

INVx1_ASAP7_75t_SL g1741 ( 
.A(n_1511),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1517),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1562),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1562),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1492),
.Y(n_1745)
);

INVxp33_ASAP7_75t_L g1746 ( 
.A(n_1607),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_SL g1747 ( 
.A(n_1638),
.B(n_1115),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1577),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1520),
.B(n_1455),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1461),
.A2(n_997),
.B(n_956),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1581),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1534),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1460),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1646),
.Y(n_1754)
);

CKINVDCx16_ASAP7_75t_R g1755 ( 
.A(n_1649),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1533),
.Y(n_1756)
);

INVxp33_ASAP7_75t_SL g1757 ( 
.A(n_1459),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1646),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1660),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1540),
.B(n_1467),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1472),
.B(n_1116),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1660),
.B(n_1118),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1566),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1642),
.A2(n_1001),
.B(n_1000),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1503),
.B(n_1125),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1570),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1603),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1454),
.A2(n_1040),
.B(n_1001),
.Y(n_1768)
);

XOR2x2_ASAP7_75t_L g1769 ( 
.A(n_1643),
.B(n_27),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1637),
.B(n_1048),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1575),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1475),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1575),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1587),
.Y(n_1774)
);

AND2x6_ASAP7_75t_L g1775 ( 
.A(n_1518),
.B(n_1499),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1587),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1569),
.B(n_1308),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1548),
.B(n_1102),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1608),
.Y(n_1779)
);

NOR2xp67_ASAP7_75t_L g1780 ( 
.A(n_1572),
.B(n_766),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1608),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1488),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1557),
.B(n_1308),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1629),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1503),
.B(n_1126),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1592),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1593),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1504),
.B(n_1129),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1596),
.Y(n_1789)
);

CKINVDCx16_ASAP7_75t_R g1790 ( 
.A(n_1633),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1512),
.B(n_1130),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1576),
.B(n_1057),
.Y(n_1792)
);

NAND2xp33_ASAP7_75t_R g1793 ( 
.A(n_1557),
.B(n_1134),
.Y(n_1793)
);

NOR2xp67_ASAP7_75t_L g1794 ( 
.A(n_1507),
.B(n_767),
.Y(n_1794)
);

CKINVDCx20_ASAP7_75t_R g1795 ( 
.A(n_1647),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1580),
.B(n_1061),
.Y(n_1796)
);

XNOR2x2_ASAP7_75t_L g1797 ( 
.A(n_1476),
.B(n_1069),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1601),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1539),
.B(n_1137),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1480),
.Y(n_1800)
);

BUFx8_ASAP7_75t_L g1801 ( 
.A(n_1498),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1541),
.B(n_1653),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1542),
.B(n_1138),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1492),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1506),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1508),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1514),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1506),
.Y(n_1808)
);

CKINVDCx20_ASAP7_75t_R g1809 ( 
.A(n_1654),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1563),
.B(n_1140),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1471),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1471),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1450),
.B(n_1141),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1564),
.B(n_1145),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1583),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1449),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1611),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1618),
.Y(n_1818)
);

INVxp67_ASAP7_75t_SL g1819 ( 
.A(n_1585),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1630),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1521),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1522),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1513),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1632),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1568),
.B(n_1148),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1476),
.B(n_1149),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1659),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1478),
.B(n_1150),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1635),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1604),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1621),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_SL g1832 ( 
.A(n_1470),
.B(n_1151),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1588),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1610),
.Y(n_1834)
);

NOR2x1p5_ASAP7_75t_L g1835 ( 
.A(n_1464),
.B(n_1152),
.Y(n_1835)
);

INVx2_ASAP7_75t_SL g1836 ( 
.A(n_1652),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1617),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1631),
.Y(n_1838)
);

INVxp33_ASAP7_75t_L g1839 ( 
.A(n_1478),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1655),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1590),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1574),
.B(n_1153),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1579),
.B(n_1154),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1606),
.Y(n_1844)
);

XNOR2xp5_ASAP7_75t_L g1845 ( 
.A(n_1538),
.B(n_1537),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1620),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1560),
.B(n_1157),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1623),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1626),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1513),
.Y(n_1850)
);

AND2x2_ASAP7_75t_SL g1851 ( 
.A(n_1547),
.B(n_1040),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1567),
.B(n_1162),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1597),
.B(n_1089),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1525),
.B(n_1164),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1523),
.Y(n_1855)
);

INVxp33_ASAP7_75t_L g1856 ( 
.A(n_1490),
.Y(n_1856)
);

XOR2xp5_ASAP7_75t_L g1857 ( 
.A(n_1554),
.B(n_1296),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_SL g1858 ( 
.A(n_1545),
.B(n_1165),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1490),
.B(n_1166),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1526),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1532),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1536),
.Y(n_1862)
);

CKINVDCx20_ASAP7_75t_R g1863 ( 
.A(n_1565),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1473),
.B(n_1169),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1561),
.B(n_1171),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1552),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1556),
.B(n_1175),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1474),
.B(n_1176),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1558),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1466),
.B(n_1177),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1559),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1591),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1636),
.A2(n_1071),
.B(n_1060),
.Y(n_1873)
);

XNOR2xp5_ASAP7_75t_L g1874 ( 
.A(n_1465),
.B(n_1178),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1640),
.B(n_1180),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1578),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1573),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1656),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1591),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1481),
.B(n_1182),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1493),
.B(n_1183),
.Y(n_1881)
);

XOR2x2_ASAP7_75t_L g1882 ( 
.A(n_1494),
.B(n_29),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1582),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1605),
.Y(n_1884)
);

OAI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1589),
.A2(n_1600),
.B(n_1599),
.Y(n_1885)
);

XNOR2x2_ASAP7_75t_L g1886 ( 
.A(n_1501),
.B(n_1092),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1584),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1612),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1616),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1619),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1625),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1609),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1615),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1627),
.B(n_1184),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1594),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1594),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1528),
.B(n_1185),
.Y(n_1897)
);

BUFx3_ASAP7_75t_L g1898 ( 
.A(n_1658),
.Y(n_1898)
);

INVxp67_ASAP7_75t_SL g1899 ( 
.A(n_1613),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1657),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1657),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1657),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1595),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1641),
.B(n_1189),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1528),
.B(n_1192),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1657),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1528),
.B(n_1194),
.Y(n_1907)
);

CKINVDCx20_ASAP7_75t_R g1908 ( 
.A(n_1495),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1528),
.B(n_1255),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1528),
.A2(n_1094),
.B(n_1093),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1657),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1657),
.Y(n_1912)
);

XNOR2x1_ASAP7_75t_L g1913 ( 
.A(n_1446),
.B(n_1197),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1657),
.Y(n_1914)
);

CKINVDCx20_ASAP7_75t_R g1915 ( 
.A(n_1495),
.Y(n_1915)
);

OAI21x1_ASAP7_75t_L g1916 ( 
.A1(n_1480),
.A2(n_1071),
.B(n_1060),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1657),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1528),
.B(n_1198),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1657),
.Y(n_1919)
);

BUFx3_ASAP7_75t_L g1920 ( 
.A(n_1658),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1657),
.Y(n_1921)
);

INVxp67_ASAP7_75t_SL g1922 ( 
.A(n_1613),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1658),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1657),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1657),
.Y(n_1925)
);

INVxp33_ASAP7_75t_L g1926 ( 
.A(n_1607),
.Y(n_1926)
);

BUFx6f_ASAP7_75t_L g1927 ( 
.A(n_1575),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1527),
.A2(n_1104),
.B(n_1072),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1657),
.Y(n_1929)
);

OAI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1528),
.A2(n_1133),
.B(n_1121),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1657),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1657),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1657),
.Y(n_1933)
);

XOR2xp5_ASAP7_75t_L g1934 ( 
.A(n_1446),
.B(n_1278),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1657),
.Y(n_1935)
);

BUFx3_ASAP7_75t_L g1936 ( 
.A(n_1658),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1657),
.Y(n_1937)
);

INVx2_ASAP7_75t_SL g1938 ( 
.A(n_1515),
.Y(n_1938)
);

OAI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1527),
.A2(n_1104),
.B(n_1072),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1657),
.Y(n_1940)
);

OAI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1528),
.A2(n_1144),
.B(n_1143),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1528),
.B(n_1199),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1657),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1657),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1479),
.B(n_1147),
.Y(n_1945)
);

BUFx2_ASAP7_75t_L g1946 ( 
.A(n_1479),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1528),
.B(n_1204),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1641),
.B(n_1216),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1657),
.Y(n_1949)
);

XNOR2x2_ASAP7_75t_L g1950 ( 
.A(n_1476),
.B(n_1156),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1657),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1657),
.Y(n_1952)
);

INVxp33_ASAP7_75t_SL g1953 ( 
.A(n_1505),
.Y(n_1953)
);

INVxp67_ASAP7_75t_SL g1954 ( 
.A(n_1613),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1641),
.B(n_1217),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1872),
.Y(n_1956)
);

INVx2_ASAP7_75t_SL g1957 ( 
.A(n_1741),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1741),
.B(n_1675),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1731),
.B(n_1221),
.Y(n_1959)
);

OAI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1916),
.A2(n_1168),
.B(n_1167),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1743),
.B(n_1170),
.Y(n_1961)
);

AND2x4_ASAP7_75t_L g1962 ( 
.A(n_1744),
.B(n_1172),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1667),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1676),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1706),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1669),
.Y(n_1966)
);

INVx2_ASAP7_75t_SL g1967 ( 
.A(n_1706),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1872),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1872),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1721),
.B(n_1223),
.Y(n_1970)
);

AND2x4_ASAP7_75t_L g1971 ( 
.A(n_1737),
.B(n_1174),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1701),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1739),
.B(n_1868),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1721),
.B(n_1224),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1704),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1927),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1711),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1736),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1672),
.B(n_1181),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1721),
.B(n_1227),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1880),
.B(n_1231),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1677),
.Y(n_1982)
);

INVx2_ASAP7_75t_SL g1983 ( 
.A(n_1706),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1927),
.B(n_1234),
.Y(n_1984)
);

INVx4_ASAP7_75t_L g1985 ( 
.A(n_1927),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1729),
.Y(n_1986)
);

AND2x4_ASAP7_75t_L g1987 ( 
.A(n_1938),
.B(n_1187),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1721),
.B(n_1238),
.Y(n_1988)
);

HB1xp67_ASAP7_75t_L g1989 ( 
.A(n_1664),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1946),
.Y(n_1990)
);

INVxp67_ASAP7_75t_L g1991 ( 
.A(n_1899),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1662),
.Y(n_1992)
);

CKINVDCx20_ASAP7_75t_R g1993 ( 
.A(n_1755),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1881),
.B(n_1717),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1663),
.Y(n_1995)
);

OAI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1800),
.A2(n_1195),
.B(n_1191),
.Y(n_1996)
);

AND2x4_ASAP7_75t_L g1997 ( 
.A(n_1697),
.B(n_1200),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1697),
.B(n_1203),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1681),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1683),
.B(n_1206),
.Y(n_2000)
);

INVx3_ASAP7_75t_L g2001 ( 
.A(n_1879),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1762),
.B(n_1240),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1900),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1756),
.B(n_1666),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1901),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1688),
.B(n_1247),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1709),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1756),
.B(n_1699),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1902),
.Y(n_2009)
);

OR2x2_ASAP7_75t_L g2010 ( 
.A(n_1913),
.B(n_1248),
.Y(n_2010)
);

INVx1_ASAP7_75t_SL g2011 ( 
.A(n_1772),
.Y(n_2011)
);

INVx3_ASAP7_75t_L g2012 ( 
.A(n_1806),
.Y(n_2012)
);

OAI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1714),
.A2(n_1212),
.B(n_1208),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1689),
.B(n_1250),
.Y(n_2014)
);

AND2x4_ASAP7_75t_L g2015 ( 
.A(n_1684),
.B(n_1214),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1722),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_1685),
.B(n_1222),
.Y(n_2017)
);

BUFx3_ASAP7_75t_L g2018 ( 
.A(n_1898),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1906),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_1945),
.Y(n_2020)
);

AND2x6_ASAP7_75t_L g2021 ( 
.A(n_1710),
.B(n_1113),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1911),
.Y(n_2022)
);

INVx4_ASAP7_75t_L g2023 ( 
.A(n_1702),
.Y(n_2023)
);

BUFx4f_ASAP7_75t_L g2024 ( 
.A(n_1770),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1904),
.B(n_1948),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1682),
.Y(n_2026)
);

BUFx3_ASAP7_75t_L g2027 ( 
.A(n_1920),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1955),
.B(n_1251),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1691),
.B(n_1253),
.Y(n_2029)
);

AND2x2_ASAP7_75t_SL g2030 ( 
.A(n_1790),
.B(n_963),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1749),
.B(n_1256),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1912),
.Y(n_2032)
);

AND2x6_ASAP7_75t_L g2033 ( 
.A(n_1712),
.B(n_1113),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1826),
.B(n_1259),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1828),
.B(n_1260),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1807),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1821),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1692),
.B(n_1261),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1694),
.B(n_1695),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_1945),
.Y(n_2040)
);

BUFx3_ASAP7_75t_L g2041 ( 
.A(n_1936),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1705),
.B(n_1262),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1822),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1859),
.B(n_1264),
.Y(n_2044)
);

BUFx5_ASAP7_75t_L g2045 ( 
.A(n_1727),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1813),
.B(n_1265),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1835),
.B(n_1266),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1698),
.B(n_1268),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1914),
.Y(n_2049)
);

INVx3_ASAP7_75t_L g2050 ( 
.A(n_1855),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1876),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1815),
.B(n_1269),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1917),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_1922),
.Y(n_2054)
);

INVx3_ASAP7_75t_L g2055 ( 
.A(n_1730),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1910),
.B(n_1270),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1817),
.B(n_1271),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1673),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1910),
.B(n_1272),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1674),
.Y(n_2060)
);

AND2x6_ASAP7_75t_L g2061 ( 
.A(n_1713),
.B(n_1122),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1678),
.B(n_1799),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_1923),
.Y(n_2063)
);

INVxp67_ASAP7_75t_L g2064 ( 
.A(n_1954),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_1757),
.B(n_1274),
.Y(n_2065)
);

OAI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1928),
.A2(n_1233),
.B(n_1225),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1818),
.B(n_1276),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1930),
.B(n_1280),
.Y(n_2068)
);

OAI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_1930),
.A2(n_1237),
.B(n_1236),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1865),
.B(n_1282),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1680),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1941),
.B(n_1286),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1919),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_1687),
.B(n_1239),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1845),
.B(n_1297),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1874),
.B(n_1299),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1765),
.B(n_1302),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_1860),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_1857),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_1766),
.B(n_1241),
.Y(n_2080)
);

BUFx6f_ASAP7_75t_L g2081 ( 
.A(n_1861),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1941),
.B(n_1303),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1921),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1785),
.B(n_1307),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1753),
.B(n_1243),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_1754),
.B(n_1245),
.Y(n_2086)
);

INVxp67_ASAP7_75t_L g2087 ( 
.A(n_1905),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1918),
.B(n_1947),
.Y(n_2088)
);

AND2x2_ASAP7_75t_SL g2089 ( 
.A(n_1745),
.B(n_1122),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1924),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1878),
.B(n_1246),
.Y(n_2091)
);

OAI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1728),
.A2(n_1254),
.B(n_1249),
.Y(n_2092)
);

INVx4_ASAP7_75t_L g2093 ( 
.A(n_1702),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_1758),
.B(n_1263),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1680),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1925),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_1759),
.B(n_1267),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1929),
.Y(n_2098)
);

BUFx3_ASAP7_75t_L g2099 ( 
.A(n_1801),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1738),
.B(n_1275),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1931),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_1707),
.A2(n_1281),
.B1(n_1277),
.B2(n_1193),
.Y(n_2102)
);

AND2x2_ASAP7_75t_SL g2103 ( 
.A(n_1832),
.B(n_1190),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1680),
.Y(n_2104)
);

NAND2x1p5_ASAP7_75t_L g2105 ( 
.A(n_1708),
.B(n_1193),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1680),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1932),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_1724),
.B(n_1210),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_1851),
.B(n_1210),
.Y(n_2109)
);

INVx2_ASAP7_75t_SL g2110 ( 
.A(n_1724),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1738),
.B(n_1215),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1933),
.Y(n_2112)
);

INVx3_ASAP7_75t_L g2113 ( 
.A(n_1752),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1935),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1784),
.B(n_1215),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1786),
.B(n_1242),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1862),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1937),
.Y(n_2118)
);

BUFx6f_ASAP7_75t_L g2119 ( 
.A(n_1866),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1680),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1940),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1943),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1735),
.B(n_1242),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_L g2124 ( 
.A(n_1788),
.B(n_1283),
.Y(n_2124)
);

OAI21x1_ASAP7_75t_L g2125 ( 
.A1(n_1885),
.A2(n_1287),
.B(n_1283),
.Y(n_2125)
);

INVx3_ASAP7_75t_L g2126 ( 
.A(n_1869),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1871),
.Y(n_2127)
);

OR2x2_ASAP7_75t_L g2128 ( 
.A(n_1700),
.B(n_29),
.Y(n_2128)
);

AND2x4_ASAP7_75t_L g2129 ( 
.A(n_1748),
.B(n_1255),
.Y(n_2129)
);

INVx2_ASAP7_75t_SL g2130 ( 
.A(n_1853),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_1751),
.B(n_1255),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_1671),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_1734),
.B(n_1255),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1787),
.B(n_1257),
.Y(n_2134)
);

OAI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_1939),
.A2(n_1257),
.B(n_756),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1715),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_1801),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1839),
.B(n_1856),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1882),
.B(n_1257),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_1703),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1716),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1789),
.B(n_1257),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1863),
.B(n_30),
.Y(n_2143)
);

AND2x4_ASAP7_75t_L g2144 ( 
.A(n_1782),
.B(n_30),
.Y(n_2144)
);

OAI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_1726),
.A2(n_757),
.B(n_755),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1944),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_1934),
.B(n_31),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_1897),
.B(n_32),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1665),
.Y(n_2149)
);

HB1xp67_ASAP7_75t_L g2150 ( 
.A(n_1703),
.Y(n_2150)
);

AND2x6_ASAP7_75t_L g2151 ( 
.A(n_1740),
.B(n_758),
.Y(n_2151)
);

OAI21xp5_ASAP7_75t_L g2152 ( 
.A1(n_1873),
.A2(n_1783),
.B(n_1733),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1949),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1951),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1798),
.B(n_1838),
.Y(n_2155)
);

HB1xp67_ASAP7_75t_L g2156 ( 
.A(n_1772),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1841),
.B(n_33),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_1907),
.B(n_33),
.Y(n_2158)
);

NAND2x1p5_ASAP7_75t_L g2159 ( 
.A(n_1771),
.B(n_34),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1844),
.B(n_35),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1846),
.B(n_36),
.Y(n_2161)
);

INVx1_ASAP7_75t_SL g2162 ( 
.A(n_1805),
.Y(n_2162)
);

INVx2_ASAP7_75t_SL g2163 ( 
.A(n_1853),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_1942),
.B(n_36),
.Y(n_2164)
);

BUFx3_ASAP7_75t_L g2165 ( 
.A(n_1953),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1848),
.B(n_37),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1849),
.B(n_37),
.Y(n_2167)
);

INVx3_ASAP7_75t_SL g2168 ( 
.A(n_1732),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1903),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_1793),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1952),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_R g2172 ( 
.A(n_1679),
.B(n_1832),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_1773),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_1791),
.B(n_38),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_1792),
.B(n_1796),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1718),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_1792),
.B(n_38),
.Y(n_2177)
);

INVx2_ASAP7_75t_SL g2178 ( 
.A(n_1774),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1796),
.B(n_40),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1720),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1894),
.Y(n_2181)
);

HB1xp67_ASAP7_75t_L g2182 ( 
.A(n_1805),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1767),
.Y(n_2183)
);

BUFx6f_ASAP7_75t_L g2184 ( 
.A(n_1909),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1819),
.B(n_1764),
.Y(n_2185)
);

BUFx6f_ASAP7_75t_L g2186 ( 
.A(n_1776),
.Y(n_2186)
);

INVx8_ASAP7_75t_L g2187 ( 
.A(n_1775),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_1816),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1895),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_1823),
.B(n_41),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1887),
.B(n_41),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1742),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1670),
.B(n_42),
.Y(n_2193)
);

INVx2_ASAP7_75t_SL g2194 ( 
.A(n_1779),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1895),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1888),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_1823),
.B(n_42),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_1802),
.B(n_43),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1778),
.B(n_44),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1750),
.Y(n_2200)
);

INVx3_ASAP7_75t_L g2201 ( 
.A(n_1781),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1833),
.Y(n_2202)
);

OAI21x1_ASAP7_75t_L g2203 ( 
.A1(n_1885),
.A2(n_761),
.B(n_760),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_1814),
.B(n_45),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1760),
.B(n_45),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_1768),
.B(n_46),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1890),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1891),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_1825),
.B(n_47),
.Y(n_2209)
);

XOR2xp5_ASAP7_75t_L g2210 ( 
.A(n_1723),
.B(n_47),
.Y(n_2210)
);

INVx4_ASAP7_75t_L g2211 ( 
.A(n_1827),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_1797),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1834),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_1747),
.B(n_49),
.Y(n_2214)
);

INVx3_ASAP7_75t_L g2215 ( 
.A(n_1884),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1837),
.Y(n_2216)
);

INVx3_ASAP7_75t_L g2217 ( 
.A(n_1877),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_1747),
.B(n_49),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1811),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1812),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_1668),
.Y(n_2221)
);

INVx1_ASAP7_75t_SL g2222 ( 
.A(n_1847),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1840),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_1864),
.B(n_50),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1883),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1896),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_1836),
.Y(n_2227)
);

INVx2_ASAP7_75t_SL g2228 ( 
.A(n_1690),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1889),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_1686),
.B(n_50),
.Y(n_2230)
);

OAI21xp33_ASAP7_75t_L g2231 ( 
.A1(n_1804),
.A2(n_1808),
.B(n_1725),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1829),
.Y(n_2232)
);

INVx2_ASAP7_75t_SL g2233 ( 
.A(n_1886),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1850),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1852),
.Y(n_2235)
);

BUFx6f_ASAP7_75t_L g2236 ( 
.A(n_1777),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1693),
.B(n_51),
.Y(n_2237)
);

INVx2_ASAP7_75t_SL g2238 ( 
.A(n_1696),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1775),
.B(n_53),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_SL g2240 ( 
.A(n_1820),
.B(n_53),
.Y(n_2240)
);

AND2x4_ASAP7_75t_L g2241 ( 
.A(n_1824),
.B(n_54),
.Y(n_2241)
);

NAND2x1p5_ASAP7_75t_L g2242 ( 
.A(n_1830),
.B(n_54),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1892),
.Y(n_2243)
);

OAI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_1780),
.A2(n_769),
.B(n_763),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1950),
.Y(n_2245)
);

AND2x4_ASAP7_75t_L g2246 ( 
.A(n_1831),
.B(n_55),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1893),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_1875),
.B(n_55),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1803),
.Y(n_2249)
);

AND2x4_ASAP7_75t_L g2250 ( 
.A(n_1761),
.B(n_56),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1810),
.Y(n_2251)
);

INVxp67_ASAP7_75t_L g2252 ( 
.A(n_1858),
.Y(n_2252)
);

INVx2_ASAP7_75t_SL g2253 ( 
.A(n_1775),
.Y(n_2253)
);

AND2x4_ASAP7_75t_L g2254 ( 
.A(n_1775),
.B(n_57),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1867),
.B(n_57),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1854),
.Y(n_2256)
);

INVxp67_ASAP7_75t_L g2257 ( 
.A(n_1858),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1870),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_L g2259 ( 
.A(n_1842),
.B(n_58),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1843),
.Y(n_2260)
);

BUFx3_ASAP7_75t_L g2261 ( 
.A(n_1795),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1780),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1794),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_1719),
.B(n_58),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1769),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1794),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1809),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1763),
.B(n_59),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1746),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_1926),
.B(n_59),
.Y(n_2270)
);

BUFx3_ASAP7_75t_L g2271 ( 
.A(n_1908),
.Y(n_2271)
);

INVx4_ASAP7_75t_L g2272 ( 
.A(n_1915),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_1741),
.B(n_60),
.Y(n_2273)
);

BUFx2_ASAP7_75t_L g2274 ( 
.A(n_1675),
.Y(n_2274)
);

BUFx3_ASAP7_75t_L g2275 ( 
.A(n_1729),
.Y(n_2275)
);

INVxp67_ASAP7_75t_SL g2276 ( 
.A(n_1899),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_1741),
.B(n_60),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_1741),
.B(n_61),
.Y(n_2278)
);

AND2x2_ASAP7_75t_SL g2279 ( 
.A(n_1755),
.B(n_62),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_1741),
.B(n_62),
.Y(n_2280)
);

BUFx4f_ASAP7_75t_L g2281 ( 
.A(n_1706),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_1741),
.B(n_63),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_SL g2283 ( 
.A(n_1927),
.B(n_63),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1676),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1667),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_1741),
.B(n_64),
.Y(n_2286)
);

HB1xp67_ASAP7_75t_L g2287 ( 
.A(n_1741),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_1676),
.Y(n_2288)
);

HB1xp67_ASAP7_75t_L g2289 ( 
.A(n_1741),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_1741),
.B(n_64),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1721),
.B(n_65),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_1743),
.B(n_65),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1667),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_1741),
.B(n_66),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1721),
.B(n_66),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_1741),
.B(n_68),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2136),
.Y(n_2297)
);

INVx3_ASAP7_75t_L g2298 ( 
.A(n_1976),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_2062),
.B(n_68),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2141),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_1964),
.Y(n_2301)
);

NOR2xp33_ASAP7_75t_SL g2302 ( 
.A(n_2103),
.B(n_771),
.Y(n_2302)
);

OR2x6_ASAP7_75t_L g2303 ( 
.A(n_2099),
.B(n_69),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1972),
.Y(n_2304)
);

AND2x4_ASAP7_75t_L g2305 ( 
.A(n_1957),
.B(n_70),
.Y(n_2305)
);

CKINVDCx6p67_ASAP7_75t_R g2306 ( 
.A(n_2137),
.Y(n_2306)
);

NAND2x1p5_ASAP7_75t_L g2307 ( 
.A(n_2281),
.B(n_71),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2284),
.Y(n_2308)
);

NAND2x1_ASAP7_75t_L g2309 ( 
.A(n_1976),
.B(n_773),
.Y(n_2309)
);

OR2x6_ASAP7_75t_L g2310 ( 
.A(n_2023),
.B(n_70),
.Y(n_2310)
);

NAND2x1p5_ASAP7_75t_L g2311 ( 
.A(n_2281),
.B(n_73),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_1958),
.B(n_72),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2039),
.Y(n_2313)
);

AND2x4_ASAP7_75t_L g2314 ( 
.A(n_2287),
.B(n_72),
.Y(n_2314)
);

BUFx6f_ASAP7_75t_L g2315 ( 
.A(n_1976),
.Y(n_2315)
);

BUFx3_ASAP7_75t_L g2316 ( 
.A(n_2275),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2289),
.B(n_74),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2288),
.Y(n_2318)
);

BUFx6f_ASAP7_75t_L g2319 ( 
.A(n_1969),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_1994),
.B(n_74),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2175),
.B(n_75),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2039),
.Y(n_2322)
);

INVx3_ASAP7_75t_L g2323 ( 
.A(n_1969),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2045),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_SL g2325 ( 
.A(n_2151),
.B(n_774),
.Y(n_2325)
);

INVx4_ASAP7_75t_L g2326 ( 
.A(n_1969),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2232),
.Y(n_2327)
);

AND2x6_ASAP7_75t_L g2328 ( 
.A(n_2254),
.B(n_76),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2011),
.B(n_76),
.Y(n_2329)
);

BUFx4f_ASAP7_75t_L g2330 ( 
.A(n_2279),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2011),
.B(n_77),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2088),
.B(n_77),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1982),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2004),
.B(n_78),
.Y(n_2334)
);

CKINVDCx20_ASAP7_75t_R g2335 ( 
.A(n_1993),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_2274),
.B(n_78),
.Y(n_2336)
);

OR2x6_ASAP7_75t_L g2337 ( 
.A(n_2023),
.B(n_79),
.Y(n_2337)
);

CKINVDCx11_ASAP7_75t_R g2338 ( 
.A(n_2093),
.Y(n_2338)
);

BUFx6f_ASAP7_75t_L g2339 ( 
.A(n_1985),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2008),
.B(n_79),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_SL g2341 ( 
.A(n_2151),
.B(n_779),
.Y(n_2341)
);

BUFx2_ASAP7_75t_L g2342 ( 
.A(n_1989),
.Y(n_2342)
);

AND2x4_ASAP7_75t_L g2343 ( 
.A(n_2253),
.B(n_80),
.Y(n_2343)
);

BUFx3_ASAP7_75t_L g2344 ( 
.A(n_2018),
.Y(n_2344)
);

OR2x2_ASAP7_75t_L g2345 ( 
.A(n_2010),
.B(n_80),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2045),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2045),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2045),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1999),
.Y(n_2349)
);

AND2x4_ASAP7_75t_L g2350 ( 
.A(n_2235),
.B(n_82),
.Y(n_2350)
);

NOR2x1_ASAP7_75t_L g2351 ( 
.A(n_2239),
.B(n_84),
.Y(n_2351)
);

AND2x4_ASAP7_75t_L g2352 ( 
.A(n_2217),
.B(n_85),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2196),
.Y(n_2353)
);

AND2x4_ASAP7_75t_L g2354 ( 
.A(n_2217),
.B(n_86),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2075),
.B(n_87),
.Y(n_2355)
);

INVx3_ASAP7_75t_L g2356 ( 
.A(n_1985),
.Y(n_2356)
);

HB1xp67_ASAP7_75t_L g2357 ( 
.A(n_2156),
.Y(n_2357)
);

BUFx2_ASAP7_75t_L g2358 ( 
.A(n_1990),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_2078),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_1986),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2031),
.B(n_88),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_1973),
.B(n_88),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2045),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_2020),
.Y(n_2364)
);

INVx5_ASAP7_75t_L g2365 ( 
.A(n_2093),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2046),
.B(n_1981),
.Y(n_2366)
);

INVx3_ASAP7_75t_L g2367 ( 
.A(n_2078),
.Y(n_2367)
);

BUFx2_ASAP7_75t_L g2368 ( 
.A(n_1965),
.Y(n_2368)
);

BUFx6f_ASAP7_75t_L g2369 ( 
.A(n_2078),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_L g2370 ( 
.A(n_2087),
.B(n_89),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2207),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2172),
.B(n_90),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2026),
.Y(n_2373)
);

BUFx3_ASAP7_75t_L g2374 ( 
.A(n_2027),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2208),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2192),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2139),
.B(n_90),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2007),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2155),
.B(n_91),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2007),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2007),
.Y(n_2381)
);

BUFx2_ASAP7_75t_L g2382 ( 
.A(n_1965),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2087),
.B(n_91),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2134),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2025),
.B(n_92),
.Y(n_2385)
);

INVx3_ASAP7_75t_L g2386 ( 
.A(n_2081),
.Y(n_2386)
);

BUFx6f_ASAP7_75t_L g2387 ( 
.A(n_2081),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2109),
.B(n_92),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2058),
.Y(n_2389)
);

AND2x4_ASAP7_75t_L g2390 ( 
.A(n_1967),
.B(n_93),
.Y(n_2390)
);

INVx3_ASAP7_75t_L g2391 ( 
.A(n_2081),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2060),
.Y(n_2392)
);

BUFx12f_ASAP7_75t_L g2393 ( 
.A(n_2140),
.Y(n_2393)
);

NAND2x1p5_ASAP7_75t_L g2394 ( 
.A(n_2041),
.B(n_2024),
.Y(n_2394)
);

AND2x4_ASAP7_75t_L g2395 ( 
.A(n_1983),
.B(n_94),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2134),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2142),
.Y(n_2397)
);

AND2x4_ASAP7_75t_L g2398 ( 
.A(n_2222),
.B(n_94),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2056),
.B(n_95),
.Y(n_2399)
);

AND2x6_ASAP7_75t_L g2400 ( 
.A(n_2254),
.B(n_96),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2056),
.B(n_96),
.Y(n_2401)
);

NAND2x1p5_ASAP7_75t_L g2402 ( 
.A(n_2024),
.B(n_98),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2059),
.B(n_2068),
.Y(n_2403)
);

OR2x2_ASAP7_75t_L g2404 ( 
.A(n_2267),
.B(n_97),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_2222),
.B(n_97),
.Y(n_2405)
);

INVx5_ASAP7_75t_L g2406 ( 
.A(n_2151),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2142),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2002),
.B(n_99),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2206),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2206),
.Y(n_2410)
);

BUFx6f_ASAP7_75t_L g2411 ( 
.A(n_2117),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2059),
.B(n_100),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2125),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2076),
.B(n_100),
.Y(n_2414)
);

OR2x6_ASAP7_75t_L g2415 ( 
.A(n_2187),
.B(n_102),
.Y(n_2415)
);

BUFx8_ASAP7_75t_SL g2416 ( 
.A(n_2016),
.Y(n_2416)
);

NAND2x1p5_ASAP7_75t_L g2417 ( 
.A(n_2063),
.B(n_2165),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2070),
.B(n_102),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2127),
.Y(n_2419)
);

AND2x4_ASAP7_75t_L g2420 ( 
.A(n_2130),
.B(n_103),
.Y(n_2420)
);

INVxp67_ASAP7_75t_L g2421 ( 
.A(n_2040),
.Y(n_2421)
);

AND2x4_ASAP7_75t_L g2422 ( 
.A(n_2163),
.B(n_2228),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2219),
.Y(n_2423)
);

BUFx3_ASAP7_75t_L g2424 ( 
.A(n_2150),
.Y(n_2424)
);

BUFx2_ASAP7_75t_L g2425 ( 
.A(n_2292),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_SL g2426 ( 
.A(n_2151),
.B(n_780),
.Y(n_2426)
);

AND2x4_ASAP7_75t_L g2427 ( 
.A(n_2181),
.B(n_104),
.Y(n_2427)
);

BUFx6f_ASAP7_75t_L g2428 ( 
.A(n_2117),
.Y(n_2428)
);

NOR2x1_ASAP7_75t_L g2429 ( 
.A(n_2239),
.B(n_2291),
.Y(n_2429)
);

BUFx4f_ASAP7_75t_L g2430 ( 
.A(n_2030),
.Y(n_2430)
);

BUFx2_ASAP7_75t_L g2431 ( 
.A(n_2292),
.Y(n_2431)
);

BUFx4_ASAP7_75t_SL g2432 ( 
.A(n_2269),
.Y(n_2432)
);

INVx3_ASAP7_75t_L g2433 ( 
.A(n_2117),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2068),
.B(n_106),
.Y(n_2434)
);

AND2x4_ASAP7_75t_L g2435 ( 
.A(n_2256),
.B(n_106),
.Y(n_2435)
);

AND2x4_ASAP7_75t_L g2436 ( 
.A(n_2149),
.B(n_107),
.Y(n_2436)
);

INVxp67_ASAP7_75t_L g2437 ( 
.A(n_2273),
.Y(n_2437)
);

INVx3_ASAP7_75t_L g2438 ( 
.A(n_2119),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2072),
.B(n_2082),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2243),
.Y(n_2440)
);

NAND2x1p5_ASAP7_75t_L g2441 ( 
.A(n_1956),
.B(n_109),
.Y(n_2441)
);

NAND2x1p5_ASAP7_75t_L g2442 ( 
.A(n_1956),
.B(n_110),
.Y(n_2442)
);

NAND2x1p5_ASAP7_75t_L g2443 ( 
.A(n_1968),
.B(n_111),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2072),
.B(n_107),
.Y(n_2444)
);

BUFx6f_ASAP7_75t_L g2445 ( 
.A(n_2119),
.Y(n_2445)
);

HB1xp67_ASAP7_75t_L g2446 ( 
.A(n_2110),
.Y(n_2446)
);

OR2x2_ASAP7_75t_L g2447 ( 
.A(n_2079),
.B(n_112),
.Y(n_2447)
);

AND2x4_ASAP7_75t_L g2448 ( 
.A(n_2173),
.B(n_112),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2247),
.Y(n_2449)
);

INVx3_ASAP7_75t_L g2450 ( 
.A(n_2119),
.Y(n_2450)
);

INVx3_ASAP7_75t_L g2451 ( 
.A(n_2186),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_2065),
.B(n_113),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2082),
.B(n_113),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2220),
.Y(n_2454)
);

BUFx3_ASAP7_75t_L g2455 ( 
.A(n_1968),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2036),
.Y(n_2456)
);

AND2x4_ASAP7_75t_L g2457 ( 
.A(n_2173),
.B(n_114),
.Y(n_2457)
);

AND2x2_ASAP7_75t_SL g2458 ( 
.A(n_2089),
.B(n_115),
.Y(n_2458)
);

NOR2x1_ASAP7_75t_L g2459 ( 
.A(n_2291),
.B(n_115),
.Y(n_2459)
);

CKINVDCx6p67_ASAP7_75t_R g2460 ( 
.A(n_2168),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2143),
.B(n_116),
.Y(n_2461)
);

AND2x4_ASAP7_75t_L g2462 ( 
.A(n_2201),
.B(n_117),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_1959),
.B(n_117),
.Y(n_2463)
);

INVxp67_ASAP7_75t_L g2464 ( 
.A(n_2277),
.Y(n_2464)
);

AND2x2_ASAP7_75t_SL g2465 ( 
.A(n_2241),
.B(n_2246),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2037),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2069),
.B(n_2198),
.Y(n_2467)
);

BUFx8_ASAP7_75t_L g2468 ( 
.A(n_2241),
.Y(n_2468)
);

NAND2x1p5_ASAP7_75t_L g2469 ( 
.A(n_2144),
.B(n_120),
.Y(n_2469)
);

INVx5_ASAP7_75t_L g2470 ( 
.A(n_2021),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2043),
.Y(n_2471)
);

AND2x4_ASAP7_75t_L g2472 ( 
.A(n_2201),
.B(n_119),
.Y(n_2472)
);

OR2x2_ASAP7_75t_L g2473 ( 
.A(n_2128),
.B(n_120),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2028),
.B(n_122),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2051),
.Y(n_2475)
);

BUFx3_ASAP7_75t_L g2476 ( 
.A(n_2261),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2034),
.B(n_122),
.Y(n_2477)
);

BUFx6f_ASAP7_75t_L g2478 ( 
.A(n_2132),
.Y(n_2478)
);

NAND2x1p5_ASAP7_75t_L g2479 ( 
.A(n_2144),
.B(n_2246),
.Y(n_2479)
);

CKINVDCx20_ASAP7_75t_R g2480 ( 
.A(n_2170),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2200),
.Y(n_2481)
);

INVxp67_ASAP7_75t_L g2482 ( 
.A(n_2278),
.Y(n_2482)
);

BUFx2_ASAP7_75t_L g2483 ( 
.A(n_1979),
.Y(n_2483)
);

INVxp67_ASAP7_75t_SL g2484 ( 
.A(n_1991),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_1963),
.Y(n_2485)
);

OR2x2_ASAP7_75t_L g2486 ( 
.A(n_2265),
.B(n_123),
.Y(n_2486)
);

INVx1_ASAP7_75t_SL g2487 ( 
.A(n_2054),
.Y(n_2487)
);

HB1xp67_ASAP7_75t_L g2488 ( 
.A(n_2296),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_1966),
.Y(n_2489)
);

CKINVDCx8_ASAP7_75t_R g2490 ( 
.A(n_2187),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2069),
.B(n_123),
.Y(n_2491)
);

BUFx2_ASAP7_75t_L g2492 ( 
.A(n_1979),
.Y(n_2492)
);

AND2x4_ASAP7_75t_L g2493 ( 
.A(n_2249),
.B(n_124),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2202),
.B(n_126),
.Y(n_2494)
);

NOR2x1_ASAP7_75t_L g2495 ( 
.A(n_2295),
.B(n_126),
.Y(n_2495)
);

INVxp67_ASAP7_75t_L g2496 ( 
.A(n_2280),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_2258),
.B(n_127),
.Y(n_2497)
);

NOR2xp33_ASAP7_75t_L g2498 ( 
.A(n_2260),
.B(n_2077),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2213),
.B(n_128),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2035),
.B(n_129),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2234),
.Y(n_2501)
);

BUFx12f_ASAP7_75t_L g2502 ( 
.A(n_2227),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_SL g2503 ( 
.A(n_2187),
.B(n_781),
.Y(n_2503)
);

CKINVDCx6p67_ASAP7_75t_R g2504 ( 
.A(n_2271),
.Y(n_2504)
);

BUFx2_ASAP7_75t_L g2505 ( 
.A(n_1987),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2216),
.B(n_129),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2251),
.B(n_2085),
.Y(n_2507)
);

AND2x6_ASAP7_75t_L g2508 ( 
.A(n_2295),
.B(n_130),
.Y(n_2508)
);

OR2x6_ASAP7_75t_L g2509 ( 
.A(n_2159),
.B(n_130),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2044),
.B(n_2177),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2179),
.B(n_2147),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2085),
.B(n_131),
.Y(n_2512)
);

NAND2x1p5_ASAP7_75t_L g2513 ( 
.A(n_2186),
.B(n_134),
.Y(n_2513)
);

INVxp67_ASAP7_75t_L g2514 ( 
.A(n_2282),
.Y(n_2514)
);

AND2x4_ASAP7_75t_L g2515 ( 
.A(n_2086),
.B(n_133),
.Y(n_2515)
);

BUFx2_ASAP7_75t_L g2516 ( 
.A(n_1987),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_1992),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_SL g2518 ( 
.A(n_1991),
.B(n_782),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2155),
.B(n_135),
.Y(n_2519)
);

OR2x6_ASAP7_75t_L g2520 ( 
.A(n_2159),
.B(n_2242),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_1995),
.Y(n_2521)
);

HB1xp67_ASAP7_75t_L g2522 ( 
.A(n_2294),
.Y(n_2522)
);

NOR2xp33_ASAP7_75t_SL g2523 ( 
.A(n_2064),
.B(n_783),
.Y(n_2523)
);

BUFx6f_ASAP7_75t_L g2524 ( 
.A(n_2132),
.Y(n_2524)
);

BUFx4f_ASAP7_75t_L g2525 ( 
.A(n_2242),
.Y(n_2525)
);

AND2x4_ASAP7_75t_L g2526 ( 
.A(n_2086),
.B(n_135),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_SL g2527 ( 
.A(n_2064),
.B(n_784),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2185),
.B(n_137),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2094),
.B(n_137),
.Y(n_2529)
);

OR2x6_ASAP7_75t_L g2530 ( 
.A(n_2272),
.B(n_140),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2094),
.B(n_140),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2003),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2097),
.B(n_141),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2285),
.Y(n_2534)
);

BUFx4f_ASAP7_75t_L g2535 ( 
.A(n_2227),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2084),
.B(n_142),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2005),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2052),
.B(n_142),
.Y(n_2538)
);

BUFx4f_ASAP7_75t_L g2539 ( 
.A(n_2227),
.Y(n_2539)
);

CKINVDCx20_ASAP7_75t_R g2540 ( 
.A(n_2221),
.Y(n_2540)
);

BUFx2_ASAP7_75t_L g2541 ( 
.A(n_2286),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2097),
.B(n_143),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2009),
.Y(n_2543)
);

INVx4_ASAP7_75t_L g2544 ( 
.A(n_2021),
.Y(n_2544)
);

OR2x6_ASAP7_75t_L g2545 ( 
.A(n_2272),
.B(n_143),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2123),
.B(n_145),
.Y(n_2546)
);

BUFx2_ASAP7_75t_L g2547 ( 
.A(n_2290),
.Y(n_2547)
);

NOR2xp33_ASAP7_75t_SL g2548 ( 
.A(n_2252),
.B(n_785),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2185),
.B(n_145),
.Y(n_2549)
);

INVx6_ASAP7_75t_L g2550 ( 
.A(n_2186),
.Y(n_2550)
);

INVxp67_ASAP7_75t_SL g2551 ( 
.A(n_2276),
.Y(n_2551)
);

OR2x2_ASAP7_75t_L g2552 ( 
.A(n_2108),
.B(n_146),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2293),
.Y(n_2553)
);

NAND2xp33_ASAP7_75t_L g2554 ( 
.A(n_2021),
.B(n_787),
.Y(n_2554)
);

CKINVDCx8_ASAP7_75t_R g2555 ( 
.A(n_2188),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2057),
.B(n_146),
.Y(n_2556)
);

INVx1_ASAP7_75t_SL g2557 ( 
.A(n_2162),
.Y(n_2557)
);

OR2x2_ASAP7_75t_L g2558 ( 
.A(n_2108),
.B(n_147),
.Y(n_2558)
);

INVx3_ASAP7_75t_L g2559 ( 
.A(n_2132),
.Y(n_2559)
);

AND2x2_ASAP7_75t_SL g2560 ( 
.A(n_2214),
.B(n_147),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_2067),
.B(n_148),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2091),
.B(n_148),
.Y(n_2562)
);

AND2x4_ASAP7_75t_L g2563 ( 
.A(n_2215),
.B(n_149),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2225),
.Y(n_2564)
);

INVxp67_ASAP7_75t_L g2565 ( 
.A(n_2182),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_L g2566 ( 
.A(n_2238),
.B(n_150),
.Y(n_2566)
);

BUFx3_ASAP7_75t_L g2567 ( 
.A(n_2001),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2229),
.Y(n_2568)
);

INVx3_ASAP7_75t_L g2569 ( 
.A(n_2169),
.Y(n_2569)
);

AND2x4_ASAP7_75t_L g2570 ( 
.A(n_2215),
.B(n_150),
.Y(n_2570)
);

OR2x2_ASAP7_75t_L g2571 ( 
.A(n_2138),
.B(n_151),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2204),
.B(n_153),
.Y(n_2572)
);

OR2x6_ASAP7_75t_L g2573 ( 
.A(n_2211),
.B(n_153),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2209),
.B(n_155),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2248),
.B(n_155),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2006),
.B(n_2014),
.Y(n_2576)
);

NAND2x1p5_ASAP7_75t_L g2577 ( 
.A(n_2055),
.B(n_157),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_2211),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2133),
.B(n_156),
.Y(n_2579)
);

BUFx3_ASAP7_75t_L g2580 ( 
.A(n_2001),
.Y(n_2580)
);

BUFx2_ASAP7_75t_L g2581 ( 
.A(n_2021),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2019),
.Y(n_2582)
);

BUFx12f_ASAP7_75t_L g2583 ( 
.A(n_1997),
.Y(n_2583)
);

AND2x4_ASAP7_75t_L g2584 ( 
.A(n_2148),
.B(n_156),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2006),
.B(n_157),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2022),
.Y(n_2586)
);

BUFx6f_ASAP7_75t_L g2587 ( 
.A(n_2169),
.Y(n_2587)
);

NOR2x1_ASAP7_75t_L g2588 ( 
.A(n_2255),
.B(n_158),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2233),
.B(n_159),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_1975),
.Y(n_2590)
);

NOR2xp33_ASAP7_75t_L g2591 ( 
.A(n_2014),
.B(n_159),
.Y(n_2591)
);

INVx2_ASAP7_75t_SL g2592 ( 
.A(n_1997),
.Y(n_2592)
);

NOR2x1_ASAP7_75t_L g2593 ( 
.A(n_2255),
.B(n_160),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_1977),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2029),
.B(n_160),
.Y(n_2595)
);

INVx4_ASAP7_75t_L g2596 ( 
.A(n_2033),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_1998),
.B(n_1971),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_1998),
.B(n_162),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2029),
.B(n_162),
.Y(n_2599)
);

NOR2xp33_ASAP7_75t_L g2600 ( 
.A(n_2038),
.B(n_163),
.Y(n_2600)
);

AND2x4_ASAP7_75t_L g2601 ( 
.A(n_2158),
.B(n_163),
.Y(n_2601)
);

BUFx2_ASAP7_75t_L g2602 ( 
.A(n_2033),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_1971),
.B(n_164),
.Y(n_2603)
);

BUFx6f_ASAP7_75t_L g2604 ( 
.A(n_2169),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2080),
.B(n_164),
.Y(n_2605)
);

NAND2x1p5_ASAP7_75t_L g2606 ( 
.A(n_2055),
.B(n_167),
.Y(n_2606)
);

BUFx2_ASAP7_75t_SL g2607 ( 
.A(n_2129),
.Y(n_2607)
);

AND2x4_ASAP7_75t_L g2608 ( 
.A(n_2164),
.B(n_166),
.Y(n_2608)
);

AND2x4_ASAP7_75t_L g2609 ( 
.A(n_2223),
.B(n_166),
.Y(n_2609)
);

INVx5_ASAP7_75t_L g2610 ( 
.A(n_2033),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_1978),
.Y(n_2611)
);

BUFx2_ASAP7_75t_L g2612 ( 
.A(n_2033),
.Y(n_2612)
);

AND2x4_ASAP7_75t_L g2613 ( 
.A(n_2032),
.B(n_167),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2113),
.Y(n_2614)
);

INVx3_ASAP7_75t_L g2615 ( 
.A(n_2113),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2049),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2080),
.B(n_168),
.Y(n_2617)
);

NOR2xp33_ASAP7_75t_SL g2618 ( 
.A(n_2252),
.B(n_789),
.Y(n_2618)
);

OR2x2_ASAP7_75t_L g2619 ( 
.A(n_2038),
.B(n_2048),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2053),
.Y(n_2620)
);

INVx1_ASAP7_75t_SL g2621 ( 
.A(n_2162),
.Y(n_2621)
);

BUFx6f_ASAP7_75t_L g2622 ( 
.A(n_2226),
.Y(n_2622)
);

AND2x4_ASAP7_75t_L g2623 ( 
.A(n_2073),
.B(n_168),
.Y(n_2623)
);

AND2x4_ASAP7_75t_L g2624 ( 
.A(n_2083),
.B(n_169),
.Y(n_2624)
);

OR2x6_ASAP7_75t_L g2625 ( 
.A(n_2268),
.B(n_169),
.Y(n_2625)
);

AND2x4_ASAP7_75t_L g2626 ( 
.A(n_2090),
.B(n_170),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2157),
.B(n_171),
.Y(n_2627)
);

BUFx6f_ASAP7_75t_L g2628 ( 
.A(n_2226),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2096),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2098),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2000),
.B(n_171),
.Y(n_2631)
);

INVx3_ASAP7_75t_L g2632 ( 
.A(n_2126),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2048),
.B(n_172),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2124),
.B(n_173),
.Y(n_2634)
);

BUFx2_ASAP7_75t_L g2635 ( 
.A(n_2061),
.Y(n_2635)
);

NOR2xp33_ASAP7_75t_L g2636 ( 
.A(n_2047),
.B(n_174),
.Y(n_2636)
);

AND2x4_ASAP7_75t_L g2637 ( 
.A(n_2101),
.B(n_174),
.Y(n_2637)
);

AND2x4_ASAP7_75t_L g2638 ( 
.A(n_2107),
.B(n_175),
.Y(n_2638)
);

AND2x4_ASAP7_75t_L g2639 ( 
.A(n_2112),
.B(n_176),
.Y(n_2639)
);

BUFx4f_ASAP7_75t_L g2640 ( 
.A(n_2061),
.Y(n_2640)
);

INVx1_ASAP7_75t_SL g2641 ( 
.A(n_2129),
.Y(n_2641)
);

INVx3_ASAP7_75t_L g2642 ( 
.A(n_2126),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2000),
.B(n_176),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2114),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2102),
.B(n_177),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2102),
.B(n_177),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2100),
.B(n_178),
.Y(n_2647)
);

AND2x4_ASAP7_75t_L g2648 ( 
.A(n_2118),
.B(n_179),
.Y(n_2648)
);

NAND2x1_ASAP7_75t_SL g2649 ( 
.A(n_2218),
.B(n_179),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2100),
.B(n_180),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2178),
.B(n_180),
.Y(n_2651)
);

INVxp67_ASAP7_75t_L g2652 ( 
.A(n_2250),
.Y(n_2652)
);

CKINVDCx20_ASAP7_75t_R g2653 ( 
.A(n_2210),
.Y(n_2653)
);

INVx3_ASAP7_75t_L g2654 ( 
.A(n_2189),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2174),
.B(n_181),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2121),
.Y(n_2656)
);

OR2x6_ASAP7_75t_L g2657 ( 
.A(n_2268),
.B(n_181),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2122),
.B(n_182),
.Y(n_2658)
);

BUFx12f_ASAP7_75t_L g2659 ( 
.A(n_1961),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2146),
.Y(n_2660)
);

INVx3_ASAP7_75t_L g2661 ( 
.A(n_2195),
.Y(n_2661)
);

AND2x4_ASAP7_75t_L g2662 ( 
.A(n_2153),
.B(n_182),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2154),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2171),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2176),
.B(n_183),
.Y(n_2665)
);

AND2x4_ASAP7_75t_L g2666 ( 
.A(n_2194),
.B(n_184),
.Y(n_2666)
);

INVx4_ASAP7_75t_L g2667 ( 
.A(n_2061),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2015),
.B(n_184),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_SL g2669 ( 
.A(n_2250),
.B(n_185),
.Y(n_2669)
);

BUFx2_ASAP7_75t_L g2670 ( 
.A(n_2061),
.Y(n_2670)
);

AND2x4_ASAP7_75t_L g2671 ( 
.A(n_2183),
.B(n_2180),
.Y(n_2671)
);

BUFx3_ASAP7_75t_L g2672 ( 
.A(n_2264),
.Y(n_2672)
);

BUFx6f_ASAP7_75t_L g2673 ( 
.A(n_2226),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2131),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2191),
.Y(n_2675)
);

AND2x4_ASAP7_75t_L g2676 ( 
.A(n_1961),
.B(n_185),
.Y(n_2676)
);

OR2x2_ASAP7_75t_L g2677 ( 
.A(n_2270),
.B(n_2015),
.Y(n_2677)
);

INVx3_ASAP7_75t_L g2678 ( 
.A(n_2105),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2191),
.Y(n_2679)
);

BUFx4f_ASAP7_75t_L g2680 ( 
.A(n_2105),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_SL g2681 ( 
.A(n_1970),
.B(n_186),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2115),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2092),
.B(n_186),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2092),
.B(n_187),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2157),
.B(n_187),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2017),
.B(n_188),
.Y(n_2686)
);

OR2x6_ASAP7_75t_L g2687 ( 
.A(n_2257),
.B(n_189),
.Y(n_2687)
);

AO21x2_ASAP7_75t_L g2688 ( 
.A1(n_2135),
.A2(n_791),
.B(n_790),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2160),
.B(n_189),
.Y(n_2689)
);

INVx8_ASAP7_75t_L g2690 ( 
.A(n_2131),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2012),
.Y(n_2691)
);

BUFx6f_ASAP7_75t_L g2692 ( 
.A(n_2071),
.Y(n_2692)
);

NOR2xp33_ASAP7_75t_L g2693 ( 
.A(n_2042),
.B(n_190),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2160),
.B(n_191),
.Y(n_2694)
);

INVx4_ASAP7_75t_L g2695 ( 
.A(n_2012),
.Y(n_2695)
);

BUFx3_ASAP7_75t_L g2696 ( 
.A(n_2017),
.Y(n_2696)
);

INVx3_ASAP7_75t_L g2697 ( 
.A(n_2050),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2050),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2184),
.Y(n_2699)
);

AND2x6_ASAP7_75t_L g2700 ( 
.A(n_2095),
.B(n_2104),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2161),
.B(n_192),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2115),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2074),
.B(n_192),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2074),
.B(n_193),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_1962),
.B(n_194),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2116),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_1962),
.B(n_194),
.Y(n_2707)
);

AND2x4_ASAP7_75t_L g2708 ( 
.A(n_1984),
.B(n_195),
.Y(n_2708)
);

AND2x4_ASAP7_75t_L g2709 ( 
.A(n_2224),
.B(n_196),
.Y(n_2709)
);

AO21x2_ASAP7_75t_L g2710 ( 
.A1(n_2135),
.A2(n_794),
.B(n_792),
.Y(n_2710)
);

INVx1_ASAP7_75t_SL g2711 ( 
.A(n_1970),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2270),
.B(n_197),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2116),
.Y(n_2713)
);

AND2x4_ASAP7_75t_L g2714 ( 
.A(n_2013),
.B(n_198),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_1996),
.B(n_199),
.Y(n_2715)
);

OR2x6_ASAP7_75t_L g2716 ( 
.A(n_2257),
.B(n_199),
.Y(n_2716)
);

CKINVDCx20_ASAP7_75t_R g2717 ( 
.A(n_1974),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2184),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2161),
.Y(n_2719)
);

BUFx2_ASAP7_75t_L g2720 ( 
.A(n_1974),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2166),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2166),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2184),
.Y(n_2723)
);

INVx4_ASAP7_75t_L g2724 ( 
.A(n_2106),
.Y(n_2724)
);

NOR2xp33_ASAP7_75t_L g2725 ( 
.A(n_1980),
.B(n_1988),
.Y(n_2725)
);

NAND2x1p5_ASAP7_75t_L g2726 ( 
.A(n_2283),
.B(n_201),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2167),
.Y(n_2727)
);

AND2x4_ASAP7_75t_L g2728 ( 
.A(n_2013),
.B(n_200),
.Y(n_2728)
);

AND2x4_ASAP7_75t_L g2729 ( 
.A(n_2167),
.B(n_200),
.Y(n_2729)
);

INVx3_ASAP7_75t_L g2730 ( 
.A(n_2120),
.Y(n_2730)
);

BUFx4_ASAP7_75t_SL g2731 ( 
.A(n_2245),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2231),
.B(n_201),
.Y(n_2732)
);

BUFx5_ASAP7_75t_L g2733 ( 
.A(n_2263),
.Y(n_2733)
);

AND2x2_ASAP7_75t_L g2734 ( 
.A(n_1996),
.B(n_2190),
.Y(n_2734)
);

AND2x4_ASAP7_75t_L g2735 ( 
.A(n_2066),
.B(n_202),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2197),
.B(n_202),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2231),
.B(n_203),
.Y(n_2737)
);

BUFx2_ASAP7_75t_L g2738 ( 
.A(n_1980),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2193),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2193),
.Y(n_2740)
);

OR2x6_ASAP7_75t_L g2741 ( 
.A(n_2240),
.B(n_203),
.Y(n_2741)
);

OR2x2_ASAP7_75t_L g2742 ( 
.A(n_1988),
.B(n_204),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2259),
.B(n_204),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2066),
.B(n_205),
.Y(n_2744)
);

OR2x2_ASAP7_75t_L g2745 ( 
.A(n_2212),
.B(n_206),
.Y(n_2745)
);

NOR2xp67_ASAP7_75t_L g2746 ( 
.A(n_2199),
.B(n_795),
.Y(n_2746)
);

AND2x4_ASAP7_75t_L g2747 ( 
.A(n_2230),
.B(n_2237),
.Y(n_2747)
);

NOR2xp33_ASAP7_75t_SL g2748 ( 
.A(n_2145),
.B(n_796),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2199),
.Y(n_2749)
);

BUFx4f_ASAP7_75t_L g2750 ( 
.A(n_2236),
.Y(n_2750)
);

BUFx3_ASAP7_75t_L g2751 ( 
.A(n_2230),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2237),
.B(n_206),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2205),
.B(n_2152),
.Y(n_2753)
);

BUFx2_ASAP7_75t_L g2754 ( 
.A(n_2205),
.Y(n_2754)
);

INVx4_ASAP7_75t_L g2755 ( 
.A(n_2236),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2111),
.B(n_208),
.Y(n_2756)
);

BUFx2_ASAP7_75t_L g2757 ( 
.A(n_2145),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2203),
.Y(n_2758)
);

NAND2x1p5_ASAP7_75t_L g2759 ( 
.A(n_2236),
.B(n_211),
.Y(n_2759)
);

INVx3_ASAP7_75t_L g2760 ( 
.A(n_2266),
.Y(n_2760)
);

NOR2x1_ASAP7_75t_L g2761 ( 
.A(n_2152),
.B(n_209),
.Y(n_2761)
);

BUFx3_ASAP7_75t_L g2762 ( 
.A(n_2111),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2262),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_1960),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_1960),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2244),
.B(n_209),
.Y(n_2766)
);

NOR2x1_ASAP7_75t_L g2767 ( 
.A(n_2244),
.B(n_211),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_1972),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_1972),
.Y(n_2769)
);

AND2x4_ASAP7_75t_L g2770 ( 
.A(n_1957),
.B(n_212),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2136),
.Y(n_2771)
);

BUFx8_ASAP7_75t_L g2772 ( 
.A(n_2099),
.Y(n_2772)
);

BUFx4f_ASAP7_75t_L g2773 ( 
.A(n_2279),
.Y(n_2773)
);

INVx4_ASAP7_75t_L g2774 ( 
.A(n_1976),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_1972),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2136),
.Y(n_2776)
);

AND2x4_ASAP7_75t_L g2777 ( 
.A(n_1957),
.B(n_212),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_1958),
.B(n_213),
.Y(n_2778)
);

NAND2x1_ASAP7_75t_SL g2779 ( 
.A(n_2287),
.B(n_213),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_1958),
.B(n_214),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_1958),
.B(n_214),
.Y(n_2781)
);

AND2x4_ASAP7_75t_L g2782 ( 
.A(n_1957),
.B(n_215),
.Y(n_2782)
);

INVx8_ASAP7_75t_L g2783 ( 
.A(n_1976),
.Y(n_2783)
);

BUFx3_ASAP7_75t_L g2784 ( 
.A(n_2275),
.Y(n_2784)
);

CKINVDCx6p67_ASAP7_75t_R g2785 ( 
.A(n_2099),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_1958),
.B(n_216),
.Y(n_2786)
);

INVx3_ASAP7_75t_L g2787 ( 
.A(n_1976),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_1972),
.B(n_216),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_1958),
.B(n_217),
.Y(n_2789)
);

AND2x4_ASAP7_75t_L g2790 ( 
.A(n_1957),
.B(n_217),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_1958),
.B(n_218),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_1958),
.B(n_218),
.Y(n_2792)
);

NOR2xp33_ASAP7_75t_L g2793 ( 
.A(n_2062),
.B(n_219),
.Y(n_2793)
);

INVx3_ASAP7_75t_L g2794 ( 
.A(n_1976),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_1958),
.B(n_221),
.Y(n_2795)
);

NOR2xp67_ASAP7_75t_L g2796 ( 
.A(n_2252),
.B(n_797),
.Y(n_2796)
);

INVx4_ASAP7_75t_L g2797 ( 
.A(n_1976),
.Y(n_2797)
);

BUFx6f_ASAP7_75t_L g2798 ( 
.A(n_1976),
.Y(n_2798)
);

BUFx3_ASAP7_75t_L g2799 ( 
.A(n_2275),
.Y(n_2799)
);

AND2x2_ASAP7_75t_L g2800 ( 
.A(n_1958),
.B(n_221),
.Y(n_2800)
);

BUFx12f_ASAP7_75t_L g2801 ( 
.A(n_2772),
.Y(n_2801)
);

BUFx3_ASAP7_75t_L g2802 ( 
.A(n_2772),
.Y(n_2802)
);

INVxp67_ASAP7_75t_SL g2803 ( 
.A(n_2313),
.Y(n_2803)
);

BUFx2_ASAP7_75t_L g2804 ( 
.A(n_2583),
.Y(n_2804)
);

INVx4_ASAP7_75t_L g2805 ( 
.A(n_2502),
.Y(n_2805)
);

NAND2x1p5_ASAP7_75t_L g2806 ( 
.A(n_2680),
.B(n_222),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2327),
.Y(n_2807)
);

CKINVDCx11_ASAP7_75t_R g2808 ( 
.A(n_2306),
.Y(n_2808)
);

INVx3_ASAP7_75t_L g2809 ( 
.A(n_2680),
.Y(n_2809)
);

BUFx3_ASAP7_75t_L g2810 ( 
.A(n_2316),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_2416),
.Y(n_2811)
);

BUFx6f_ASAP7_75t_L g2812 ( 
.A(n_2319),
.Y(n_2812)
);

AOI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_2735),
.A2(n_226),
.B1(n_223),
.B2(n_225),
.Y(n_2813)
);

BUFx12f_ASAP7_75t_L g2814 ( 
.A(n_2338),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2313),
.Y(n_2815)
);

INVx4_ASAP7_75t_L g2816 ( 
.A(n_2785),
.Y(n_2816)
);

AND2x4_ASAP7_75t_L g2817 ( 
.A(n_2322),
.B(n_227),
.Y(n_2817)
);

INVxp67_ASAP7_75t_SL g2818 ( 
.A(n_2322),
.Y(n_2818)
);

BUFx12f_ASAP7_75t_L g2819 ( 
.A(n_2393),
.Y(n_2819)
);

INVx3_ASAP7_75t_SL g2820 ( 
.A(n_2303),
.Y(n_2820)
);

INVx1_ASAP7_75t_SL g2821 ( 
.A(n_2487),
.Y(n_2821)
);

BUFx3_ASAP7_75t_L g2822 ( 
.A(n_2784),
.Y(n_2822)
);

INVx1_ASAP7_75t_SL g2823 ( 
.A(n_2487),
.Y(n_2823)
);

INVx4_ASAP7_75t_L g2824 ( 
.A(n_2783),
.Y(n_2824)
);

AOI22xp33_ASAP7_75t_L g2825 ( 
.A1(n_2458),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.Y(n_2825)
);

INVx6_ASAP7_75t_SL g2826 ( 
.A(n_2303),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2682),
.B(n_228),
.Y(n_2827)
);

INVx4_ASAP7_75t_L g2828 ( 
.A(n_2783),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2682),
.B(n_230),
.Y(n_2829)
);

NAND2x1p5_ASAP7_75t_L g2830 ( 
.A(n_2640),
.B(n_2535),
.Y(n_2830)
);

NAND2x1p5_ASAP7_75t_L g2831 ( 
.A(n_2640),
.B(n_230),
.Y(n_2831)
);

INVxp67_ASAP7_75t_SL g2832 ( 
.A(n_2735),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2327),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2465),
.B(n_231),
.Y(n_2834)
);

AOI22xp33_ASAP7_75t_L g2835 ( 
.A1(n_2330),
.A2(n_235),
.B1(n_232),
.B2(n_233),
.Y(n_2835)
);

CKINVDCx16_ASAP7_75t_R g2836 ( 
.A(n_2335),
.Y(n_2836)
);

INVx5_ASAP7_75t_SL g2837 ( 
.A(n_2310),
.Y(n_2837)
);

CKINVDCx5p33_ASAP7_75t_R g2838 ( 
.A(n_2540),
.Y(n_2838)
);

NAND2x1p5_ASAP7_75t_L g2839 ( 
.A(n_2535),
.B(n_232),
.Y(n_2839)
);

NOR2xp33_ASAP7_75t_L g2840 ( 
.A(n_2619),
.B(n_233),
.Y(n_2840)
);

AOI22xp33_ASAP7_75t_L g2841 ( 
.A1(n_2330),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2702),
.B(n_237),
.Y(n_2842)
);

BUFx6f_ASAP7_75t_L g2843 ( 
.A(n_2319),
.Y(n_2843)
);

BUFx3_ASAP7_75t_L g2844 ( 
.A(n_2799),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2304),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2297),
.Y(n_2846)
);

BUFx6f_ASAP7_75t_L g2847 ( 
.A(n_2319),
.Y(n_2847)
);

BUFx2_ASAP7_75t_R g2848 ( 
.A(n_2555),
.Y(n_2848)
);

BUFx3_ASAP7_75t_L g2849 ( 
.A(n_2344),
.Y(n_2849)
);

BUFx3_ASAP7_75t_L g2850 ( 
.A(n_2374),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2304),
.Y(n_2851)
);

BUFx2_ASAP7_75t_SL g2852 ( 
.A(n_2365),
.Y(n_2852)
);

CKINVDCx5p33_ASAP7_75t_R g2853 ( 
.A(n_2468),
.Y(n_2853)
);

INVxp67_ASAP7_75t_SL g2854 ( 
.A(n_2714),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2300),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2771),
.Y(n_2856)
);

INVxp67_ASAP7_75t_SL g2857 ( 
.A(n_2714),
.Y(n_2857)
);

INVx5_ASAP7_75t_L g2858 ( 
.A(n_2783),
.Y(n_2858)
);

OR2x2_ASAP7_75t_L g2859 ( 
.A(n_2342),
.B(n_238),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2702),
.B(n_239),
.Y(n_2860)
);

INVx1_ASAP7_75t_SL g2861 ( 
.A(n_2557),
.Y(n_2861)
);

CKINVDCx20_ASAP7_75t_R g2862 ( 
.A(n_2468),
.Y(n_2862)
);

BUFx3_ASAP7_75t_L g2863 ( 
.A(n_2365),
.Y(n_2863)
);

BUFx3_ASAP7_75t_L g2864 ( 
.A(n_2365),
.Y(n_2864)
);

INVx5_ASAP7_75t_SL g2865 ( 
.A(n_2310),
.Y(n_2865)
);

AND2x2_ASAP7_75t_L g2866 ( 
.A(n_2366),
.B(n_239),
.Y(n_2866)
);

CKINVDCx5p33_ASAP7_75t_R g2867 ( 
.A(n_2460),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2768),
.Y(n_2868)
);

INVx2_ASAP7_75t_SL g2869 ( 
.A(n_2539),
.Y(n_2869)
);

INVx5_ASAP7_75t_L g2870 ( 
.A(n_2415),
.Y(n_2870)
);

INVx4_ASAP7_75t_L g2871 ( 
.A(n_2539),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2706),
.B(n_2713),
.Y(n_2872)
);

BUFx6f_ASAP7_75t_L g2873 ( 
.A(n_2315),
.Y(n_2873)
);

CKINVDCx16_ASAP7_75t_R g2874 ( 
.A(n_2659),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2776),
.Y(n_2875)
);

BUFx2_ASAP7_75t_L g2876 ( 
.A(n_2358),
.Y(n_2876)
);

INVx3_ASAP7_75t_L g2877 ( 
.A(n_2750),
.Y(n_2877)
);

NAND2x1p5_ASAP7_75t_L g2878 ( 
.A(n_2470),
.B(n_2610),
.Y(n_2878)
);

INVx3_ASAP7_75t_L g2879 ( 
.A(n_2750),
.Y(n_2879)
);

INVxp67_ASAP7_75t_L g2880 ( 
.A(n_2357),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2597),
.B(n_240),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2706),
.B(n_240),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2373),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2768),
.Y(n_2884)
);

BUFx3_ASAP7_75t_L g2885 ( 
.A(n_2476),
.Y(n_2885)
);

BUFx12f_ASAP7_75t_L g2886 ( 
.A(n_2337),
.Y(n_2886)
);

BUFx2_ASAP7_75t_L g2887 ( 
.A(n_2360),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2389),
.Y(n_2888)
);

OR2x2_ASAP7_75t_L g2889 ( 
.A(n_2479),
.B(n_2483),
.Y(n_2889)
);

BUFx2_ASAP7_75t_L g2890 ( 
.A(n_2415),
.Y(n_2890)
);

NOR2xp33_ASAP7_75t_L g2891 ( 
.A(n_2511),
.B(n_241),
.Y(n_2891)
);

BUFx3_ASAP7_75t_L g2892 ( 
.A(n_2417),
.Y(n_2892)
);

INVx6_ASAP7_75t_SL g2893 ( 
.A(n_2337),
.Y(n_2893)
);

BUFx3_ASAP7_75t_L g2894 ( 
.A(n_2394),
.Y(n_2894)
);

BUFx3_ASAP7_75t_L g2895 ( 
.A(n_2424),
.Y(n_2895)
);

INVx2_ASAP7_75t_SL g2896 ( 
.A(n_2525),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2492),
.B(n_2505),
.Y(n_2897)
);

BUFx12f_ASAP7_75t_L g2898 ( 
.A(n_2530),
.Y(n_2898)
);

BUFx3_ASAP7_75t_L g2899 ( 
.A(n_2504),
.Y(n_2899)
);

INVx1_ASAP7_75t_SL g2900 ( 
.A(n_2557),
.Y(n_2900)
);

INVx4_ASAP7_75t_L g2901 ( 
.A(n_2328),
.Y(n_2901)
);

NAND2x1p5_ASAP7_75t_L g2902 ( 
.A(n_2470),
.B(n_242),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2392),
.Y(n_2903)
);

BUFx4f_ASAP7_75t_SL g2904 ( 
.A(n_2653),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2773),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2769),
.Y(n_2906)
);

OAI22xp5_ASAP7_75t_L g2907 ( 
.A1(n_2728),
.A2(n_246),
.B1(n_243),
.B2(n_244),
.Y(n_2907)
);

BUFx2_ASAP7_75t_L g2908 ( 
.A(n_2328),
.Y(n_2908)
);

INVxp67_ASAP7_75t_SL g2909 ( 
.A(n_2728),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2419),
.Y(n_2910)
);

AND2x2_ASAP7_75t_L g2911 ( 
.A(n_2516),
.B(n_2510),
.Y(n_2911)
);

INVx1_ASAP7_75t_SL g2912 ( 
.A(n_2621),
.Y(n_2912)
);

BUFx4_ASAP7_75t_SL g2913 ( 
.A(n_2530),
.Y(n_2913)
);

BUFx3_ASAP7_75t_L g2914 ( 
.A(n_2339),
.Y(n_2914)
);

AND2x2_ASAP7_75t_L g2915 ( 
.A(n_2560),
.B(n_246),
.Y(n_2915)
);

INVx2_ASAP7_75t_SL g2916 ( 
.A(n_2525),
.Y(n_2916)
);

BUFx2_ASAP7_75t_L g2917 ( 
.A(n_2328),
.Y(n_2917)
);

INVx2_ASAP7_75t_SL g2918 ( 
.A(n_2432),
.Y(n_2918)
);

INVx4_ASAP7_75t_L g2919 ( 
.A(n_2328),
.Y(n_2919)
);

INVx2_ASAP7_75t_SL g2920 ( 
.A(n_2690),
.Y(n_2920)
);

AND2x2_ASAP7_75t_L g2921 ( 
.A(n_2676),
.B(n_247),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2440),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2769),
.Y(n_2923)
);

BUFx2_ASAP7_75t_SL g2924 ( 
.A(n_2490),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2775),
.Y(n_2925)
);

BUFx6f_ASAP7_75t_L g2926 ( 
.A(n_2315),
.Y(n_2926)
);

CKINVDCx16_ASAP7_75t_R g2927 ( 
.A(n_2545),
.Y(n_2927)
);

BUFx2_ASAP7_75t_SL g2928 ( 
.A(n_2400),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2775),
.Y(n_2929)
);

HB1xp67_ASAP7_75t_L g2930 ( 
.A(n_2352),
.Y(n_2930)
);

BUFx3_ASAP7_75t_L g2931 ( 
.A(n_2339),
.Y(n_2931)
);

OR2x6_ASAP7_75t_L g2932 ( 
.A(n_2469),
.B(n_248),
.Y(n_2932)
);

BUFx2_ASAP7_75t_L g2933 ( 
.A(n_2400),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2353),
.Y(n_2934)
);

BUFx5_ASAP7_75t_L g2935 ( 
.A(n_2700),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2353),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2713),
.B(n_249),
.Y(n_2937)
);

BUFx12f_ASAP7_75t_L g2938 ( 
.A(n_2545),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2371),
.Y(n_2939)
);

BUFx2_ASAP7_75t_SL g2940 ( 
.A(n_2400),
.Y(n_2940)
);

INVx1_ASAP7_75t_SL g2941 ( 
.A(n_2621),
.Y(n_2941)
);

INVx5_ASAP7_75t_L g2942 ( 
.A(n_2315),
.Y(n_2942)
);

BUFx3_ASAP7_75t_L g2943 ( 
.A(n_2339),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_SL g2944 ( 
.A(n_2325),
.B(n_799),
.Y(n_2944)
);

INVx1_ASAP7_75t_SL g2945 ( 
.A(n_2607),
.Y(n_2945)
);

NAND2x1p5_ASAP7_75t_L g2946 ( 
.A(n_2470),
.B(n_251),
.Y(n_2946)
);

BUFx3_ASAP7_75t_L g2947 ( 
.A(n_2430),
.Y(n_2947)
);

INVx2_ASAP7_75t_SL g2948 ( 
.A(n_2690),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2676),
.B(n_251),
.Y(n_2949)
);

INVx5_ASAP7_75t_L g2950 ( 
.A(n_2798),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2449),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2719),
.B(n_2721),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2371),
.Y(n_2953)
);

BUFx2_ASAP7_75t_L g2954 ( 
.A(n_2400),
.Y(n_2954)
);

BUFx3_ASAP7_75t_L g2955 ( 
.A(n_2430),
.Y(n_2955)
);

BUFx2_ASAP7_75t_L g2956 ( 
.A(n_2520),
.Y(n_2956)
);

BUFx12f_ASAP7_75t_L g2957 ( 
.A(n_2578),
.Y(n_2957)
);

BUFx3_ASAP7_75t_L g2958 ( 
.A(n_2696),
.Y(n_2958)
);

BUFx12f_ASAP7_75t_L g2959 ( 
.A(n_2573),
.Y(n_2959)
);

BUFx6f_ASAP7_75t_SL g2960 ( 
.A(n_2573),
.Y(n_2960)
);

BUFx2_ASAP7_75t_L g2961 ( 
.A(n_2520),
.Y(n_2961)
);

INVx4_ASAP7_75t_L g2962 ( 
.A(n_2509),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2375),
.Y(n_2963)
);

OR2x2_ASAP7_75t_L g2964 ( 
.A(n_2345),
.B(n_252),
.Y(n_2964)
);

INVx6_ASAP7_75t_SL g2965 ( 
.A(n_2509),
.Y(n_2965)
);

BUFx6f_ASAP7_75t_SL g2966 ( 
.A(n_2687),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2375),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2355),
.B(n_252),
.Y(n_2968)
);

INVx3_ASAP7_75t_SL g2969 ( 
.A(n_2687),
.Y(n_2969)
);

INVx8_ASAP7_75t_L g2970 ( 
.A(n_2690),
.Y(n_2970)
);

AND2x2_ASAP7_75t_L g2971 ( 
.A(n_2425),
.B(n_253),
.Y(n_2971)
);

BUFx2_ASAP7_75t_L g2972 ( 
.A(n_2551),
.Y(n_2972)
);

INVx1_ASAP7_75t_SL g2973 ( 
.A(n_2352),
.Y(n_2973)
);

BUFx3_ASAP7_75t_L g2974 ( 
.A(n_2480),
.Y(n_2974)
);

BUFx6f_ASAP7_75t_L g2975 ( 
.A(n_2798),
.Y(n_2975)
);

INVx1_ASAP7_75t_SL g2976 ( 
.A(n_2354),
.Y(n_2976)
);

AND2x2_ASAP7_75t_L g2977 ( 
.A(n_2431),
.B(n_2603),
.Y(n_2977)
);

BUFx6f_ASAP7_75t_L g2978 ( 
.A(n_2798),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2719),
.B(n_255),
.Y(n_2979)
);

INVx8_ASAP7_75t_L g2980 ( 
.A(n_2716),
.Y(n_2980)
);

INVx5_ASAP7_75t_L g2981 ( 
.A(n_2544),
.Y(n_2981)
);

INVx1_ASAP7_75t_SL g2982 ( 
.A(n_2354),
.Y(n_2982)
);

INVx4_ASAP7_75t_L g2983 ( 
.A(n_2610),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2333),
.Y(n_2984)
);

BUFx3_ASAP7_75t_L g2985 ( 
.A(n_2567),
.Y(n_2985)
);

INVx1_ASAP7_75t_SL g2986 ( 
.A(n_2563),
.Y(n_2986)
);

BUFx6f_ASAP7_75t_L g2987 ( 
.A(n_2369),
.Y(n_2987)
);

AND2x2_ASAP7_75t_L g2988 ( 
.A(n_2631),
.B(n_256),
.Y(n_2988)
);

AND2x4_ASAP7_75t_L g2989 ( 
.A(n_2544),
.B(n_259),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2721),
.B(n_259),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2485),
.Y(n_2991)
);

BUFx2_ASAP7_75t_L g2992 ( 
.A(n_2755),
.Y(n_2992)
);

INVx8_ASAP7_75t_L g2993 ( 
.A(n_2716),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2489),
.Y(n_2994)
);

BUFx3_ASAP7_75t_L g2995 ( 
.A(n_2580),
.Y(n_2995)
);

BUFx3_ASAP7_75t_L g2996 ( 
.A(n_2314),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2534),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2553),
.Y(n_2998)
);

INVx5_ASAP7_75t_L g2999 ( 
.A(n_2369),
.Y(n_2999)
);

CKINVDCx16_ASAP7_75t_R g3000 ( 
.A(n_2717),
.Y(n_3000)
);

BUFx2_ASAP7_75t_SL g3001 ( 
.A(n_2610),
.Y(n_3001)
);

BUFx2_ASAP7_75t_L g3002 ( 
.A(n_2755),
.Y(n_3002)
);

BUFx6f_ASAP7_75t_L g3003 ( 
.A(n_2369),
.Y(n_3003)
);

CKINVDCx20_ASAP7_75t_R g3004 ( 
.A(n_2773),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2333),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2788),
.Y(n_3006)
);

BUFx6f_ASAP7_75t_L g3007 ( 
.A(n_2387),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2788),
.Y(n_3008)
);

BUFx3_ASAP7_75t_L g3009 ( 
.A(n_2314),
.Y(n_3009)
);

BUFx2_ASAP7_75t_L g3010 ( 
.A(n_2402),
.Y(n_3010)
);

INVx8_ASAP7_75t_L g3011 ( 
.A(n_2515),
.Y(n_3011)
);

BUFx6f_ASAP7_75t_L g3012 ( 
.A(n_2387),
.Y(n_3012)
);

BUFx3_ASAP7_75t_L g3013 ( 
.A(n_2550),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2349),
.Y(n_3014)
);

NAND2x1p5_ASAP7_75t_L g3015 ( 
.A(n_2596),
.B(n_260),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2349),
.Y(n_3016)
);

AOI22xp33_ASAP7_75t_L g3017 ( 
.A1(n_2722),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_3017)
);

BUFx3_ASAP7_75t_L g3018 ( 
.A(n_2550),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2616),
.Y(n_3019)
);

AND2x2_ASAP7_75t_L g3020 ( 
.A(n_2643),
.B(n_262),
.Y(n_3020)
);

CKINVDCx6p67_ASAP7_75t_R g3021 ( 
.A(n_2625),
.Y(n_3021)
);

BUFx3_ASAP7_75t_L g3022 ( 
.A(n_2356),
.Y(n_3022)
);

CKINVDCx6p67_ASAP7_75t_R g3023 ( 
.A(n_2625),
.Y(n_3023)
);

INVx1_ASAP7_75t_SL g3024 ( 
.A(n_2563),
.Y(n_3024)
);

BUFx4f_ASAP7_75t_L g3025 ( 
.A(n_2307),
.Y(n_3025)
);

BUFx3_ASAP7_75t_L g3026 ( 
.A(n_2356),
.Y(n_3026)
);

BUFx12f_ASAP7_75t_L g3027 ( 
.A(n_2311),
.Y(n_3027)
);

INVx5_ASAP7_75t_L g3028 ( 
.A(n_2596),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2722),
.B(n_263),
.Y(n_3029)
);

INVx2_ASAP7_75t_SL g3030 ( 
.A(n_2350),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2436),
.Y(n_3031)
);

INVx5_ASAP7_75t_L g3032 ( 
.A(n_2667),
.Y(n_3032)
);

INVx1_ASAP7_75t_SL g3033 ( 
.A(n_2570),
.Y(n_3033)
);

NAND2x1p5_ASAP7_75t_L g3034 ( 
.A(n_2667),
.B(n_263),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2436),
.Y(n_3035)
);

BUFx2_ASAP7_75t_R g3036 ( 
.A(n_2576),
.Y(n_3036)
);

AOI22xp33_ASAP7_75t_L g3037 ( 
.A1(n_2727),
.A2(n_2747),
.B1(n_2679),
.B2(n_2675),
.Y(n_3037)
);

BUFx12f_ASAP7_75t_L g3038 ( 
.A(n_2447),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2620),
.Y(n_3039)
);

BUFx6f_ASAP7_75t_L g3040 ( 
.A(n_2387),
.Y(n_3040)
);

INVx8_ASAP7_75t_L g3041 ( 
.A(n_2515),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2629),
.Y(n_3042)
);

BUFx2_ASAP7_75t_R g3043 ( 
.A(n_2372),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_2668),
.B(n_264),
.Y(n_3044)
);

INVx3_ASAP7_75t_L g3045 ( 
.A(n_2326),
.Y(n_3045)
);

CKINVDCx5p33_ASAP7_75t_R g3046 ( 
.A(n_2731),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2663),
.Y(n_3047)
);

BUFx3_ASAP7_75t_L g3048 ( 
.A(n_2422),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2301),
.Y(n_3049)
);

BUFx2_ASAP7_75t_L g3050 ( 
.A(n_2350),
.Y(n_3050)
);

CKINVDCx12_ASAP7_75t_R g3051 ( 
.A(n_2657),
.Y(n_3051)
);

BUFx6f_ASAP7_75t_L g3052 ( 
.A(n_2411),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2308),
.Y(n_3053)
);

BUFx3_ASAP7_75t_L g3054 ( 
.A(n_2422),
.Y(n_3054)
);

INVx2_ASAP7_75t_SL g3055 ( 
.A(n_2570),
.Y(n_3055)
);

BUFx12f_ASAP7_75t_L g3056 ( 
.A(n_2526),
.Y(n_3056)
);

BUFx2_ASAP7_75t_R g3057 ( 
.A(n_2669),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2686),
.B(n_264),
.Y(n_3058)
);

INVx3_ASAP7_75t_L g3059 ( 
.A(n_2326),
.Y(n_3059)
);

BUFx2_ASAP7_75t_L g3060 ( 
.A(n_2448),
.Y(n_3060)
);

CKINVDCx5p33_ASAP7_75t_R g3061 ( 
.A(n_2657),
.Y(n_3061)
);

INVx3_ASAP7_75t_L g3062 ( 
.A(n_2774),
.Y(n_3062)
);

INVx6_ASAP7_75t_SL g3063 ( 
.A(n_2526),
.Y(n_3063)
);

AND2x4_ASAP7_75t_L g3064 ( 
.A(n_2406),
.B(n_265),
.Y(n_3064)
);

CKINVDCx20_ASAP7_75t_R g3065 ( 
.A(n_2336),
.Y(n_3065)
);

INVx3_ASAP7_75t_L g3066 ( 
.A(n_2774),
.Y(n_3066)
);

BUFx3_ASAP7_75t_L g3067 ( 
.A(n_2455),
.Y(n_3067)
);

CKINVDCx5p33_ASAP7_75t_R g3068 ( 
.A(n_2741),
.Y(n_3068)
);

INVx1_ASAP7_75t_SL g3069 ( 
.A(n_2641),
.Y(n_3069)
);

BUFx3_ASAP7_75t_L g3070 ( 
.A(n_2427),
.Y(n_3070)
);

INVx2_ASAP7_75t_SL g3071 ( 
.A(n_2448),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2517),
.Y(n_3072)
);

NOR2xp33_ASAP7_75t_L g3073 ( 
.A(n_2652),
.B(n_265),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2318),
.Y(n_3074)
);

CKINVDCx5p33_ASAP7_75t_R g3075 ( 
.A(n_2741),
.Y(n_3075)
);

HB1xp67_ASAP7_75t_L g3076 ( 
.A(n_2493),
.Y(n_3076)
);

BUFx2_ASAP7_75t_SL g3077 ( 
.A(n_2406),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2727),
.B(n_266),
.Y(n_3078)
);

BUFx2_ASAP7_75t_SL g3079 ( 
.A(n_2406),
.Y(n_3079)
);

BUFx2_ASAP7_75t_L g3080 ( 
.A(n_2457),
.Y(n_3080)
);

CKINVDCx5p33_ASAP7_75t_R g3081 ( 
.A(n_2672),
.Y(n_3081)
);

BUFx3_ASAP7_75t_L g3082 ( 
.A(n_2427),
.Y(n_3082)
);

AO21x2_ASAP7_75t_L g3083 ( 
.A1(n_2758),
.A2(n_806),
.B(n_800),
.Y(n_3083)
);

BUFx3_ASAP7_75t_L g3084 ( 
.A(n_2368),
.Y(n_3084)
);

INVx2_ASAP7_75t_SL g3085 ( 
.A(n_2457),
.Y(n_3085)
);

INVx5_ASAP7_75t_L g3086 ( 
.A(n_2411),
.Y(n_3086)
);

INVx2_ASAP7_75t_SL g3087 ( 
.A(n_2462),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2517),
.Y(n_3088)
);

NOR2xp33_ASAP7_75t_L g3089 ( 
.A(n_2677),
.B(n_266),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2521),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2564),
.Y(n_3091)
);

BUFx4f_ASAP7_75t_SL g3092 ( 
.A(n_2797),
.Y(n_3092)
);

INVx2_ASAP7_75t_SL g3093 ( 
.A(n_2462),
.Y(n_3093)
);

INVx5_ASAP7_75t_L g3094 ( 
.A(n_2411),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2568),
.Y(n_3095)
);

INVx5_ASAP7_75t_L g3096 ( 
.A(n_2428),
.Y(n_3096)
);

BUFx3_ASAP7_75t_L g3097 ( 
.A(n_2382),
.Y(n_3097)
);

INVx2_ASAP7_75t_SL g3098 ( 
.A(n_2472),
.Y(n_3098)
);

BUFx4_ASAP7_75t_SL g3099 ( 
.A(n_2552),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2739),
.B(n_267),
.Y(n_3100)
);

BUFx4f_ASAP7_75t_L g3101 ( 
.A(n_2577),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_2703),
.B(n_267),
.Y(n_3102)
);

INVx6_ASAP7_75t_L g3103 ( 
.A(n_2708),
.Y(n_3103)
);

INVx5_ASAP7_75t_L g3104 ( 
.A(n_2428),
.Y(n_3104)
);

NAND2x1p5_ASAP7_75t_L g3105 ( 
.A(n_2678),
.B(n_268),
.Y(n_3105)
);

BUFx6f_ASAP7_75t_L g3106 ( 
.A(n_2428),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2521),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2532),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2532),
.Y(n_3109)
);

NAND2x1p5_ASAP7_75t_L g3110 ( 
.A(n_2678),
.B(n_268),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2537),
.Y(n_3111)
);

INVx1_ASAP7_75t_SL g3112 ( 
.A(n_2641),
.Y(n_3112)
);

INVx3_ASAP7_75t_L g3113 ( 
.A(n_2797),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2537),
.Y(n_3114)
);

BUFx12f_ASAP7_75t_L g3115 ( 
.A(n_2390),
.Y(n_3115)
);

BUFx4f_ASAP7_75t_SL g3116 ( 
.A(n_2472),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2543),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_2704),
.B(n_269),
.Y(n_3118)
);

INVx1_ASAP7_75t_SL g3119 ( 
.A(n_2445),
.Y(n_3119)
);

CKINVDCx20_ASAP7_75t_R g3120 ( 
.A(n_2446),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_2414),
.B(n_269),
.Y(n_3121)
);

BUFx6f_ASAP7_75t_L g3122 ( 
.A(n_2445),
.Y(n_3122)
);

BUFx12f_ASAP7_75t_L g3123 ( 
.A(n_2390),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_2543),
.Y(n_3124)
);

NAND2x1p5_ASAP7_75t_L g3125 ( 
.A(n_2581),
.B(n_270),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2582),
.Y(n_3126)
);

INVx3_ASAP7_75t_SL g3127 ( 
.A(n_2613),
.Y(n_3127)
);

BUFx6f_ASAP7_75t_L g3128 ( 
.A(n_2445),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2582),
.Y(n_3129)
);

NAND2x1p5_ASAP7_75t_L g3130 ( 
.A(n_2602),
.B(n_270),
.Y(n_3130)
);

INVx3_ASAP7_75t_L g3131 ( 
.A(n_2695),
.Y(n_3131)
);

BUFx2_ASAP7_75t_L g3132 ( 
.A(n_2493),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2586),
.Y(n_3133)
);

BUFx3_ASAP7_75t_L g3134 ( 
.A(n_2398),
.Y(n_3134)
);

INVx1_ASAP7_75t_SL g3135 ( 
.A(n_2558),
.Y(n_3135)
);

OR2x2_ASAP7_75t_L g3136 ( 
.A(n_2592),
.B(n_272),
.Y(n_3136)
);

BUFx3_ASAP7_75t_L g3137 ( 
.A(n_2398),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2586),
.Y(n_3138)
);

BUFx12f_ASAP7_75t_L g3139 ( 
.A(n_2395),
.Y(n_3139)
);

INVx2_ASAP7_75t_SL g3140 ( 
.A(n_2666),
.Y(n_3140)
);

BUFx5_ASAP7_75t_L g3141 ( 
.A(n_2700),
.Y(n_3141)
);

INVx3_ASAP7_75t_L g3142 ( 
.A(n_2695),
.Y(n_3142)
);

BUFx12f_ASAP7_75t_L g3143 ( 
.A(n_2395),
.Y(n_3143)
);

BUFx3_ASAP7_75t_L g3144 ( 
.A(n_2405),
.Y(n_3144)
);

BUFx2_ASAP7_75t_SL g3145 ( 
.A(n_2613),
.Y(n_3145)
);

BUFx6f_ASAP7_75t_SL g3146 ( 
.A(n_2623),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2630),
.Y(n_3147)
);

INVx3_ASAP7_75t_L g3148 ( 
.A(n_2632),
.Y(n_3148)
);

INVx2_ASAP7_75t_SL g3149 ( 
.A(n_2666),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2630),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2644),
.Y(n_3151)
);

BUFx2_ASAP7_75t_L g3152 ( 
.A(n_2405),
.Y(n_3152)
);

BUFx6f_ASAP7_75t_SL g3153 ( 
.A(n_2623),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2644),
.Y(n_3154)
);

BUFx6f_ASAP7_75t_L g3155 ( 
.A(n_2622),
.Y(n_3155)
);

BUFx10_ASAP7_75t_L g3156 ( 
.A(n_2624),
.Y(n_3156)
);

INVx3_ASAP7_75t_L g3157 ( 
.A(n_2632),
.Y(n_3157)
);

NOR2xp33_ASAP7_75t_L g3158 ( 
.A(n_2498),
.B(n_273),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_2656),
.Y(n_3159)
);

INVx5_ASAP7_75t_L g3160 ( 
.A(n_2622),
.Y(n_3160)
);

BUFx2_ASAP7_75t_SL g3161 ( 
.A(n_2624),
.Y(n_3161)
);

INVx3_ASAP7_75t_SL g3162 ( 
.A(n_2626),
.Y(n_3162)
);

NAND2x1p5_ASAP7_75t_L g3163 ( 
.A(n_2612),
.B(n_2635),
.Y(n_3163)
);

INVx8_ASAP7_75t_L g3164 ( 
.A(n_2626),
.Y(n_3164)
);

BUFx6f_ASAP7_75t_L g3165 ( 
.A(n_2622),
.Y(n_3165)
);

INVx8_ASAP7_75t_L g3166 ( 
.A(n_2637),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2656),
.Y(n_3167)
);

BUFx6f_ASAP7_75t_L g3168 ( 
.A(n_2628),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2660),
.Y(n_3169)
);

BUFx3_ASAP7_75t_L g3170 ( 
.A(n_2441),
.Y(n_3170)
);

NAND2x1p5_ASAP7_75t_L g3171 ( 
.A(n_2670),
.B(n_273),
.Y(n_3171)
);

OR2x2_ASAP7_75t_L g3172 ( 
.A(n_2473),
.B(n_274),
.Y(n_3172)
);

BUFx3_ASAP7_75t_L g3173 ( 
.A(n_2442),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2660),
.Y(n_3174)
);

INVx6_ASAP7_75t_L g3175 ( 
.A(n_2708),
.Y(n_3175)
);

HB1xp67_ASAP7_75t_L g3176 ( 
.A(n_2305),
.Y(n_3176)
);

BUFx3_ASAP7_75t_L g3177 ( 
.A(n_2443),
.Y(n_3177)
);

INVx1_ASAP7_75t_SL g3178 ( 
.A(n_2606),
.Y(n_3178)
);

INVx6_ASAP7_75t_L g3179 ( 
.A(n_2637),
.Y(n_3179)
);

OR2x6_ASAP7_75t_L g3180 ( 
.A(n_2638),
.B(n_274),
.Y(n_3180)
);

HB1xp67_ASAP7_75t_L g3181 ( 
.A(n_2305),
.Y(n_3181)
);

BUFx12f_ASAP7_75t_L g3182 ( 
.A(n_2420),
.Y(n_3182)
);

CKINVDCx20_ASAP7_75t_R g3183 ( 
.A(n_2565),
.Y(n_3183)
);

BUFx3_ASAP7_75t_L g3184 ( 
.A(n_2638),
.Y(n_3184)
);

BUFx4_ASAP7_75t_SL g3185 ( 
.A(n_2664),
.Y(n_3185)
);

CKINVDCx16_ASAP7_75t_R g3186 ( 
.A(n_2325),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2739),
.B(n_275),
.Y(n_3187)
);

AND2x2_ASAP7_75t_L g3188 ( 
.A(n_2461),
.B(n_275),
.Y(n_3188)
);

INVx2_ASAP7_75t_SL g3189 ( 
.A(n_2639),
.Y(n_3189)
);

NAND2x1p5_ASAP7_75t_L g3190 ( 
.A(n_2639),
.B(n_276),
.Y(n_3190)
);

BUFx6f_ASAP7_75t_SL g3191 ( 
.A(n_2648),
.Y(n_3191)
);

BUFx4f_ASAP7_75t_SL g3192 ( 
.A(n_2700),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2664),
.Y(n_3193)
);

BUFx2_ASAP7_75t_L g3194 ( 
.A(n_2484),
.Y(n_3194)
);

INVx1_ASAP7_75t_SL g3195 ( 
.A(n_2786),
.Y(n_3195)
);

BUFx6f_ASAP7_75t_L g3196 ( 
.A(n_2628),
.Y(n_3196)
);

BUFx3_ASAP7_75t_L g3197 ( 
.A(n_2648),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2456),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_2466),
.Y(n_3199)
);

BUFx3_ASAP7_75t_L g3200 ( 
.A(n_2662),
.Y(n_3200)
);

INVx2_ASAP7_75t_SL g3201 ( 
.A(n_2662),
.Y(n_3201)
);

BUFx3_ASAP7_75t_L g3202 ( 
.A(n_2451),
.Y(n_3202)
);

CKINVDCx5p33_ASAP7_75t_R g3203 ( 
.A(n_2609),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2740),
.B(n_277),
.Y(n_3204)
);

INVx3_ASAP7_75t_L g3205 ( 
.A(n_2642),
.Y(n_3205)
);

INVx2_ASAP7_75t_SL g3206 ( 
.A(n_2420),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2671),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2671),
.Y(n_3208)
);

INVxp67_ASAP7_75t_SL g3209 ( 
.A(n_2341),
.Y(n_3209)
);

INVx4_ASAP7_75t_L g3210 ( 
.A(n_2323),
.Y(n_3210)
);

BUFx6f_ASAP7_75t_L g3211 ( 
.A(n_2628),
.Y(n_3211)
);

INVx3_ASAP7_75t_L g3212 ( 
.A(n_2642),
.Y(n_3212)
);

INVx3_ASAP7_75t_L g3213 ( 
.A(n_2615),
.Y(n_3213)
);

BUFx3_ASAP7_75t_L g3214 ( 
.A(n_2451),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2376),
.Y(n_3215)
);

INVx5_ASAP7_75t_L g3216 ( 
.A(n_2673),
.Y(n_3216)
);

BUFx2_ASAP7_75t_L g3217 ( 
.A(n_2770),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_2362),
.B(n_277),
.Y(n_3218)
);

BUFx2_ASAP7_75t_R g3219 ( 
.A(n_2507),
.Y(n_3219)
);

BUFx6f_ASAP7_75t_L g3220 ( 
.A(n_2673),
.Y(n_3220)
);

BUFx6f_ASAP7_75t_SL g3221 ( 
.A(n_2609),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2471),
.Y(n_3222)
);

BUFx6f_ASAP7_75t_L g3223 ( 
.A(n_2673),
.Y(n_3223)
);

INVx1_ASAP7_75t_SL g3224 ( 
.A(n_2789),
.Y(n_3224)
);

NAND2x1p5_ASAP7_75t_L g3225 ( 
.A(n_2323),
.B(n_279),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_2475),
.Y(n_3226)
);

INVxp67_ASAP7_75t_SL g3227 ( 
.A(n_2341),
.Y(n_3227)
);

CKINVDCx20_ASAP7_75t_R g3228 ( 
.A(n_2364),
.Y(n_3228)
);

BUFx6f_ASAP7_75t_L g3229 ( 
.A(n_2478),
.Y(n_3229)
);

CKINVDCx6p67_ASAP7_75t_R g3230 ( 
.A(n_2770),
.Y(n_3230)
);

BUFx6f_ASAP7_75t_L g3231 ( 
.A(n_2478),
.Y(n_3231)
);

BUFx3_ASAP7_75t_L g3232 ( 
.A(n_2777),
.Y(n_3232)
);

BUFx2_ASAP7_75t_L g3233 ( 
.A(n_2777),
.Y(n_3233)
);

BUFx3_ASAP7_75t_L g3234 ( 
.A(n_2782),
.Y(n_3234)
);

BUFx12f_ASAP7_75t_L g3235 ( 
.A(n_2782),
.Y(n_3235)
);

BUFx3_ASAP7_75t_L g3236 ( 
.A(n_2790),
.Y(n_3236)
);

BUFx6f_ASAP7_75t_L g3237 ( 
.A(n_2478),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2376),
.Y(n_3238)
);

INVx1_ASAP7_75t_SL g3239 ( 
.A(n_2791),
.Y(n_3239)
);

CKINVDCx11_ASAP7_75t_R g3240 ( 
.A(n_2801),
.Y(n_3240)
);

INVx3_ASAP7_75t_L g3241 ( 
.A(n_2901),
.Y(n_3241)
);

INVx3_ASAP7_75t_L g3242 ( 
.A(n_2901),
.Y(n_3242)
);

BUFx2_ASAP7_75t_R g3243 ( 
.A(n_2838),
.Y(n_3243)
);

CKINVDCx11_ASAP7_75t_R g3244 ( 
.A(n_2808),
.Y(n_3244)
);

CKINVDCx20_ASAP7_75t_R g3245 ( 
.A(n_2808),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_2803),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2991),
.Y(n_3247)
);

OAI22xp5_ASAP7_75t_L g3248 ( 
.A1(n_2832),
.A2(n_2467),
.B1(n_2435),
.B2(n_2790),
.Y(n_3248)
);

AOI22xp33_ASAP7_75t_L g3249 ( 
.A1(n_2966),
.A2(n_2299),
.B1(n_2793),
.B2(n_2452),
.Y(n_3249)
);

INVx1_ASAP7_75t_SL g3250 ( 
.A(n_3185),
.Y(n_3250)
);

AOI22xp33_ASAP7_75t_L g3251 ( 
.A1(n_2966),
.A2(n_2747),
.B1(n_2751),
.B2(n_2754),
.Y(n_3251)
);

INVx3_ASAP7_75t_L g3252 ( 
.A(n_2919),
.Y(n_3252)
);

INVxp67_ASAP7_75t_SL g3253 ( 
.A(n_2803),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2994),
.Y(n_3254)
);

OAI22xp5_ASAP7_75t_SL g3255 ( 
.A1(n_2927),
.A2(n_2636),
.B1(n_2370),
.B2(n_2486),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_2997),
.Y(n_3256)
);

AOI22xp5_ASAP7_75t_L g3257 ( 
.A1(n_3180),
.A2(n_2600),
.B1(n_2591),
.B2(n_2377),
.Y(n_3257)
);

INVx2_ASAP7_75t_L g3258 ( 
.A(n_2815),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_2840),
.B(n_2321),
.Y(n_3259)
);

BUFx4f_ASAP7_75t_SL g3260 ( 
.A(n_2814),
.Y(n_3260)
);

OAI22xp33_ASAP7_75t_L g3261 ( 
.A1(n_3116),
.A2(n_2426),
.B1(n_2302),
.B2(n_2503),
.Y(n_3261)
);

INVx6_ASAP7_75t_L g3262 ( 
.A(n_2816),
.Y(n_3262)
);

CKINVDCx11_ASAP7_75t_R g3263 ( 
.A(n_2819),
.Y(n_3263)
);

AOI22xp33_ASAP7_75t_SL g3264 ( 
.A1(n_3116),
.A2(n_2426),
.B1(n_2302),
.B2(n_2503),
.Y(n_3264)
);

AOI22xp33_ASAP7_75t_SL g3265 ( 
.A1(n_3164),
.A2(n_3166),
.B1(n_3161),
.B2(n_3145),
.Y(n_3265)
);

BUFx12f_ASAP7_75t_L g3266 ( 
.A(n_2811),
.Y(n_3266)
);

BUFx10_ASAP7_75t_L g3267 ( 
.A(n_2960),
.Y(n_3267)
);

CKINVDCx10_ASAP7_75t_R g3268 ( 
.A(n_2836),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2998),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3039),
.Y(n_3270)
);

INVx2_ASAP7_75t_SL g3271 ( 
.A(n_3185),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3047),
.Y(n_3272)
);

OAI22xp33_ASAP7_75t_R g3273 ( 
.A1(n_2913),
.A2(n_2745),
.B1(n_2404),
.B2(n_2571),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_2845),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2851),
.Y(n_3275)
);

CKINVDCx11_ASAP7_75t_R g3276 ( 
.A(n_2862),
.Y(n_3276)
);

CKINVDCx20_ASAP7_75t_R g3277 ( 
.A(n_2874),
.Y(n_3277)
);

NAND2x1p5_ASAP7_75t_L g3278 ( 
.A(n_2858),
.B(n_2343),
.Y(n_3278)
);

OAI22xp5_ASAP7_75t_L g3279 ( 
.A1(n_2832),
.A2(n_2857),
.B1(n_2909),
.B2(n_2854),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_2984),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2840),
.B(n_2361),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2868),
.Y(n_3282)
);

OAI22xp5_ASAP7_75t_SL g3283 ( 
.A1(n_3051),
.A2(n_2709),
.B1(n_2435),
.B2(n_2601),
.Y(n_3283)
);

INVxp67_ASAP7_75t_SL g3284 ( 
.A(n_2818),
.Y(n_3284)
);

AOI22xp33_ASAP7_75t_L g3285 ( 
.A1(n_2960),
.A2(n_2729),
.B1(n_2679),
.B2(n_2675),
.Y(n_3285)
);

INVx2_ASAP7_75t_L g3286 ( 
.A(n_3005),
.Y(n_3286)
);

BUFx4f_ASAP7_75t_SL g3287 ( 
.A(n_2802),
.Y(n_3287)
);

AOI22xp33_ASAP7_75t_SL g3288 ( 
.A1(n_3164),
.A2(n_2508),
.B1(n_2748),
.B2(n_2523),
.Y(n_3288)
);

AOI22xp33_ASAP7_75t_L g3289 ( 
.A1(n_2962),
.A2(n_2729),
.B1(n_2709),
.B2(n_2740),
.Y(n_3289)
);

CKINVDCx20_ASAP7_75t_R g3290 ( 
.A(n_2904),
.Y(n_3290)
);

INVx6_ASAP7_75t_L g3291 ( 
.A(n_2816),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_2884),
.Y(n_3292)
);

INVx3_ASAP7_75t_L g3293 ( 
.A(n_2919),
.Y(n_3293)
);

AOI22xp33_ASAP7_75t_SL g3294 ( 
.A1(n_3164),
.A2(n_2508),
.B1(n_2748),
.B2(n_2523),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3158),
.B(n_2792),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_3158),
.B(n_2795),
.Y(n_3296)
);

CKINVDCx11_ASAP7_75t_R g3297 ( 
.A(n_2820),
.Y(n_3297)
);

CKINVDCx11_ASAP7_75t_R g3298 ( 
.A(n_2820),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_2906),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_2923),
.Y(n_3300)
);

OAI22xp5_ASAP7_75t_L g3301 ( 
.A1(n_2854),
.A2(n_2584),
.B1(n_2608),
.B2(n_2601),
.Y(n_3301)
);

OAI22xp33_ASAP7_75t_L g3302 ( 
.A1(n_3180),
.A2(n_2646),
.B1(n_2645),
.B2(n_2527),
.Y(n_3302)
);

AND2x2_ASAP7_75t_L g3303 ( 
.A(n_2911),
.B(n_2800),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3014),
.Y(n_3304)
);

BUFx12f_ASAP7_75t_L g3305 ( 
.A(n_2867),
.Y(n_3305)
);

CKINVDCx6p67_ASAP7_75t_R g3306 ( 
.A(n_2959),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2925),
.Y(n_3307)
);

AOI22xp33_ASAP7_75t_L g3308 ( 
.A1(n_2962),
.A2(n_2608),
.B1(n_2584),
.B2(n_2418),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_2972),
.B(n_2403),
.Y(n_3309)
);

INVx2_ASAP7_75t_SL g3310 ( 
.A(n_2970),
.Y(n_3310)
);

OAI22xp33_ASAP7_75t_L g3311 ( 
.A1(n_3180),
.A2(n_2518),
.B1(n_2527),
.B2(n_2439),
.Y(n_3311)
);

CKINVDCx20_ASAP7_75t_R g3312 ( 
.A(n_2904),
.Y(n_3312)
);

BUFx2_ASAP7_75t_L g3313 ( 
.A(n_2965),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_2929),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3072),
.Y(n_3315)
);

OAI22xp33_ASAP7_75t_L g3316 ( 
.A1(n_2932),
.A2(n_3162),
.B1(n_3127),
.B2(n_3011),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_3016),
.Y(n_3317)
);

AOI22xp33_ASAP7_75t_L g3318 ( 
.A1(n_2965),
.A2(n_2993),
.B1(n_2980),
.B2(n_2898),
.Y(n_3318)
);

BUFx2_ASAP7_75t_L g3319 ( 
.A(n_3063),
.Y(n_3319)
);

AOI22xp33_ASAP7_75t_SL g3320 ( 
.A1(n_3166),
.A2(n_2508),
.B1(n_2518),
.B2(n_2548),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3088),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3019),
.Y(n_3322)
);

OAI22xp33_ASAP7_75t_L g3323 ( 
.A1(n_2932),
.A2(n_2720),
.B1(n_2738),
.B2(n_2589),
.Y(n_3323)
);

CKINVDCx20_ASAP7_75t_R g3324 ( 
.A(n_2853),
.Y(n_3324)
);

BUFx3_ASAP7_75t_L g3325 ( 
.A(n_2895),
.Y(n_3325)
);

BUFx12f_ASAP7_75t_L g3326 ( 
.A(n_2918),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3090),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3108),
.Y(n_3328)
);

OR2x2_ASAP7_75t_L g3329 ( 
.A(n_2821),
.B(n_2589),
.Y(n_3329)
);

AOI22xp33_ASAP7_75t_L g3330 ( 
.A1(n_2980),
.A2(n_2497),
.B1(n_2477),
.B2(n_2408),
.Y(n_3330)
);

BUFx12f_ASAP7_75t_L g3331 ( 
.A(n_3046),
.Y(n_3331)
);

BUFx2_ASAP7_75t_L g3332 ( 
.A(n_3063),
.Y(n_3332)
);

AOI22xp33_ASAP7_75t_L g3333 ( 
.A1(n_2980),
.A2(n_2500),
.B1(n_2561),
.B2(n_2538),
.Y(n_3333)
);

AOI22xp33_ASAP7_75t_L g3334 ( 
.A1(n_2993),
.A2(n_2536),
.B1(n_2410),
.B2(n_2409),
.Y(n_3334)
);

AOI22xp33_ASAP7_75t_SL g3335 ( 
.A1(n_3166),
.A2(n_2508),
.B1(n_2618),
.B2(n_2548),
.Y(n_3335)
);

CKINVDCx20_ASAP7_75t_R g3336 ( 
.A(n_3183),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3109),
.Y(n_3337)
);

AOI22xp33_ASAP7_75t_L g3338 ( 
.A1(n_2993),
.A2(n_2410),
.B1(n_2409),
.B2(n_2734),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_3042),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3111),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3114),
.Y(n_3341)
);

CKINVDCx6p67_ASAP7_75t_R g3342 ( 
.A(n_2886),
.Y(n_3342)
);

INVx3_ASAP7_75t_L g3343 ( 
.A(n_2981),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3117),
.Y(n_3344)
);

BUFx2_ASAP7_75t_L g3345 ( 
.A(n_2893),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3133),
.Y(n_3346)
);

BUFx3_ASAP7_75t_L g3347 ( 
.A(n_2892),
.Y(n_3347)
);

INVx3_ASAP7_75t_L g3348 ( 
.A(n_2981),
.Y(n_3348)
);

OAI22xp5_ASAP7_75t_L g3349 ( 
.A1(n_2857),
.A2(n_2343),
.B1(n_2762),
.B2(n_2684),
.Y(n_3349)
);

NAND2x1_ASAP7_75t_L g3350 ( 
.A(n_2908),
.B(n_2700),
.Y(n_3350)
);

NAND2x1p5_ASAP7_75t_L g3351 ( 
.A(n_2858),
.B(n_2298),
.Y(n_3351)
);

OAI22xp33_ASAP7_75t_L g3352 ( 
.A1(n_2932),
.A2(n_3162),
.B1(n_3127),
.B2(n_3011),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3138),
.Y(n_3353)
);

AOI22xp33_ASAP7_75t_L g3354 ( 
.A1(n_2938),
.A2(n_2969),
.B1(n_3153),
.B2(n_3146),
.Y(n_3354)
);

OAI22xp5_ASAP7_75t_L g3355 ( 
.A1(n_2909),
.A2(n_2683),
.B1(n_2701),
.B2(n_2627),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3150),
.Y(n_3356)
);

BUFx12f_ASAP7_75t_L g3357 ( 
.A(n_2805),
.Y(n_3357)
);

INVx2_ASAP7_75t_R g3358 ( 
.A(n_2942),
.Y(n_3358)
);

OAI22xp5_ASAP7_75t_L g3359 ( 
.A1(n_3186),
.A2(n_2701),
.B1(n_2627),
.B2(n_2711),
.Y(n_3359)
);

BUFx12f_ASAP7_75t_L g3360 ( 
.A(n_2805),
.Y(n_3360)
);

CKINVDCx20_ASAP7_75t_R g3361 ( 
.A(n_3228),
.Y(n_3361)
);

OAI22xp33_ASAP7_75t_SL g3362 ( 
.A1(n_3190),
.A2(n_2618),
.B1(n_2759),
.B2(n_2726),
.Y(n_3362)
);

OAI22xp5_ASAP7_75t_L g3363 ( 
.A1(n_2818),
.A2(n_2711),
.B1(n_2541),
.B2(n_2547),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3154),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3169),
.Y(n_3365)
);

AOI22xp33_ASAP7_75t_L g3366 ( 
.A1(n_2969),
.A2(n_3146),
.B1(n_3191),
.B2(n_3153),
.Y(n_3366)
);

BUFx3_ASAP7_75t_L g3367 ( 
.A(n_2810),
.Y(n_3367)
);

AOI22xp33_ASAP7_75t_SL g3368 ( 
.A1(n_3011),
.A2(n_2715),
.B1(n_2757),
.B2(n_2605),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3174),
.Y(n_3369)
);

AOI22xp5_ASAP7_75t_L g3370 ( 
.A1(n_3191),
.A2(n_2579),
.B1(n_2617),
.B2(n_2725),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3107),
.Y(n_3371)
);

AOI22xp33_ASAP7_75t_L g3372 ( 
.A1(n_3221),
.A2(n_2870),
.B1(n_3023),
.B2(n_3021),
.Y(n_3372)
);

INVx6_ASAP7_75t_L g3373 ( 
.A(n_2858),
.Y(n_3373)
);

AOI22xp33_ASAP7_75t_SL g3374 ( 
.A1(n_3041),
.A2(n_2554),
.B1(n_2707),
.B2(n_2705),
.Y(n_3374)
);

BUFx3_ASAP7_75t_L g3375 ( 
.A(n_2822),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3193),
.Y(n_3376)
);

BUFx3_ASAP7_75t_L g3377 ( 
.A(n_2844),
.Y(n_3377)
);

CKINVDCx11_ASAP7_75t_R g3378 ( 
.A(n_2957),
.Y(n_3378)
);

AOI22xp33_ASAP7_75t_SL g3379 ( 
.A1(n_3041),
.A2(n_2463),
.B1(n_2474),
.B2(n_2598),
.Y(n_3379)
);

AOI22xp33_ASAP7_75t_L g3380 ( 
.A1(n_3221),
.A2(n_2593),
.B1(n_2588),
.B2(n_2693),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3215),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3238),
.Y(n_3382)
);

AOI22xp33_ASAP7_75t_L g3383 ( 
.A1(n_2870),
.A2(n_2593),
.B1(n_2588),
.B2(n_2351),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3124),
.Y(n_3384)
);

CKINVDCx20_ASAP7_75t_R g3385 ( 
.A(n_3120),
.Y(n_3385)
);

AOI22xp33_ASAP7_75t_SL g3386 ( 
.A1(n_3041),
.A2(n_2513),
.B1(n_2522),
.B2(n_2488),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_2952),
.B(n_2423),
.Y(n_3387)
);

AOI22xp33_ASAP7_75t_L g3388 ( 
.A1(n_2870),
.A2(n_2351),
.B1(n_2712),
.B2(n_2556),
.Y(n_3388)
);

OAI22xp33_ASAP7_75t_L g3389 ( 
.A1(n_3203),
.A2(n_2383),
.B1(n_2491),
.B2(n_2529),
.Y(n_3389)
);

INVx6_ASAP7_75t_L g3390 ( 
.A(n_2970),
.Y(n_3390)
);

INVxp67_ASAP7_75t_L g3391 ( 
.A(n_2876),
.Y(n_3391)
);

OAI22xp33_ASAP7_75t_L g3392 ( 
.A1(n_3068),
.A2(n_2533),
.B1(n_2542),
.B2(n_2531),
.Y(n_3392)
);

BUFx6f_ASAP7_75t_L g3393 ( 
.A(n_2942),
.Y(n_3393)
);

AOI22xp33_ASAP7_75t_L g3394 ( 
.A1(n_3103),
.A2(n_2332),
.B1(n_2753),
.B2(n_2634),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3126),
.Y(n_3395)
);

OAI22xp5_ASAP7_75t_L g3396 ( 
.A1(n_3195),
.A2(n_2512),
.B1(n_2744),
.B2(n_2767),
.Y(n_3396)
);

BUFx8_ASAP7_75t_L g3397 ( 
.A(n_2804),
.Y(n_3397)
);

BUFx12f_ASAP7_75t_L g3398 ( 
.A(n_3027),
.Y(n_3398)
);

BUFx2_ASAP7_75t_L g3399 ( 
.A(n_2893),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_2952),
.B(n_2423),
.Y(n_3400)
);

AOI22xp33_ASAP7_75t_L g3401 ( 
.A1(n_3103),
.A2(n_2753),
.B1(n_2566),
.B2(n_2655),
.Y(n_3401)
);

BUFx4f_ASAP7_75t_SL g3402 ( 
.A(n_2826),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3129),
.Y(n_3403)
);

BUFx12f_ASAP7_75t_L g3404 ( 
.A(n_2899),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_3147),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_3151),
.Y(n_3406)
);

INVx1_ASAP7_75t_SL g3407 ( 
.A(n_2913),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3159),
.Y(n_3408)
);

AOI22xp5_ASAP7_75t_SL g3409 ( 
.A1(n_3075),
.A2(n_2317),
.B1(n_2651),
.B2(n_2320),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3167),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_2807),
.Y(n_3411)
);

INVx4_ASAP7_75t_L g3412 ( 
.A(n_2970),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_2833),
.Y(n_3413)
);

OAI22xp5_ASAP7_75t_L g3414 ( 
.A1(n_3195),
.A2(n_2767),
.B1(n_2459),
.B2(n_2495),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_2934),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_2936),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_2846),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_2939),
.Y(n_3418)
);

INVx1_ASAP7_75t_SL g3419 ( 
.A(n_2852),
.Y(n_3419)
);

BUFx3_ASAP7_75t_L g3420 ( 
.A(n_2849),
.Y(n_3420)
);

BUFx8_ASAP7_75t_L g3421 ( 
.A(n_2890),
.Y(n_3421)
);

AOI22xp5_ASAP7_75t_L g3422 ( 
.A1(n_3065),
.A2(n_2437),
.B1(n_2482),
.B2(n_2464),
.Y(n_3422)
);

INVx6_ASAP7_75t_L g3423 ( 
.A(n_2824),
.Y(n_3423)
);

BUFx2_ASAP7_75t_L g3424 ( 
.A(n_2826),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_2855),
.Y(n_3425)
);

INVx5_ASAP7_75t_L g3426 ( 
.A(n_2809),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_2872),
.Y(n_3427)
);

BUFx3_ASAP7_75t_L g3428 ( 
.A(n_2850),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_2872),
.Y(n_3429)
);

INVx5_ASAP7_75t_L g3430 ( 
.A(n_2809),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3135),
.B(n_2454),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_2953),
.Y(n_3432)
);

CKINVDCx20_ASAP7_75t_R g3433 ( 
.A(n_3000),
.Y(n_3433)
);

CKINVDCx11_ASAP7_75t_R g3434 ( 
.A(n_2974),
.Y(n_3434)
);

INVx2_ASAP7_75t_SL g3435 ( 
.A(n_3025),
.Y(n_3435)
);

AOI22xp33_ASAP7_75t_L g3436 ( 
.A1(n_3175),
.A2(n_2459),
.B1(n_2495),
.B2(n_2736),
.Y(n_3436)
);

BUFx2_ASAP7_75t_L g3437 ( 
.A(n_3092),
.Y(n_3437)
);

AOI22xp33_ASAP7_75t_L g3438 ( 
.A1(n_3175),
.A2(n_2429),
.B1(n_2401),
.B2(n_2412),
.Y(n_3438)
);

INVx6_ASAP7_75t_L g3439 ( 
.A(n_2824),
.Y(n_3439)
);

BUFx3_ASAP7_75t_L g3440 ( 
.A(n_2885),
.Y(n_3440)
);

AOI22xp33_ASAP7_75t_L g3441 ( 
.A1(n_3056),
.A2(n_2429),
.B1(n_2434),
.B2(n_2399),
.Y(n_3441)
);

BUFx3_ASAP7_75t_L g3442 ( 
.A(n_2894),
.Y(n_3442)
);

OAI21xp5_ASAP7_75t_SL g3443 ( 
.A1(n_2825),
.A2(n_2761),
.B(n_2514),
.Y(n_3443)
);

INVx3_ASAP7_75t_L g3444 ( 
.A(n_2981),
.Y(n_3444)
);

INVx1_ASAP7_75t_SL g3445 ( 
.A(n_2887),
.Y(n_3445)
);

AOI22xp33_ASAP7_75t_L g3446 ( 
.A1(n_2837),
.A2(n_2453),
.B1(n_2444),
.B2(n_2585),
.Y(n_3446)
);

INVx4_ASAP7_75t_L g3447 ( 
.A(n_3092),
.Y(n_3447)
);

OAI22xp5_ASAP7_75t_L g3448 ( 
.A1(n_3224),
.A2(n_3239),
.B1(n_3190),
.B2(n_3230),
.Y(n_3448)
);

OAI22xp33_ASAP7_75t_L g3449 ( 
.A1(n_3061),
.A2(n_2742),
.B1(n_2496),
.B2(n_2519),
.Y(n_3449)
);

CKINVDCx11_ASAP7_75t_R g3450 ( 
.A(n_3004),
.Y(n_3450)
);

INVx6_ASAP7_75t_L g3451 ( 
.A(n_2828),
.Y(n_3451)
);

AOI22xp33_ASAP7_75t_L g3452 ( 
.A1(n_2837),
.A2(n_2865),
.B1(n_3025),
.B2(n_3235),
.Y(n_3452)
);

BUFx2_ASAP7_75t_L g3453 ( 
.A(n_2863),
.Y(n_3453)
);

BUFx10_ASAP7_75t_L g3454 ( 
.A(n_2896),
.Y(n_3454)
);

AOI22xp33_ASAP7_75t_L g3455 ( 
.A1(n_2837),
.A2(n_2599),
.B1(n_2633),
.B2(n_2595),
.Y(n_3455)
);

AOI22xp33_ASAP7_75t_SL g3456 ( 
.A1(n_2865),
.A2(n_2766),
.B1(n_2710),
.B2(n_2688),
.Y(n_3456)
);

INVxp67_ASAP7_75t_SL g3457 ( 
.A(n_2930),
.Y(n_3457)
);

CKINVDCx5p33_ASAP7_75t_R g3458 ( 
.A(n_2848),
.Y(n_3458)
);

CKINVDCx6p67_ASAP7_75t_R g3459 ( 
.A(n_2924),
.Y(n_3459)
);

OAI22x1_ASAP7_75t_L g3460 ( 
.A1(n_2813),
.A2(n_2806),
.B1(n_2915),
.B2(n_3105),
.Y(n_3460)
);

BUFx3_ASAP7_75t_L g3461 ( 
.A(n_2985),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_2963),
.Y(n_3462)
);

CKINVDCx11_ASAP7_75t_R g3463 ( 
.A(n_3038),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_2967),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_2856),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_2875),
.Y(n_3466)
);

AND2x4_ASAP7_75t_L g3467 ( 
.A(n_2981),
.B(n_2454),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_2883),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_2888),
.Y(n_3469)
);

CKINVDCx20_ASAP7_75t_R g3470 ( 
.A(n_2865),
.Y(n_3470)
);

AOI22xp33_ASAP7_75t_L g3471 ( 
.A1(n_3152),
.A2(n_2689),
.B1(n_2694),
.B2(n_2685),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_2903),
.Y(n_3472)
);

AOI22xp33_ASAP7_75t_SL g3473 ( 
.A1(n_2928),
.A2(n_2710),
.B1(n_2688),
.B2(n_2384),
.Y(n_3473)
);

BUFx3_ASAP7_75t_L g3474 ( 
.A(n_2995),
.Y(n_3474)
);

OAI22xp5_ASAP7_75t_L g3475 ( 
.A1(n_3239),
.A2(n_2519),
.B1(n_2379),
.B2(n_2572),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_2910),
.Y(n_3476)
);

BUFx3_ASAP7_75t_L g3477 ( 
.A(n_2864),
.Y(n_3477)
);

BUFx6f_ASAP7_75t_L g3478 ( 
.A(n_2942),
.Y(n_3478)
);

CKINVDCx5p33_ASAP7_75t_R g3479 ( 
.A(n_2848),
.Y(n_3479)
);

OAI22xp33_ASAP7_75t_L g3480 ( 
.A1(n_2813),
.A2(n_3101),
.B1(n_2806),
.B2(n_3050),
.Y(n_3480)
);

BUFx6f_ASAP7_75t_L g3481 ( 
.A(n_2942),
.Y(n_3481)
);

INVx6_ASAP7_75t_L g3482 ( 
.A(n_2828),
.Y(n_3482)
);

OAI22xp5_ASAP7_75t_L g3483 ( 
.A1(n_3224),
.A2(n_2379),
.B1(n_2574),
.B2(n_2331),
.Y(n_3483)
);

BUFx2_ASAP7_75t_SL g3484 ( 
.A(n_2916),
.Y(n_3484)
);

INVx6_ASAP7_75t_L g3485 ( 
.A(n_2871),
.Y(n_3485)
);

OAI21xp5_ASAP7_75t_SL g3486 ( 
.A1(n_2825),
.A2(n_2761),
.B(n_2743),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3135),
.B(n_2501),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_2922),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_2951),
.Y(n_3489)
);

INVx4_ASAP7_75t_L g3490 ( 
.A(n_3028),
.Y(n_3490)
);

HB1xp67_ASAP7_75t_L g3491 ( 
.A(n_3194),
.Y(n_3491)
);

INVxp67_ASAP7_75t_SL g3492 ( 
.A(n_2930),
.Y(n_3492)
);

BUFx6f_ASAP7_75t_L g3493 ( 
.A(n_2950),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3089),
.B(n_2891),
.Y(n_3494)
);

INVx2_ASAP7_75t_SL g3495 ( 
.A(n_3101),
.Y(n_3495)
);

INVx1_ASAP7_75t_SL g3496 ( 
.A(n_2821),
.Y(n_3496)
);

INVx4_ASAP7_75t_L g3497 ( 
.A(n_3028),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3089),
.B(n_2501),
.Y(n_3498)
);

BUFx12f_ASAP7_75t_L g3499 ( 
.A(n_3081),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3049),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_2891),
.B(n_2421),
.Y(n_3501)
);

BUFx8_ASAP7_75t_L g3502 ( 
.A(n_3010),
.Y(n_3502)
);

BUFx12f_ASAP7_75t_L g3503 ( 
.A(n_3115),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_L g3504 ( 
.A1(n_3182),
.A2(n_2388),
.B1(n_2385),
.B2(n_2681),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3037),
.B(n_2334),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_SL g3506 ( 
.A(n_2917),
.B(n_2796),
.Y(n_3506)
);

AOI22xp33_ASAP7_75t_L g3507 ( 
.A1(n_3123),
.A2(n_2340),
.B1(n_2562),
.B2(n_2546),
.Y(n_3507)
);

AOI22xp33_ASAP7_75t_L g3508 ( 
.A1(n_3139),
.A2(n_2575),
.B1(n_2778),
.B2(n_2312),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3037),
.B(n_2780),
.Y(n_3509)
);

OAI22xp33_ASAP7_75t_SL g3510 ( 
.A1(n_3179),
.A2(n_2329),
.B1(n_2781),
.B2(n_2499),
.Y(n_3510)
);

CKINVDCx20_ASAP7_75t_R g3511 ( 
.A(n_3084),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3053),
.Y(n_3512)
);

AOI22xp33_ASAP7_75t_L g3513 ( 
.A1(n_3143),
.A2(n_2752),
.B1(n_2650),
.B2(n_2647),
.Y(n_3513)
);

INVx6_ASAP7_75t_L g3514 ( 
.A(n_2871),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3074),
.Y(n_3515)
);

BUFx12f_ASAP7_75t_L g3516 ( 
.A(n_3156),
.Y(n_3516)
);

INVx6_ASAP7_75t_L g3517 ( 
.A(n_3156),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3091),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3095),
.Y(n_3519)
);

INVx4_ASAP7_75t_L g3520 ( 
.A(n_3028),
.Y(n_3520)
);

CKINVDCx11_ASAP7_75t_R g3521 ( 
.A(n_2947),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3198),
.Y(n_3522)
);

INVx1_ASAP7_75t_SL g3523 ( 
.A(n_2823),
.Y(n_3523)
);

OAI22xp5_ASAP7_75t_L g3524 ( 
.A1(n_2973),
.A2(n_2384),
.B1(n_2397),
.B2(n_2396),
.Y(n_3524)
);

BUFx12f_ASAP7_75t_L g3525 ( 
.A(n_2839),
.Y(n_3525)
);

BUFx2_ASAP7_75t_SL g3526 ( 
.A(n_3028),
.Y(n_3526)
);

BUFx2_ASAP7_75t_SL g3527 ( 
.A(n_3032),
.Y(n_3527)
);

BUFx6f_ASAP7_75t_L g3528 ( 
.A(n_2950),
.Y(n_3528)
);

INVx6_ASAP7_75t_L g3529 ( 
.A(n_2958),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3199),
.Y(n_3530)
);

HB1xp67_ASAP7_75t_L g3531 ( 
.A(n_2823),
.Y(n_3531)
);

INVx3_ASAP7_75t_L g3532 ( 
.A(n_3032),
.Y(n_3532)
);

HB1xp67_ASAP7_75t_L g3533 ( 
.A(n_2880),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3222),
.Y(n_3534)
);

HB1xp67_ASAP7_75t_L g3535 ( 
.A(n_2880),
.Y(n_3535)
);

CKINVDCx20_ASAP7_75t_R g3536 ( 
.A(n_3097),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3226),
.Y(n_3537)
);

BUFx12f_ASAP7_75t_L g3538 ( 
.A(n_2839),
.Y(n_3538)
);

BUFx10_ASAP7_75t_L g3539 ( 
.A(n_2989),
.Y(n_3539)
);

INVx3_ASAP7_75t_L g3540 ( 
.A(n_3032),
.Y(n_3540)
);

AOI22xp33_ASAP7_75t_SL g3541 ( 
.A1(n_2940),
.A2(n_2396),
.B1(n_2407),
.B2(n_2397),
.Y(n_3541)
);

BUFx4f_ASAP7_75t_SL g3542 ( 
.A(n_2955),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_2827),
.Y(n_3543)
);

CKINVDCx5p33_ASAP7_75t_R g3544 ( 
.A(n_3099),
.Y(n_3544)
);

AOI22xp33_ASAP7_75t_SL g3545 ( 
.A1(n_3179),
.A2(n_2407),
.B1(n_2615),
.B2(n_2549),
.Y(n_3545)
);

OAI22xp33_ASAP7_75t_L g3546 ( 
.A1(n_3184),
.A2(n_2665),
.B1(n_2658),
.B2(n_2506),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_SL g3547 ( 
.A1(n_3209),
.A2(n_2549),
.B(n_2528),
.Y(n_3547)
);

CKINVDCx5p33_ASAP7_75t_R g3548 ( 
.A(n_3099),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_2897),
.B(n_2494),
.Y(n_3549)
);

AOI22xp33_ASAP7_75t_SL g3550 ( 
.A1(n_3060),
.A2(n_2528),
.B1(n_2737),
.B2(n_2732),
.Y(n_3550)
);

OAI22xp5_ASAP7_75t_L g3551 ( 
.A1(n_2973),
.A2(n_2756),
.B1(n_2765),
.B2(n_2749),
.Y(n_3551)
);

OAI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_3006),
.A2(n_2765),
.B(n_2796),
.Y(n_3552)
);

BUFx6f_ASAP7_75t_L g3553 ( 
.A(n_2950),
.Y(n_3553)
);

CKINVDCx20_ASAP7_75t_R g3554 ( 
.A(n_3067),
.Y(n_3554)
);

CKINVDCx11_ASAP7_75t_R g3555 ( 
.A(n_2956),
.Y(n_3555)
);

BUFx12f_ASAP7_75t_L g3556 ( 
.A(n_2961),
.Y(n_3556)
);

AOI22xp33_ASAP7_75t_L g3557 ( 
.A1(n_3132),
.A2(n_2481),
.B1(n_2674),
.B2(n_2760),
.Y(n_3557)
);

BUFx10_ASAP7_75t_L g3558 ( 
.A(n_2989),
.Y(n_3558)
);

INVx8_ASAP7_75t_L g3559 ( 
.A(n_3032),
.Y(n_3559)
);

BUFx3_ASAP7_75t_L g3560 ( 
.A(n_2914),
.Y(n_3560)
);

AOI22xp33_ASAP7_75t_L g3561 ( 
.A1(n_2817),
.A2(n_2481),
.B1(n_2760),
.B2(n_2763),
.Y(n_3561)
);

INVx2_ASAP7_75t_SL g3562 ( 
.A(n_2931),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_2979),
.Y(n_3563)
);

BUFx8_ASAP7_75t_SL g3564 ( 
.A(n_3080),
.Y(n_3564)
);

INVx2_ASAP7_75t_L g3565 ( 
.A(n_2827),
.Y(n_3565)
);

BUFx10_ASAP7_75t_L g3566 ( 
.A(n_3064),
.Y(n_3566)
);

BUFx10_ASAP7_75t_L g3567 ( 
.A(n_3064),
.Y(n_3567)
);

OAI22xp5_ASAP7_75t_L g3568 ( 
.A1(n_2976),
.A2(n_2764),
.B1(n_2654),
.B2(n_2661),
.Y(n_3568)
);

OAI22xp5_ASAP7_75t_L g3569 ( 
.A1(n_2976),
.A2(n_2654),
.B1(n_2661),
.B2(n_2614),
.Y(n_3569)
);

INVx1_ASAP7_75t_SL g3570 ( 
.A(n_2992),
.Y(n_3570)
);

CKINVDCx11_ASAP7_75t_R g3571 ( 
.A(n_3170),
.Y(n_3571)
);

AOI22xp33_ASAP7_75t_L g3572 ( 
.A1(n_2817),
.A2(n_2697),
.B1(n_2698),
.B2(n_2691),
.Y(n_3572)
);

AOI22xp33_ASAP7_75t_L g3573 ( 
.A1(n_3217),
.A2(n_2697),
.B1(n_2733),
.B2(n_2594),
.Y(n_3573)
);

INVx1_ASAP7_75t_SL g3574 ( 
.A(n_3002),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_2979),
.Y(n_3575)
);

INVx4_ASAP7_75t_L g3576 ( 
.A(n_3192),
.Y(n_3576)
);

BUFx10_ASAP7_75t_L g3577 ( 
.A(n_2869),
.Y(n_3577)
);

BUFx3_ASAP7_75t_L g3578 ( 
.A(n_2943),
.Y(n_3578)
);

INVx6_ASAP7_75t_L g3579 ( 
.A(n_3048),
.Y(n_3579)
);

INVx2_ASAP7_75t_SL g3580 ( 
.A(n_3173),
.Y(n_3580)
);

OAI22xp5_ASAP7_75t_L g3581 ( 
.A1(n_2982),
.A2(n_2324),
.B1(n_2347),
.B2(n_2346),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_2990),
.Y(n_3582)
);

BUFx10_ASAP7_75t_L g3583 ( 
.A(n_2920),
.Y(n_3583)
);

INVx2_ASAP7_75t_L g3584 ( 
.A(n_2829),
.Y(n_3584)
);

AOI22xp33_ASAP7_75t_L g3585 ( 
.A1(n_3233),
.A2(n_2733),
.B1(n_2611),
.B2(n_2590),
.Y(n_3585)
);

CKINVDCx11_ASAP7_75t_R g3586 ( 
.A(n_3177),
.Y(n_3586)
);

AOI22xp33_ASAP7_75t_L g3587 ( 
.A1(n_3134),
.A2(n_2733),
.B1(n_2348),
.B2(n_2363),
.Y(n_3587)
);

AOI22xp33_ASAP7_75t_SL g3588 ( 
.A1(n_2933),
.A2(n_2733),
.B1(n_2779),
.B2(n_2359),
.Y(n_3588)
);

INVx2_ASAP7_75t_SL g3589 ( 
.A(n_3054),
.Y(n_3589)
);

AOI22xp33_ASAP7_75t_L g3590 ( 
.A1(n_3137),
.A2(n_2733),
.B1(n_2746),
.B2(n_2724),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_2829),
.Y(n_3591)
);

BUFx3_ASAP7_75t_L g3592 ( 
.A(n_2948),
.Y(n_3592)
);

BUFx3_ASAP7_75t_L g3593 ( 
.A(n_3022),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_2842),
.Y(n_3594)
);

INVx1_ASAP7_75t_SL g3595 ( 
.A(n_2861),
.Y(n_3595)
);

OAI22xp5_ASAP7_75t_L g3596 ( 
.A1(n_2982),
.A2(n_2359),
.B1(n_2386),
.B2(n_2367),
.Y(n_3596)
);

AOI22xp33_ASAP7_75t_L g3597 ( 
.A1(n_3144),
.A2(n_2746),
.B1(n_2724),
.B2(n_2413),
.Y(n_3597)
);

INVx1_ASAP7_75t_SL g3598 ( 
.A(n_2861),
.Y(n_3598)
);

BUFx2_ASAP7_75t_SL g3599 ( 
.A(n_2996),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3008),
.Y(n_3600)
);

OAI22xp5_ASAP7_75t_L g3601 ( 
.A1(n_3264),
.A2(n_3219),
.B1(n_3036),
.B2(n_3024),
.Y(n_3601)
);

AND2x2_ASAP7_75t_L g3602 ( 
.A(n_3303),
.B(n_2866),
.Y(n_3602)
);

HB1xp67_ASAP7_75t_L g3603 ( 
.A(n_3491),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3247),
.Y(n_3604)
);

BUFx12f_ASAP7_75t_L g3605 ( 
.A(n_3240),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3254),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3600),
.B(n_2900),
.Y(n_3607)
);

BUFx6f_ASAP7_75t_L g3608 ( 
.A(n_3559),
.Y(n_3608)
);

BUFx4f_ASAP7_75t_SL g3609 ( 
.A(n_3398),
.Y(n_3609)
);

INVx2_ASAP7_75t_SL g3610 ( 
.A(n_3397),
.Y(n_3610)
);

OAI22xp5_ASAP7_75t_L g3611 ( 
.A1(n_3301),
.A2(n_3219),
.B1(n_3036),
.B2(n_3024),
.Y(n_3611)
);

BUFx8_ASAP7_75t_SL g3612 ( 
.A(n_3245),
.Y(n_3612)
);

NAND3xp33_ASAP7_75t_L g3613 ( 
.A(n_3249),
.B(n_2841),
.C(n_2835),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3256),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3269),
.Y(n_3615)
);

INVx2_ASAP7_75t_L g3616 ( 
.A(n_3322),
.Y(n_3616)
);

AOI22xp33_ASAP7_75t_L g3617 ( 
.A1(n_3460),
.A2(n_2907),
.B1(n_2834),
.B2(n_2841),
.Y(n_3617)
);

BUFx6f_ASAP7_75t_L g3618 ( 
.A(n_3559),
.Y(n_3618)
);

AOI22xp33_ASAP7_75t_L g3619 ( 
.A1(n_3480),
.A2(n_2907),
.B1(n_2835),
.B2(n_2905),
.Y(n_3619)
);

HB1xp67_ASAP7_75t_L g3620 ( 
.A(n_3533),
.Y(n_3620)
);

OAI21xp33_ASAP7_75t_L g3621 ( 
.A1(n_3443),
.A2(n_2905),
.B(n_3017),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3270),
.Y(n_3622)
);

BUFx6f_ASAP7_75t_L g3623 ( 
.A(n_3393),
.Y(n_3623)
);

INVx2_ASAP7_75t_SL g3624 ( 
.A(n_3397),
.Y(n_3624)
);

AND2x2_ASAP7_75t_L g3625 ( 
.A(n_3570),
.B(n_2921),
.Y(n_3625)
);

BUFx3_ASAP7_75t_L g3626 ( 
.A(n_3554),
.Y(n_3626)
);

AOI22xp33_ASAP7_75t_L g3627 ( 
.A1(n_3273),
.A2(n_2954),
.B1(n_3030),
.B2(n_3197),
.Y(n_3627)
);

OAI21xp5_ASAP7_75t_SL g3628 ( 
.A1(n_3250),
.A2(n_2831),
.B(n_3105),
.Y(n_3628)
);

OAI22xp33_ASAP7_75t_L g3629 ( 
.A1(n_3271),
.A2(n_3110),
.B1(n_3033),
.B2(n_2986),
.Y(n_3629)
);

OAI22xp5_ASAP7_75t_L g3630 ( 
.A1(n_3320),
.A2(n_3033),
.B1(n_2986),
.B2(n_3200),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3339),
.Y(n_3631)
);

AOI22xp33_ASAP7_75t_L g3632 ( 
.A1(n_3255),
.A2(n_3234),
.B1(n_3236),
.B2(n_3232),
.Y(n_3632)
);

OAI22xp5_ASAP7_75t_L g3633 ( 
.A1(n_3288),
.A2(n_3209),
.B1(n_3227),
.B2(n_3110),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3272),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3274),
.Y(n_3635)
);

AOI22xp33_ASAP7_75t_L g3636 ( 
.A1(n_3283),
.A2(n_3189),
.B1(n_3201),
.B2(n_2949),
.Y(n_3636)
);

AOI22xp33_ASAP7_75t_L g3637 ( 
.A1(n_3494),
.A2(n_3070),
.B1(n_3082),
.B2(n_3176),
.Y(n_3637)
);

BUFx4f_ASAP7_75t_SL g3638 ( 
.A(n_3357),
.Y(n_3638)
);

AOI22xp33_ASAP7_75t_L g3639 ( 
.A1(n_3368),
.A2(n_3181),
.B1(n_3176),
.B2(n_3076),
.Y(n_3639)
);

AOI22xp33_ASAP7_75t_SL g3640 ( 
.A1(n_3448),
.A2(n_3009),
.B1(n_3178),
.B2(n_3181),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3275),
.Y(n_3641)
);

CKINVDCx5p33_ASAP7_75t_R g3642 ( 
.A(n_3276),
.Y(n_3642)
);

AOI22xp33_ASAP7_75t_SL g3643 ( 
.A1(n_3525),
.A2(n_3178),
.B1(n_3227),
.B2(n_3076),
.Y(n_3643)
);

OAI21xp5_ASAP7_75t_SL g3644 ( 
.A1(n_3407),
.A2(n_2831),
.B(n_3015),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3282),
.Y(n_3645)
);

AOI22xp33_ASAP7_75t_L g3646 ( 
.A1(n_3389),
.A2(n_3140),
.B1(n_3149),
.B2(n_3206),
.Y(n_3646)
);

BUFx2_ASAP7_75t_L g3647 ( 
.A(n_3437),
.Y(n_3647)
);

AOI22xp33_ASAP7_75t_L g3648 ( 
.A1(n_3323),
.A2(n_2977),
.B1(n_3121),
.B2(n_2968),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3292),
.Y(n_3649)
);

NOR2xp33_ASAP7_75t_L g3650 ( 
.A(n_3361),
.B(n_3057),
.Y(n_3650)
);

OAI22xp5_ASAP7_75t_L g3651 ( 
.A1(n_3294),
.A2(n_3034),
.B1(n_3015),
.B2(n_3125),
.Y(n_3651)
);

AOI22xp33_ASAP7_75t_L g3652 ( 
.A1(n_3449),
.A2(n_3055),
.B1(n_3085),
.B2(n_3071),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3600),
.B(n_2900),
.Y(n_3653)
);

AOI22xp33_ASAP7_75t_SL g3654 ( 
.A1(n_3538),
.A2(n_3034),
.B1(n_3192),
.B2(n_3130),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_L g3655 ( 
.A(n_3336),
.B(n_3057),
.Y(n_3655)
);

AOI22xp33_ASAP7_75t_L g3656 ( 
.A1(n_3302),
.A2(n_3087),
.B1(n_3098),
.B2(n_3093),
.Y(n_3656)
);

OAI21xp5_ASAP7_75t_SL g3657 ( 
.A1(n_3265),
.A2(n_3130),
.B(n_3125),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3280),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_3574),
.B(n_2912),
.Y(n_3659)
);

BUFx12f_ASAP7_75t_L g3660 ( 
.A(n_3263),
.Y(n_3660)
);

AOI222xp33_ASAP7_75t_L g3661 ( 
.A1(n_3316),
.A2(n_3073),
.B1(n_3017),
.B2(n_2988),
.C1(n_3058),
.C2(n_3044),
.Y(n_3661)
);

HB1xp67_ASAP7_75t_L g3662 ( 
.A(n_3535),
.Y(n_3662)
);

NOR2xp33_ASAP7_75t_L g3663 ( 
.A(n_3385),
.B(n_2859),
.Y(n_3663)
);

AOI22xp33_ASAP7_75t_L g3664 ( 
.A1(n_3359),
.A2(n_3188),
.B1(n_3218),
.B2(n_2881),
.Y(n_3664)
);

AOI22xp33_ASAP7_75t_L g3665 ( 
.A1(n_3394),
.A2(n_3102),
.B1(n_3118),
.B2(n_3020),
.Y(n_3665)
);

AOI22xp33_ASAP7_75t_L g3666 ( 
.A1(n_3295),
.A2(n_3073),
.B1(n_3035),
.B2(n_3031),
.Y(n_3666)
);

AOI22xp33_ASAP7_75t_L g3667 ( 
.A1(n_3296),
.A2(n_2971),
.B1(n_3208),
.B2(n_3207),
.Y(n_3667)
);

OAI22xp5_ASAP7_75t_L g3668 ( 
.A1(n_3335),
.A2(n_3171),
.B1(n_2946),
.B2(n_2902),
.Y(n_3668)
);

NOR2xp33_ASAP7_75t_L g3669 ( 
.A(n_3435),
.B(n_3172),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3427),
.B(n_2912),
.Y(n_3670)
);

OAI21xp5_ASAP7_75t_SL g3671 ( 
.A1(n_3352),
.A2(n_3171),
.B(n_2946),
.Y(n_3671)
);

BUFx3_ASAP7_75t_L g3672 ( 
.A(n_3325),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3299),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3300),
.Y(n_3674)
);

AOI22xp33_ASAP7_75t_L g3675 ( 
.A1(n_3546),
.A2(n_2964),
.B1(n_2941),
.B2(n_3100),
.Y(n_3675)
);

AOI22xp5_ASAP7_75t_L g3676 ( 
.A1(n_3281),
.A2(n_3187),
.B1(n_3204),
.B2(n_3100),
.Y(n_3676)
);

OAI22xp5_ASAP7_75t_L g3677 ( 
.A1(n_3289),
.A2(n_2902),
.B1(n_3225),
.B2(n_3043),
.Y(n_3677)
);

BUFx4f_ASAP7_75t_SL g3678 ( 
.A(n_3360),
.Y(n_3678)
);

OAI21xp33_ASAP7_75t_L g3679 ( 
.A1(n_3510),
.A2(n_2649),
.B(n_2941),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_3286),
.Y(n_3680)
);

BUFx8_ASAP7_75t_L g3681 ( 
.A(n_3305),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3427),
.B(n_3187),
.Y(n_3682)
);

BUFx12f_ASAP7_75t_L g3683 ( 
.A(n_3244),
.Y(n_3683)
);

INVx2_ASAP7_75t_SL g3684 ( 
.A(n_3262),
.Y(n_3684)
);

OAI22xp5_ASAP7_75t_L g3685 ( 
.A1(n_3308),
.A2(n_3225),
.B1(n_3043),
.B2(n_2945),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3307),
.Y(n_3686)
);

OAI22xp5_ASAP7_75t_L g3687 ( 
.A1(n_3261),
.A2(n_3561),
.B1(n_3253),
.B2(n_3284),
.Y(n_3687)
);

AOI22xp33_ASAP7_75t_L g3688 ( 
.A1(n_3259),
.A2(n_3392),
.B1(n_3475),
.B2(n_3401),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3314),
.Y(n_3689)
);

OAI22xp33_ASAP7_75t_SL g3690 ( 
.A1(n_3419),
.A2(n_2945),
.B1(n_2944),
.B2(n_3204),
.Y(n_3690)
);

BUFx5_ASAP7_75t_L g3691 ( 
.A(n_3467),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3531),
.B(n_3026),
.Y(n_3692)
);

OAI21xp5_ASAP7_75t_L g3693 ( 
.A1(n_3486),
.A2(n_3029),
.B(n_2990),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3315),
.Y(n_3694)
);

NOR2xp33_ASAP7_75t_L g3695 ( 
.A(n_3495),
.B(n_2889),
.Y(n_3695)
);

INVx3_ASAP7_75t_L g3696 ( 
.A(n_3490),
.Y(n_3696)
);

AOI22xp33_ASAP7_75t_SL g3697 ( 
.A1(n_3539),
.A2(n_3077),
.B1(n_3079),
.B2(n_3001),
.Y(n_3697)
);

AOI22xp33_ASAP7_75t_SL g3698 ( 
.A1(n_3539),
.A2(n_3142),
.B1(n_3131),
.B2(n_2935),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3304),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_SL g3700 ( 
.A(n_3311),
.B(n_2935),
.Y(n_3700)
);

OAI22xp33_ASAP7_75t_L g3701 ( 
.A1(n_3370),
.A2(n_3078),
.B1(n_3029),
.B2(n_2842),
.Y(n_3701)
);

OAI22xp33_ASAP7_75t_L g3702 ( 
.A1(n_3257),
.A2(n_3078),
.B1(n_2860),
.B2(n_2937),
.Y(n_3702)
);

OAI21xp5_ASAP7_75t_SL g3703 ( 
.A1(n_3452),
.A2(n_2830),
.B(n_2878),
.Y(n_3703)
);

AOI22xp33_ASAP7_75t_SL g3704 ( 
.A1(n_3558),
.A2(n_3142),
.B1(n_3131),
.B2(n_3141),
.Y(n_3704)
);

AOI22xp33_ASAP7_75t_L g3705 ( 
.A1(n_3338),
.A2(n_2882),
.B1(n_2937),
.B2(n_2860),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3321),
.Y(n_3706)
);

INVx3_ASAP7_75t_L g3707 ( 
.A(n_3490),
.Y(n_3707)
);

OAI21xp5_ASAP7_75t_SL g3708 ( 
.A1(n_3366),
.A2(n_2830),
.B(n_2878),
.Y(n_3708)
);

OAI21xp5_ASAP7_75t_SL g3709 ( 
.A1(n_3372),
.A2(n_3354),
.B(n_3318),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3327),
.Y(n_3710)
);

OAI222xp33_ASAP7_75t_L g3711 ( 
.A1(n_3363),
.A2(n_2944),
.B1(n_2882),
.B2(n_3112),
.C1(n_3069),
.C2(n_3163),
.Y(n_3711)
);

AOI22xp33_ASAP7_75t_SL g3712 ( 
.A1(n_3558),
.A2(n_3141),
.B1(n_2935),
.B2(n_3163),
.Y(n_3712)
);

INVx4_ASAP7_75t_L g3713 ( 
.A(n_3447),
.Y(n_3713)
);

OAI21xp5_ASAP7_75t_SL g3714 ( 
.A1(n_3374),
.A2(n_2879),
.B(n_2877),
.Y(n_3714)
);

OAI22xp33_ASAP7_75t_L g3715 ( 
.A1(n_3248),
.A2(n_2983),
.B1(n_3136),
.B2(n_2879),
.Y(n_3715)
);

AOI22xp33_ASAP7_75t_SL g3716 ( 
.A1(n_3362),
.A2(n_2935),
.B1(n_3141),
.B2(n_2983),
.Y(n_3716)
);

BUFx4f_ASAP7_75t_SL g3717 ( 
.A(n_3331),
.Y(n_3717)
);

HB1xp67_ASAP7_75t_L g3718 ( 
.A(n_3496),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3328),
.Y(n_3719)
);

OAI22xp5_ASAP7_75t_L g3720 ( 
.A1(n_3285),
.A2(n_3112),
.B1(n_3069),
.B2(n_3045),
.Y(n_3720)
);

INVx1_ASAP7_75t_SL g3721 ( 
.A(n_3511),
.Y(n_3721)
);

AOI22xp33_ASAP7_75t_L g3722 ( 
.A1(n_3379),
.A2(n_2877),
.B1(n_3059),
.B2(n_3045),
.Y(n_3722)
);

OAI22xp5_ASAP7_75t_L g3723 ( 
.A1(n_3334),
.A2(n_3062),
.B1(n_3066),
.B2(n_3059),
.Y(n_3723)
);

AOI22xp33_ASAP7_75t_L g3724 ( 
.A1(n_3513),
.A2(n_3066),
.B1(n_3113),
.B2(n_3062),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3337),
.Y(n_3725)
);

AOI22xp33_ASAP7_75t_L g3726 ( 
.A1(n_3330),
.A2(n_3113),
.B1(n_3157),
.B2(n_3148),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3340),
.Y(n_3727)
);

AOI22xp33_ASAP7_75t_L g3728 ( 
.A1(n_3483),
.A2(n_3157),
.B1(n_3205),
.B2(n_3148),
.Y(n_3728)
);

OAI21xp5_ASAP7_75t_SL g3729 ( 
.A1(n_3278),
.A2(n_3212),
.B(n_3205),
.Y(n_3729)
);

OAI22xp5_ASAP7_75t_L g3730 ( 
.A1(n_3333),
.A2(n_3251),
.B1(n_3572),
.B2(n_3541),
.Y(n_3730)
);

BUFx5_ASAP7_75t_L g3731 ( 
.A(n_3467),
.Y(n_3731)
);

BUFx3_ASAP7_75t_L g3732 ( 
.A(n_3287),
.Y(n_3732)
);

OAI22xp5_ASAP7_75t_L g3733 ( 
.A1(n_3380),
.A2(n_3212),
.B1(n_3213),
.B2(n_3210),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_3317),
.Y(n_3734)
);

AND2x4_ASAP7_75t_L g3735 ( 
.A(n_3241),
.B(n_3242),
.Y(n_3735)
);

AOI22xp33_ASAP7_75t_SL g3736 ( 
.A1(n_3409),
.A2(n_3567),
.B1(n_3566),
.B2(n_3527),
.Y(n_3736)
);

AOI22xp33_ASAP7_75t_L g3737 ( 
.A1(n_3563),
.A2(n_3213),
.B1(n_3013),
.B2(n_3018),
.Y(n_3737)
);

AND2x2_ASAP7_75t_L g3738 ( 
.A(n_3453),
.B(n_280),
.Y(n_3738)
);

AOI22xp33_ASAP7_75t_L g3739 ( 
.A1(n_3575),
.A2(n_3214),
.B1(n_3202),
.B2(n_3210),
.Y(n_3739)
);

CKINVDCx20_ASAP7_75t_R g3740 ( 
.A(n_3277),
.Y(n_3740)
);

AOI22xp33_ASAP7_75t_L g3741 ( 
.A1(n_3582),
.A2(n_3141),
.B1(n_2935),
.B2(n_2367),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3341),
.Y(n_3742)
);

OAI21xp5_ASAP7_75t_SL g3743 ( 
.A1(n_3386),
.A2(n_3119),
.B(n_2787),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3417),
.Y(n_3744)
);

AOI22xp33_ASAP7_75t_L g3745 ( 
.A1(n_3349),
.A2(n_3509),
.B1(n_3505),
.B2(n_3543),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3344),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3346),
.Y(n_3747)
);

BUFx6f_ASAP7_75t_L g3748 ( 
.A(n_3393),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3353),
.Y(n_3749)
);

AOI22xp33_ASAP7_75t_L g3750 ( 
.A1(n_3565),
.A2(n_3141),
.B1(n_2391),
.B2(n_2433),
.Y(n_3750)
);

OAI22xp33_ASAP7_75t_L g3751 ( 
.A1(n_3447),
.A2(n_2999),
.B1(n_3094),
.B2(n_3086),
.Y(n_3751)
);

INVx2_ASAP7_75t_L g3752 ( 
.A(n_3425),
.Y(n_3752)
);

OAI22xp5_ASAP7_75t_L g3753 ( 
.A1(n_3383),
.A2(n_3160),
.B1(n_3216),
.B2(n_3104),
.Y(n_3753)
);

BUFx6f_ASAP7_75t_L g3754 ( 
.A(n_3393),
.Y(n_3754)
);

AOI22xp33_ASAP7_75t_L g3755 ( 
.A1(n_3584),
.A2(n_2391),
.B1(n_2433),
.B2(n_2386),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3356),
.Y(n_3756)
);

BUFx4f_ASAP7_75t_SL g3757 ( 
.A(n_3290),
.Y(n_3757)
);

AOI22xp33_ASAP7_75t_L g3758 ( 
.A1(n_3591),
.A2(n_2450),
.B1(n_2438),
.B2(n_2730),
.Y(n_3758)
);

AOI22xp33_ASAP7_75t_L g3759 ( 
.A1(n_3594),
.A2(n_3441),
.B1(n_3446),
.B2(n_3279),
.Y(n_3759)
);

OR2x2_ASAP7_75t_L g3760 ( 
.A(n_3523),
.B(n_3119),
.Y(n_3760)
);

BUFx2_ASAP7_75t_L g3761 ( 
.A(n_3536),
.Y(n_3761)
);

OAI22xp33_ASAP7_75t_L g3762 ( 
.A1(n_3402),
.A2(n_2999),
.B1(n_3094),
.B2(n_3086),
.Y(n_3762)
);

OAI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_3436),
.A2(n_3160),
.B1(n_3216),
.B2(n_3104),
.Y(n_3763)
);

OAI22xp5_ASAP7_75t_L g3764 ( 
.A1(n_3309),
.A2(n_3429),
.B1(n_3545),
.B2(n_3501),
.Y(n_3764)
);

AOI22xp33_ASAP7_75t_SL g3765 ( 
.A1(n_3566),
.A2(n_3567),
.B1(n_3526),
.B2(n_3242),
.Y(n_3765)
);

AOI22xp33_ASAP7_75t_SL g3766 ( 
.A1(n_3241),
.A2(n_3083),
.B1(n_2950),
.B2(n_3104),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3364),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3476),
.Y(n_3768)
);

AOI22xp33_ASAP7_75t_L g3769 ( 
.A1(n_3455),
.A2(n_2450),
.B1(n_2438),
.B2(n_2730),
.Y(n_3769)
);

AOI22xp5_ASAP7_75t_L g3770 ( 
.A1(n_3429),
.A2(n_2378),
.B1(n_2381),
.B2(n_2380),
.Y(n_3770)
);

AOI22xp33_ASAP7_75t_SL g3771 ( 
.A1(n_3252),
.A2(n_3293),
.B1(n_3599),
.B2(n_3414),
.Y(n_3771)
);

AOI22xp33_ASAP7_75t_L g3772 ( 
.A1(n_3471),
.A2(n_2569),
.B1(n_2559),
.B2(n_2692),
.Y(n_3772)
);

AOI22xp33_ASAP7_75t_L g3773 ( 
.A1(n_3507),
.A2(n_2569),
.B1(n_2559),
.B2(n_2692),
.Y(n_3773)
);

BUFx3_ASAP7_75t_L g3774 ( 
.A(n_3367),
.Y(n_3774)
);

BUFx8_ASAP7_75t_SL g3775 ( 
.A(n_3324),
.Y(n_3775)
);

CKINVDCx8_ASAP7_75t_R g3776 ( 
.A(n_3268),
.Y(n_3776)
);

AOI22xp33_ASAP7_75t_SL g3777 ( 
.A1(n_3252),
.A2(n_3083),
.B1(n_3160),
.B2(n_3104),
.Y(n_3777)
);

AOI22xp33_ASAP7_75t_L g3778 ( 
.A1(n_3355),
.A2(n_2692),
.B1(n_2524),
.B2(n_2604),
.Y(n_3778)
);

OAI22xp5_ASAP7_75t_L g3779 ( 
.A1(n_3388),
.A2(n_3216),
.B1(n_3160),
.B2(n_3086),
.Y(n_3779)
);

INVx3_ASAP7_75t_L g3780 ( 
.A(n_3497),
.Y(n_3780)
);

AOI22xp33_ASAP7_75t_L g3781 ( 
.A1(n_3508),
.A2(n_2524),
.B1(n_2604),
.B2(n_2587),
.Y(n_3781)
);

AOI22xp33_ASAP7_75t_SL g3782 ( 
.A1(n_3293),
.A2(n_3216),
.B1(n_3094),
.B2(n_3096),
.Y(n_3782)
);

BUFx2_ASAP7_75t_L g3783 ( 
.A(n_3477),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3365),
.Y(n_3784)
);

AOI22xp5_ASAP7_75t_L g3785 ( 
.A1(n_3498),
.A2(n_3096),
.B1(n_2999),
.B2(n_2787),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3369),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3376),
.Y(n_3787)
);

OAI22xp5_ASAP7_75t_L g3788 ( 
.A1(n_3246),
.A2(n_3096),
.B1(n_2794),
.B2(n_2298),
.Y(n_3788)
);

BUFx3_ASAP7_75t_L g3789 ( 
.A(n_3375),
.Y(n_3789)
);

AOI22xp33_ASAP7_75t_SL g3790 ( 
.A1(n_3412),
.A2(n_2812),
.B1(n_2847),
.B2(n_2843),
.Y(n_3790)
);

NOR2xp33_ASAP7_75t_L g3791 ( 
.A(n_3592),
.B(n_3445),
.Y(n_3791)
);

INVx5_ASAP7_75t_L g3792 ( 
.A(n_3412),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3381),
.Y(n_3793)
);

OAI22xp5_ASAP7_75t_L g3794 ( 
.A1(n_3246),
.A2(n_2794),
.B1(n_2524),
.B2(n_2604),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3382),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3411),
.Y(n_3796)
);

CKINVDCx5p33_ASAP7_75t_R g3797 ( 
.A(n_3378),
.Y(n_3797)
);

OAI21xp5_ASAP7_75t_SL g3798 ( 
.A1(n_3588),
.A2(n_2843),
.B(n_2812),
.Y(n_3798)
);

AND2x2_ASAP7_75t_L g3799 ( 
.A(n_3595),
.B(n_280),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3413),
.Y(n_3800)
);

OAI22xp5_ASAP7_75t_L g3801 ( 
.A1(n_3391),
.A2(n_2587),
.B1(n_3003),
.B2(n_2987),
.Y(n_3801)
);

AOI22xp33_ASAP7_75t_SL g3802 ( 
.A1(n_3390),
.A2(n_2843),
.B1(n_2847),
.B2(n_2812),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3415),
.B(n_2987),
.Y(n_3803)
);

HB1xp67_ASAP7_75t_L g3804 ( 
.A(n_3598),
.Y(n_3804)
);

BUFx4f_ASAP7_75t_SL g3805 ( 
.A(n_3312),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3560),
.B(n_283),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3416),
.Y(n_3807)
);

AOI22xp33_ASAP7_75t_SL g3808 ( 
.A1(n_3390),
.A2(n_2873),
.B1(n_2926),
.B2(n_2847),
.Y(n_3808)
);

AOI22xp33_ASAP7_75t_L g3809 ( 
.A1(n_3438),
.A2(n_2587),
.B1(n_2718),
.B2(n_2699),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3488),
.Y(n_3810)
);

AOI22xp33_ASAP7_75t_L g3811 ( 
.A1(n_3504),
.A2(n_2723),
.B1(n_3003),
.B2(n_2987),
.Y(n_3811)
);

AOI22xp33_ASAP7_75t_L g3812 ( 
.A1(n_3524),
.A2(n_3007),
.B1(n_3012),
.B2(n_3003),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3418),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3432),
.Y(n_3814)
);

OAI22xp5_ASAP7_75t_L g3815 ( 
.A1(n_3557),
.A2(n_3012),
.B1(n_3040),
.B2(n_3007),
.Y(n_3815)
);

INVx3_ASAP7_75t_L g3816 ( 
.A(n_3497),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_SL g3817 ( 
.A(n_3343),
.B(n_2873),
.Y(n_3817)
);

OAI22xp5_ASAP7_75t_L g3818 ( 
.A1(n_3387),
.A2(n_3012),
.B1(n_3040),
.B2(n_3007),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3432),
.Y(n_3819)
);

AOI22xp33_ASAP7_75t_L g3820 ( 
.A1(n_3457),
.A2(n_3492),
.B1(n_3555),
.B2(n_3396),
.Y(n_3820)
);

AOI22xp33_ASAP7_75t_L g3821 ( 
.A1(n_3549),
.A2(n_3052),
.B1(n_3106),
.B2(n_3040),
.Y(n_3821)
);

AOI22xp33_ASAP7_75t_L g3822 ( 
.A1(n_3551),
.A2(n_3106),
.B1(n_3122),
.B2(n_3052),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3462),
.Y(n_3823)
);

AOI22xp33_ASAP7_75t_L g3824 ( 
.A1(n_3329),
.A2(n_3106),
.B1(n_3122),
.B2(n_3052),
.Y(n_3824)
);

INVx3_ASAP7_75t_L g3825 ( 
.A(n_3520),
.Y(n_3825)
);

INVx1_ASAP7_75t_SL g3826 ( 
.A(n_3571),
.Y(n_3826)
);

CKINVDCx5p33_ASAP7_75t_R g3827 ( 
.A(n_3306),
.Y(n_3827)
);

AOI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3421),
.A2(n_3128),
.B1(n_3155),
.B2(n_3122),
.Y(n_3828)
);

OAI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3550),
.A2(n_2309),
.B(n_283),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3462),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3464),
.Y(n_3831)
);

OAI22xp5_ASAP7_75t_L g3832 ( 
.A1(n_3400),
.A2(n_3155),
.B1(n_3165),
.B2(n_3128),
.Y(n_3832)
);

AOI22xp33_ASAP7_75t_SL g3833 ( 
.A1(n_3520),
.A2(n_2926),
.B1(n_2975),
.B2(n_2873),
.Y(n_3833)
);

INVxp67_ASAP7_75t_L g3834 ( 
.A(n_3484),
.Y(n_3834)
);

AOI22xp33_ASAP7_75t_SL g3835 ( 
.A1(n_3343),
.A2(n_2975),
.B1(n_2978),
.B2(n_2926),
.Y(n_3835)
);

OAI21xp5_ASAP7_75t_SL g3836 ( 
.A1(n_3310),
.A2(n_2978),
.B(n_2975),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_3578),
.B(n_284),
.Y(n_3837)
);

HB1xp67_ASAP7_75t_L g3838 ( 
.A(n_3431),
.Y(n_3838)
);

AND2x2_ASAP7_75t_L g3839 ( 
.A(n_3593),
.B(n_285),
.Y(n_3839)
);

AOI222xp33_ASAP7_75t_L g3840 ( 
.A1(n_3260),
.A2(n_288),
.B1(n_291),
.B2(n_286),
.C1(n_287),
.C2(n_290),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3464),
.Y(n_3841)
);

AND2x2_ASAP7_75t_L g3842 ( 
.A(n_3562),
.B(n_3371),
.Y(n_3842)
);

CKINVDCx14_ASAP7_75t_R g3843 ( 
.A(n_3297),
.Y(n_3843)
);

AOI22xp33_ASAP7_75t_SL g3844 ( 
.A1(n_3348),
.A2(n_2978),
.B1(n_3155),
.B2(n_3128),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3487),
.Y(n_3845)
);

BUFx3_ASAP7_75t_L g3846 ( 
.A(n_3377),
.Y(n_3846)
);

AOI22xp33_ASAP7_75t_L g3847 ( 
.A1(n_3421),
.A2(n_3168),
.B1(n_3196),
.B2(n_3165),
.Y(n_3847)
);

NOR2x1_ASAP7_75t_R g3848 ( 
.A(n_3544),
.B(n_3548),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3489),
.Y(n_3849)
);

OAI22xp5_ASAP7_75t_L g3850 ( 
.A1(n_3470),
.A2(n_3422),
.B1(n_3585),
.B2(n_3439),
.Y(n_3850)
);

OAI222xp33_ASAP7_75t_L g3851 ( 
.A1(n_3350),
.A2(n_290),
.B1(n_292),
.B2(n_287),
.C1(n_288),
.C2(n_291),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3384),
.B(n_3165),
.Y(n_3852)
);

AOI22xp33_ASAP7_75t_L g3853 ( 
.A1(n_3298),
.A2(n_3196),
.B1(n_3211),
.B2(n_3168),
.Y(n_3853)
);

INVx3_ASAP7_75t_L g3854 ( 
.A(n_3478),
.Y(n_3854)
);

AOI222xp33_ASAP7_75t_L g3855 ( 
.A1(n_3267),
.A2(n_3503),
.B1(n_3434),
.B2(n_3313),
.C1(n_3479),
.C2(n_3458),
.Y(n_3855)
);

OAI21xp5_ASAP7_75t_SL g3856 ( 
.A1(n_3348),
.A2(n_3196),
.B(n_3168),
.Y(n_3856)
);

BUFx3_ASAP7_75t_L g3857 ( 
.A(n_3420),
.Y(n_3857)
);

AOI22xp33_ASAP7_75t_L g3858 ( 
.A1(n_3556),
.A2(n_3220),
.B1(n_3223),
.B2(n_3211),
.Y(n_3858)
);

OAI21xp5_ASAP7_75t_SL g3859 ( 
.A1(n_3444),
.A2(n_3540),
.B(n_3532),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3522),
.Y(n_3860)
);

OAI21xp5_ASAP7_75t_SL g3861 ( 
.A1(n_3444),
.A2(n_3220),
.B(n_3211),
.Y(n_3861)
);

AOI22xp33_ASAP7_75t_L g3862 ( 
.A1(n_3564),
.A2(n_3223),
.B1(n_3220),
.B2(n_3229),
.Y(n_3862)
);

OAI21xp33_ASAP7_75t_L g3863 ( 
.A1(n_3547),
.A2(n_3223),
.B(n_3229),
.Y(n_3863)
);

OAI21xp5_ASAP7_75t_SL g3864 ( 
.A1(n_3532),
.A2(n_3231),
.B(n_3229),
.Y(n_3864)
);

AOI22xp33_ASAP7_75t_SL g3865 ( 
.A1(n_3540),
.A2(n_3237),
.B1(n_3231),
.B2(n_294),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3395),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3405),
.B(n_292),
.Y(n_3867)
);

NOR3xp33_ASAP7_75t_L g3868 ( 
.A(n_3589),
.B(n_293),
.C(n_295),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_3258),
.Y(n_3869)
);

OAI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_3568),
.A2(n_293),
.B(n_296),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3406),
.Y(n_3871)
);

NOR2xp33_ASAP7_75t_L g3872 ( 
.A(n_3580),
.B(n_296),
.Y(n_3872)
);

AOI22xp33_ASAP7_75t_L g3873 ( 
.A1(n_3576),
.A2(n_3237),
.B1(n_3231),
.B2(n_299),
.Y(n_3873)
);

AOI22xp33_ASAP7_75t_L g3874 ( 
.A1(n_3576),
.A2(n_3237),
.B1(n_299),
.B2(n_297),
.Y(n_3874)
);

BUFx2_ASAP7_75t_L g3875 ( 
.A(n_3502),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3403),
.Y(n_3876)
);

BUFx3_ASAP7_75t_L g3877 ( 
.A(n_3428),
.Y(n_3877)
);

HB1xp67_ASAP7_75t_L g3878 ( 
.A(n_3408),
.Y(n_3878)
);

OAI22xp5_ASAP7_75t_L g3879 ( 
.A1(n_3423),
.A2(n_300),
.B1(n_297),
.B2(n_298),
.Y(n_3879)
);

AOI22xp5_ASAP7_75t_L g3880 ( 
.A1(n_3423),
.A2(n_301),
.B1(n_298),
.B2(n_300),
.Y(n_3880)
);

NOR2xp33_ASAP7_75t_L g3881 ( 
.A(n_3440),
.B(n_302),
.Y(n_3881)
);

BUFx4f_ASAP7_75t_SL g3882 ( 
.A(n_3326),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3410),
.Y(n_3883)
);

OAI22xp5_ASAP7_75t_L g3884 ( 
.A1(n_3439),
.A2(n_306),
.B1(n_303),
.B2(n_304),
.Y(n_3884)
);

OAI22xp5_ASAP7_75t_L g3885 ( 
.A1(n_3451),
.A2(n_3482),
.B1(n_3517),
.B2(n_3430),
.Y(n_3885)
);

AOI22xp33_ASAP7_75t_SL g3886 ( 
.A1(n_3517),
.A2(n_307),
.B1(n_303),
.B2(n_304),
.Y(n_3886)
);

AOI22xp33_ASAP7_75t_L g3887 ( 
.A1(n_3424),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_3887)
);

HB1xp67_ASAP7_75t_L g3888 ( 
.A(n_3465),
.Y(n_3888)
);

AOI22xp33_ASAP7_75t_SL g3889 ( 
.A1(n_3451),
.A2(n_311),
.B1(n_308),
.B2(n_310),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3466),
.Y(n_3890)
);

OAI22xp5_ASAP7_75t_L g3891 ( 
.A1(n_3482),
.A2(n_315),
.B1(n_312),
.B2(n_314),
.Y(n_3891)
);

BUFx12f_ASAP7_75t_L g3892 ( 
.A(n_3267),
.Y(n_3892)
);

OAI21xp5_ASAP7_75t_SL g3893 ( 
.A1(n_3345),
.A2(n_312),
.B(n_314),
.Y(n_3893)
);

NAND2xp33_ASAP7_75t_SL g3894 ( 
.A(n_3713),
.B(n_3433),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_3602),
.B(n_3468),
.Y(n_3895)
);

AOI22xp33_ASAP7_75t_L g3896 ( 
.A1(n_3613),
.A2(n_3399),
.B1(n_3332),
.B2(n_3319),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3878),
.Y(n_3897)
);

HB1xp67_ASAP7_75t_L g3898 ( 
.A(n_3603),
.Y(n_3898)
);

OAI222xp33_ASAP7_75t_L g3899 ( 
.A1(n_3764),
.A2(n_3601),
.B1(n_3736),
.B2(n_3611),
.C1(n_3651),
.C2(n_3771),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3838),
.B(n_3469),
.Y(n_3900)
);

OAI222xp33_ASAP7_75t_L g3901 ( 
.A1(n_3617),
.A2(n_3456),
.B1(n_3473),
.B2(n_3426),
.C1(n_3430),
.C2(n_3472),
.Y(n_3901)
);

OAI22xp5_ASAP7_75t_L g3902 ( 
.A1(n_3619),
.A2(n_3573),
.B1(n_3373),
.B2(n_3430),
.Y(n_3902)
);

AOI22xp33_ASAP7_75t_L g3903 ( 
.A1(n_3621),
.A2(n_3569),
.B1(n_3579),
.B2(n_3373),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3845),
.B(n_3500),
.Y(n_3904)
);

AOI22xp33_ASAP7_75t_L g3905 ( 
.A1(n_3621),
.A2(n_3579),
.B1(n_3485),
.B2(n_3514),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3888),
.Y(n_3906)
);

AOI22xp33_ASAP7_75t_L g3907 ( 
.A1(n_3661),
.A2(n_3485),
.B1(n_3514),
.B2(n_3581),
.Y(n_3907)
);

AOI22xp33_ASAP7_75t_L g3908 ( 
.A1(n_3688),
.A2(n_3529),
.B1(n_3516),
.B2(n_3426),
.Y(n_3908)
);

AOI22xp5_ASAP7_75t_L g3909 ( 
.A1(n_3685),
.A2(n_3459),
.B1(n_3262),
.B2(n_3291),
.Y(n_3909)
);

AOI22xp33_ASAP7_75t_SL g3910 ( 
.A1(n_3668),
.A2(n_3291),
.B1(n_3502),
.B2(n_3426),
.Y(n_3910)
);

AND2x2_ASAP7_75t_L g3911 ( 
.A(n_3659),
.B(n_3512),
.Y(n_3911)
);

AND2x2_ASAP7_75t_L g3912 ( 
.A(n_3842),
.B(n_3625),
.Y(n_3912)
);

AOI22xp33_ASAP7_75t_L g3913 ( 
.A1(n_3840),
.A2(n_3529),
.B1(n_3518),
.B2(n_3519),
.Y(n_3913)
);

AOI22xp33_ASAP7_75t_L g3914 ( 
.A1(n_3730),
.A2(n_3530),
.B1(n_3534),
.B2(n_3515),
.Y(n_3914)
);

AOI22xp33_ASAP7_75t_L g3915 ( 
.A1(n_3677),
.A2(n_3656),
.B1(n_3868),
.B2(n_3701),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3866),
.B(n_3537),
.Y(n_3916)
);

AOI22xp33_ASAP7_75t_L g3917 ( 
.A1(n_3648),
.A2(n_3474),
.B1(n_3461),
.B2(n_3552),
.Y(n_3917)
);

INVx2_ASAP7_75t_L g3918 ( 
.A(n_3658),
.Y(n_3918)
);

AOI22xp33_ASAP7_75t_L g3919 ( 
.A1(n_3759),
.A2(n_3587),
.B1(n_3597),
.B2(n_3358),
.Y(n_3919)
);

OAI22xp5_ASAP7_75t_L g3920 ( 
.A1(n_3628),
.A2(n_3342),
.B1(n_3590),
.B2(n_3243),
.Y(n_3920)
);

AND2x2_ASAP7_75t_L g3921 ( 
.A(n_3718),
.B(n_3583),
.Y(n_3921)
);

AOI22xp33_ASAP7_75t_L g3922 ( 
.A1(n_3630),
.A2(n_3478),
.B1(n_3493),
.B2(n_3481),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3876),
.B(n_3478),
.Y(n_3923)
);

AOI22xp33_ASAP7_75t_L g3924 ( 
.A1(n_3675),
.A2(n_3481),
.B1(n_3528),
.B2(n_3493),
.Y(n_3924)
);

AOI22xp33_ASAP7_75t_L g3925 ( 
.A1(n_3652),
.A2(n_3481),
.B1(n_3528),
.B2(n_3493),
.Y(n_3925)
);

BUFx2_ASAP7_75t_L g3926 ( 
.A(n_3696),
.Y(n_3926)
);

AOI22xp5_ASAP7_75t_L g3927 ( 
.A1(n_3893),
.A2(n_3586),
.B1(n_3521),
.B2(n_3404),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3883),
.B(n_3528),
.Y(n_3928)
);

AOI22xp33_ASAP7_75t_L g3929 ( 
.A1(n_3664),
.A2(n_3553),
.B1(n_3506),
.B2(n_3596),
.Y(n_3929)
);

AOI22xp33_ASAP7_75t_L g3930 ( 
.A1(n_3702),
.A2(n_3646),
.B1(n_3679),
.B2(n_3665),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3804),
.B(n_3692),
.Y(n_3931)
);

AOI22xp33_ASAP7_75t_L g3932 ( 
.A1(n_3889),
.A2(n_3553),
.B1(n_3463),
.B2(n_3347),
.Y(n_3932)
);

AND2x2_ASAP7_75t_L g3933 ( 
.A(n_3620),
.B(n_3662),
.Y(n_3933)
);

AND2x2_ASAP7_75t_L g3934 ( 
.A(n_3604),
.B(n_3583),
.Y(n_3934)
);

OAI221xp5_ASAP7_75t_SL g3935 ( 
.A1(n_3644),
.A2(n_3671),
.B1(n_3657),
.B2(n_3709),
.C(n_3636),
.Y(n_3935)
);

AOI22xp33_ASAP7_75t_SL g3936 ( 
.A1(n_3850),
.A2(n_3553),
.B1(n_3542),
.B2(n_3499),
.Y(n_3936)
);

AOI22xp33_ASAP7_75t_L g3937 ( 
.A1(n_3829),
.A2(n_3577),
.B1(n_3442),
.B2(n_3351),
.Y(n_3937)
);

AOI22xp33_ASAP7_75t_L g3938 ( 
.A1(n_3639),
.A2(n_3577),
.B1(n_3450),
.B2(n_3454),
.Y(n_3938)
);

AOI22xp33_ASAP7_75t_L g3939 ( 
.A1(n_3886),
.A2(n_3454),
.B1(n_3266),
.B2(n_318),
.Y(n_3939)
);

AOI22xp33_ASAP7_75t_L g3940 ( 
.A1(n_3715),
.A2(n_318),
.B1(n_315),
.B2(n_317),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3890),
.B(n_317),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3606),
.B(n_319),
.Y(n_3942)
);

AOI222xp33_ASAP7_75t_L g3943 ( 
.A1(n_3875),
.A2(n_3655),
.B1(n_3650),
.B2(n_3881),
.C1(n_3683),
.C2(n_3666),
.Y(n_3943)
);

OAI222xp33_ASAP7_75t_L g3944 ( 
.A1(n_3640),
.A2(n_321),
.B1(n_323),
.B2(n_319),
.C1(n_320),
.C2(n_322),
.Y(n_3944)
);

OAI22xp33_ASAP7_75t_SL g3945 ( 
.A1(n_3647),
.A2(n_323),
.B1(n_320),
.B2(n_321),
.Y(n_3945)
);

AOI22xp33_ASAP7_75t_L g3946 ( 
.A1(n_3820),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_3946)
);

AOI22xp33_ASAP7_75t_L g3947 ( 
.A1(n_3693),
.A2(n_327),
.B1(n_324),
.B2(n_325),
.Y(n_3947)
);

AOI22xp33_ASAP7_75t_SL g3948 ( 
.A1(n_3633),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_3948)
);

NOR3xp33_ASAP7_75t_L g3949 ( 
.A(n_3851),
.B(n_329),
.C(n_330),
.Y(n_3949)
);

AOI22xp33_ASAP7_75t_SL g3950 ( 
.A1(n_3687),
.A2(n_333),
.B1(n_330),
.B2(n_332),
.Y(n_3950)
);

AOI22xp33_ASAP7_75t_L g3951 ( 
.A1(n_3705),
.A2(n_337),
.B1(n_334),
.B2(n_336),
.Y(n_3951)
);

AOI222xp33_ASAP7_75t_L g3952 ( 
.A1(n_3667),
.A2(n_338),
.B1(n_340),
.B2(n_334),
.C1(n_336),
.C2(n_339),
.Y(n_3952)
);

AOI22xp33_ASAP7_75t_L g3953 ( 
.A1(n_3870),
.A2(n_341),
.B1(n_338),
.B2(n_340),
.Y(n_3953)
);

AOI22xp33_ASAP7_75t_L g3954 ( 
.A1(n_3879),
.A2(n_343),
.B1(n_341),
.B2(n_342),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3635),
.Y(n_3955)
);

OAI221xp5_ASAP7_75t_L g3956 ( 
.A1(n_3627),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.C(n_345),
.Y(n_3956)
);

AOI22xp33_ASAP7_75t_SL g3957 ( 
.A1(n_3690),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_3957)
);

AOI22xp33_ASAP7_75t_SL g3958 ( 
.A1(n_3691),
.A2(n_349),
.B1(n_346),
.B2(n_348),
.Y(n_3958)
);

AOI22xp33_ASAP7_75t_L g3959 ( 
.A1(n_3884),
.A2(n_3891),
.B1(n_3745),
.B2(n_3669),
.Y(n_3959)
);

AOI22xp33_ASAP7_75t_L g3960 ( 
.A1(n_3654),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3641),
.Y(n_3961)
);

AND2x2_ASAP7_75t_L g3962 ( 
.A(n_3614),
.B(n_350),
.Y(n_3962)
);

AOI22xp33_ASAP7_75t_L g3963 ( 
.A1(n_3663),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_3963)
);

AOI22xp33_ASAP7_75t_L g3964 ( 
.A1(n_3728),
.A2(n_3880),
.B1(n_3738),
.B2(n_3872),
.Y(n_3964)
);

OAI22xp5_ASAP7_75t_L g3965 ( 
.A1(n_3722),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_3615),
.B(n_356),
.Y(n_3966)
);

AOI22xp5_ASAP7_75t_L g3967 ( 
.A1(n_3676),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_3967)
);

INVx2_ASAP7_75t_L g3968 ( 
.A(n_3680),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3622),
.B(n_3634),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_3645),
.Y(n_3970)
);

AOI22xp33_ASAP7_75t_SL g3971 ( 
.A1(n_3691),
.A2(n_362),
.B1(n_359),
.B2(n_360),
.Y(n_3971)
);

OAI221xp5_ASAP7_75t_L g3972 ( 
.A1(n_3637),
.A2(n_365),
.B1(n_362),
.B2(n_364),
.C(n_366),
.Y(n_3972)
);

AOI22xp33_ASAP7_75t_L g3973 ( 
.A1(n_3880),
.A2(n_367),
.B1(n_364),
.B2(n_366),
.Y(n_3973)
);

OAI22xp33_ASAP7_75t_L g3974 ( 
.A1(n_3792),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_3974)
);

AOI22xp33_ASAP7_75t_SL g3975 ( 
.A1(n_3691),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_3975)
);

AOI22xp5_ASAP7_75t_L g3976 ( 
.A1(n_3676),
.A2(n_3714),
.B1(n_3703),
.B2(n_3708),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3649),
.B(n_370),
.Y(n_3977)
);

AOI22xp33_ASAP7_75t_SL g3978 ( 
.A1(n_3691),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.Y(n_3978)
);

INVx3_ASAP7_75t_L g3979 ( 
.A(n_3696),
.Y(n_3979)
);

OAI222xp33_ASAP7_75t_L g3980 ( 
.A1(n_3643),
.A2(n_375),
.B1(n_377),
.B2(n_373),
.C1(n_374),
.C2(n_376),
.Y(n_3980)
);

AOI22xp33_ASAP7_75t_L g3981 ( 
.A1(n_3865),
.A2(n_377),
.B1(n_374),
.B2(n_375),
.Y(n_3981)
);

AOI22xp33_ASAP7_75t_L g3982 ( 
.A1(n_3887),
.A2(n_381),
.B1(n_378),
.B2(n_379),
.Y(n_3982)
);

NAND3xp33_ASAP7_75t_SL g3983 ( 
.A(n_3740),
.B(n_378),
.C(n_379),
.Y(n_3983)
);

OAI221xp5_ASAP7_75t_SL g3984 ( 
.A1(n_3632),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.C(n_385),
.Y(n_3984)
);

OAI221xp5_ASAP7_75t_L g3985 ( 
.A1(n_3726),
.A2(n_385),
.B1(n_382),
.B2(n_383),
.C(n_386),
.Y(n_3985)
);

OAI211xp5_ASAP7_75t_L g3986 ( 
.A1(n_3697),
.A2(n_388),
.B(n_386),
.C(n_387),
.Y(n_3986)
);

AOI22xp33_ASAP7_75t_L g3987 ( 
.A1(n_3629),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_3987)
);

AOI22xp33_ASAP7_75t_L g3988 ( 
.A1(n_3839),
.A2(n_391),
.B1(n_389),
.B2(n_390),
.Y(n_3988)
);

AND2x2_ASAP7_75t_L g3989 ( 
.A(n_3673),
.B(n_391),
.Y(n_3989)
);

AOI22xp33_ASAP7_75t_L g3990 ( 
.A1(n_3806),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_3990)
);

OAI22xp5_ASAP7_75t_L g3991 ( 
.A1(n_3765),
.A2(n_398),
.B1(n_395),
.B2(n_396),
.Y(n_3991)
);

AOI22xp5_ASAP7_75t_L g3992 ( 
.A1(n_3773),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3674),
.B(n_399),
.Y(n_3993)
);

AOI22xp33_ASAP7_75t_L g3994 ( 
.A1(n_3837),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_3994)
);

AOI22xp33_ASAP7_75t_L g3995 ( 
.A1(n_3799),
.A2(n_3772),
.B1(n_3713),
.B2(n_3781),
.Y(n_3995)
);

AOI22xp33_ASAP7_75t_L g3996 ( 
.A1(n_3874),
.A2(n_406),
.B1(n_403),
.B2(n_404),
.Y(n_3996)
);

OAI222xp33_ASAP7_75t_L g3997 ( 
.A1(n_3716),
.A2(n_408),
.B1(n_410),
.B2(n_404),
.C1(n_406),
.C2(n_409),
.Y(n_3997)
);

AOI22xp33_ASAP7_75t_L g3998 ( 
.A1(n_3769),
.A2(n_3867),
.B1(n_3700),
.B2(n_3791),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_3686),
.B(n_409),
.Y(n_3999)
);

AOI22xp33_ASAP7_75t_L g4000 ( 
.A1(n_3735),
.A2(n_413),
.B1(n_411),
.B2(n_412),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3689),
.B(n_411),
.Y(n_4001)
);

OAI21xp5_ASAP7_75t_SL g4002 ( 
.A1(n_3843),
.A2(n_412),
.B(n_413),
.Y(n_4002)
);

AOI221xp5_ASAP7_75t_L g4003 ( 
.A1(n_3694),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.C(n_417),
.Y(n_4003)
);

BUFx6f_ASAP7_75t_L g4004 ( 
.A(n_3623),
.Y(n_4004)
);

AOI22xp33_ASAP7_75t_L g4005 ( 
.A1(n_3735),
.A2(n_418),
.B1(n_414),
.B2(n_417),
.Y(n_4005)
);

AND2x2_ASAP7_75t_L g4006 ( 
.A(n_3706),
.B(n_418),
.Y(n_4006)
);

AOI222xp33_ASAP7_75t_L g4007 ( 
.A1(n_3610),
.A2(n_422),
.B1(n_425),
.B2(n_419),
.C1(n_420),
.C2(n_423),
.Y(n_4007)
);

AOI22xp33_ASAP7_75t_L g4008 ( 
.A1(n_3682),
.A2(n_422),
.B1(n_419),
.B2(n_420),
.Y(n_4008)
);

OAI22xp33_ASAP7_75t_SL g4009 ( 
.A1(n_3834),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.Y(n_4009)
);

AND2x2_ASAP7_75t_L g4010 ( 
.A(n_3710),
.B(n_426),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3719),
.B(n_428),
.Y(n_4011)
);

AOI22xp33_ASAP7_75t_SL g4012 ( 
.A1(n_3691),
.A2(n_430),
.B1(n_428),
.B2(n_429),
.Y(n_4012)
);

OAI222xp33_ASAP7_75t_L g4013 ( 
.A1(n_3792),
.A2(n_432),
.B1(n_434),
.B2(n_430),
.C1(n_431),
.C2(n_433),
.Y(n_4013)
);

AOI22xp33_ASAP7_75t_L g4014 ( 
.A1(n_3723),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_4014)
);

AOI22xp33_ASAP7_75t_L g4015 ( 
.A1(n_3761),
.A2(n_438),
.B1(n_434),
.B2(n_436),
.Y(n_4015)
);

OAI22xp5_ASAP7_75t_L g4016 ( 
.A1(n_3792),
.A2(n_439),
.B1(n_436),
.B2(n_438),
.Y(n_4016)
);

AOI221xp5_ASAP7_75t_L g4017 ( 
.A1(n_3725),
.A2(n_442),
.B1(n_439),
.B2(n_441),
.C(n_443),
.Y(n_4017)
);

AOI22xp33_ASAP7_75t_L g4018 ( 
.A1(n_3720),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_4018)
);

OAI22xp5_ASAP7_75t_L g4019 ( 
.A1(n_3724),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.Y(n_4019)
);

AOI22xp33_ASAP7_75t_L g4020 ( 
.A1(n_3783),
.A2(n_449),
.B1(n_446),
.B2(n_448),
.Y(n_4020)
);

OAI22xp33_ASAP7_75t_L g4021 ( 
.A1(n_3608),
.A2(n_451),
.B1(n_448),
.B2(n_450),
.Y(n_4021)
);

AOI22xp33_ASAP7_75t_L g4022 ( 
.A1(n_3811),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.Y(n_4022)
);

AOI22xp33_ASAP7_75t_L g4023 ( 
.A1(n_3695),
.A2(n_455),
.B1(n_452),
.B2(n_453),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3727),
.B(n_453),
.Y(n_4024)
);

AOI22xp33_ASAP7_75t_L g4025 ( 
.A1(n_3814),
.A2(n_459),
.B1(n_456),
.B2(n_458),
.Y(n_4025)
);

OAI22xp33_ASAP7_75t_L g4026 ( 
.A1(n_3608),
.A2(n_461),
.B1(n_459),
.B2(n_460),
.Y(n_4026)
);

AOI22xp33_ASAP7_75t_L g4027 ( 
.A1(n_3819),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_4027)
);

AOI22xp33_ASAP7_75t_L g4028 ( 
.A1(n_3823),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3742),
.Y(n_4029)
);

AOI22xp33_ASAP7_75t_L g4030 ( 
.A1(n_3830),
.A2(n_3841),
.B1(n_3831),
.B2(n_3778),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3746),
.B(n_463),
.Y(n_4031)
);

AOI22xp33_ASAP7_75t_L g4032 ( 
.A1(n_3707),
.A2(n_468),
.B1(n_465),
.B2(n_466),
.Y(n_4032)
);

OAI22xp5_ASAP7_75t_L g4033 ( 
.A1(n_3698),
.A2(n_471),
.B1(n_465),
.B2(n_470),
.Y(n_4033)
);

AOI22xp33_ASAP7_75t_L g4034 ( 
.A1(n_3707),
.A2(n_474),
.B1(n_471),
.B2(n_472),
.Y(n_4034)
);

AOI22xp33_ASAP7_75t_L g4035 ( 
.A1(n_3780),
.A2(n_475),
.B1(n_472),
.B2(n_474),
.Y(n_4035)
);

NAND3xp33_ASAP7_75t_L g4036 ( 
.A(n_3859),
.B(n_475),
.C(n_477),
.Y(n_4036)
);

AOI22xp33_ASAP7_75t_L g4037 ( 
.A1(n_3780),
.A2(n_479),
.B1(n_477),
.B2(n_478),
.Y(n_4037)
);

AOI22xp33_ASAP7_75t_L g4038 ( 
.A1(n_3816),
.A2(n_3825),
.B1(n_3809),
.B2(n_3672),
.Y(n_4038)
);

NAND3xp33_ASAP7_75t_L g4039 ( 
.A(n_3737),
.B(n_479),
.C(n_480),
.Y(n_4039)
);

AOI222xp33_ASAP7_75t_L g4040 ( 
.A1(n_3624),
.A2(n_480),
.B1(n_481),
.B2(n_482),
.C1(n_483),
.C2(n_484),
.Y(n_4040)
);

INVx2_ASAP7_75t_L g4041 ( 
.A(n_3699),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_3747),
.B(n_481),
.Y(n_4042)
);

OAI22xp5_ASAP7_75t_L g4043 ( 
.A1(n_3704),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.Y(n_4043)
);

AOI22xp33_ASAP7_75t_SL g4044 ( 
.A1(n_3731),
.A2(n_487),
.B1(n_485),
.B2(n_486),
.Y(n_4044)
);

OAI22xp5_ASAP7_75t_L g4045 ( 
.A1(n_3712),
.A2(n_487),
.B1(n_485),
.B2(n_486),
.Y(n_4045)
);

AOI22xp33_ASAP7_75t_SL g4046 ( 
.A1(n_3731),
.A2(n_491),
.B1(n_488),
.B2(n_489),
.Y(n_4046)
);

OAI22xp5_ASAP7_75t_L g4047 ( 
.A1(n_3739),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.Y(n_4047)
);

AOI22xp33_ASAP7_75t_L g4048 ( 
.A1(n_3816),
.A2(n_496),
.B1(n_492),
.B2(n_495),
.Y(n_4048)
);

AOI22xp33_ASAP7_75t_SL g4049 ( 
.A1(n_3731),
.A2(n_498),
.B1(n_496),
.B2(n_497),
.Y(n_4049)
);

OAI22xp33_ASAP7_75t_L g4050 ( 
.A1(n_3608),
.A2(n_3618),
.B1(n_3825),
.B2(n_3678),
.Y(n_4050)
);

AOI22xp33_ASAP7_75t_SL g4051 ( 
.A1(n_3731),
.A2(n_499),
.B1(n_497),
.B2(n_498),
.Y(n_4051)
);

AOI22xp33_ASAP7_75t_L g4052 ( 
.A1(n_3774),
.A2(n_502),
.B1(n_499),
.B2(n_501),
.Y(n_4052)
);

BUFx2_ASAP7_75t_L g4053 ( 
.A(n_3618),
.Y(n_4053)
);

AOI22xp33_ASAP7_75t_L g4054 ( 
.A1(n_3789),
.A2(n_505),
.B1(n_503),
.B2(n_504),
.Y(n_4054)
);

AOI22xp33_ASAP7_75t_L g4055 ( 
.A1(n_3846),
.A2(n_506),
.B1(n_503),
.B2(n_504),
.Y(n_4055)
);

AOI22xp33_ASAP7_75t_L g4056 ( 
.A1(n_3857),
.A2(n_508),
.B1(n_506),
.B2(n_507),
.Y(n_4056)
);

OAI22xp5_ASAP7_75t_L g4057 ( 
.A1(n_3873),
.A2(n_510),
.B1(n_507),
.B2(n_509),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_3749),
.B(n_511),
.Y(n_4058)
);

AOI22xp33_ASAP7_75t_L g4059 ( 
.A1(n_3877),
.A2(n_513),
.B1(n_511),
.B2(n_512),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3756),
.B(n_512),
.Y(n_4060)
);

NAND3xp33_ASAP7_75t_L g4061 ( 
.A(n_3821),
.B(n_513),
.C(n_514),
.Y(n_4061)
);

OAI222xp33_ASAP7_75t_L g4062 ( 
.A1(n_3776),
.A2(n_515),
.B1(n_516),
.B2(n_517),
.C1(n_518),
.C2(n_519),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3767),
.Y(n_4063)
);

AOI22xp33_ASAP7_75t_L g4064 ( 
.A1(n_3670),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_4064)
);

AOI22xp33_ASAP7_75t_L g4065 ( 
.A1(n_3733),
.A2(n_521),
.B1(n_519),
.B2(n_520),
.Y(n_4065)
);

OR2x2_ASAP7_75t_L g4066 ( 
.A(n_3607),
.B(n_520),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3784),
.B(n_521),
.Y(n_4067)
);

AOI22xp33_ASAP7_75t_L g4068 ( 
.A1(n_3786),
.A2(n_3793),
.B1(n_3795),
.B2(n_3787),
.Y(n_4068)
);

AOI22xp33_ASAP7_75t_L g4069 ( 
.A1(n_3796),
.A2(n_524),
.B1(n_522),
.B2(n_523),
.Y(n_4069)
);

AOI22xp33_ASAP7_75t_L g4070 ( 
.A1(n_3800),
.A2(n_524),
.B1(n_522),
.B2(n_523),
.Y(n_4070)
);

AOI22xp33_ASAP7_75t_L g4071 ( 
.A1(n_3807),
.A2(n_528),
.B1(n_525),
.B2(n_526),
.Y(n_4071)
);

OAI21xp33_ASAP7_75t_SL g4072 ( 
.A1(n_3862),
.A2(n_525),
.B(n_526),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_3813),
.B(n_530),
.Y(n_4073)
);

AOI22xp33_ASAP7_75t_L g4074 ( 
.A1(n_3731),
.A2(n_532),
.B1(n_530),
.B2(n_531),
.Y(n_4074)
);

OA21x2_ASAP7_75t_L g4075 ( 
.A1(n_3863),
.A2(n_531),
.B(n_532),
.Y(n_4075)
);

AOI22xp33_ASAP7_75t_L g4076 ( 
.A1(n_3653),
.A2(n_3684),
.B1(n_3618),
.B2(n_3721),
.Y(n_4076)
);

OAI22xp5_ASAP7_75t_L g4077 ( 
.A1(n_3812),
.A2(n_537),
.B1(n_533),
.B2(n_535),
.Y(n_4077)
);

AOI22xp33_ASAP7_75t_L g4078 ( 
.A1(n_3626),
.A2(n_540),
.B1(n_538),
.B2(n_539),
.Y(n_4078)
);

OAI22xp5_ASAP7_75t_L g4079 ( 
.A1(n_3782),
.A2(n_541),
.B1(n_539),
.B2(n_540),
.Y(n_4079)
);

NAND3xp33_ASAP7_75t_L g4080 ( 
.A(n_3824),
.B(n_3760),
.C(n_3743),
.Y(n_4080)
);

OA21x2_ASAP7_75t_L g4081 ( 
.A1(n_3863),
.A2(n_3711),
.B(n_3798),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3734),
.B(n_542),
.Y(n_4082)
);

AOI22xp5_ASAP7_75t_L g4083 ( 
.A1(n_3885),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_4083)
);

OAI22xp5_ASAP7_75t_L g4084 ( 
.A1(n_3790),
.A2(n_547),
.B1(n_545),
.B2(n_546),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3897),
.B(n_3869),
.Y(n_4085)
);

OAI22xp5_ASAP7_75t_L g4086 ( 
.A1(n_3935),
.A2(n_3853),
.B1(n_3785),
.B2(n_3847),
.Y(n_4086)
);

AND2x2_ASAP7_75t_L g4087 ( 
.A(n_3931),
.B(n_3871),
.Y(n_4087)
);

NAND3xp33_ASAP7_75t_L g4088 ( 
.A(n_3896),
.B(n_3855),
.C(n_3836),
.Y(n_4088)
);

OAI221xp5_ASAP7_75t_L g4089 ( 
.A1(n_4002),
.A2(n_3826),
.B1(n_3729),
.B2(n_3828),
.C(n_3642),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3906),
.B(n_3616),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_SL g4091 ( 
.A(n_3910),
.B(n_3835),
.Y(n_4091)
);

OAI21xp5_ASAP7_75t_L g4092 ( 
.A1(n_3957),
.A2(n_3808),
.B(n_3802),
.Y(n_4092)
);

AND2x2_ASAP7_75t_L g4093 ( 
.A(n_3912),
.B(n_3631),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_4068),
.B(n_3744),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_3933),
.B(n_3752),
.Y(n_4095)
);

AND2x2_ASAP7_75t_L g4096 ( 
.A(n_3911),
.B(n_3768),
.Y(n_4096)
);

AOI22xp33_ASAP7_75t_L g4097 ( 
.A1(n_3949),
.A2(n_3815),
.B1(n_3832),
.B2(n_3818),
.Y(n_4097)
);

NAND3xp33_ASAP7_75t_L g4098 ( 
.A(n_3943),
.B(n_3822),
.C(n_3785),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3898),
.B(n_3900),
.Y(n_4099)
);

NAND3xp33_ASAP7_75t_L g4100 ( 
.A(n_3957),
.B(n_3861),
.C(n_3856),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_3955),
.B(n_3810),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_SL g4102 ( 
.A(n_3910),
.B(n_3844),
.Y(n_4102)
);

OA21x2_ASAP7_75t_L g4103 ( 
.A1(n_3976),
.A2(n_3864),
.B(n_3803),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3961),
.B(n_3849),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_L g4105 ( 
.A(n_3970),
.B(n_3860),
.Y(n_4105)
);

NAND3xp33_ASAP7_75t_L g4106 ( 
.A(n_3950),
.B(n_3858),
.C(n_3788),
.Y(n_4106)
);

OAI221xp5_ASAP7_75t_SL g4107 ( 
.A1(n_3915),
.A2(n_3762),
.B1(n_3758),
.B2(n_3751),
.C(n_3755),
.Y(n_4107)
);

AND2x2_ASAP7_75t_L g4108 ( 
.A(n_3895),
.B(n_3854),
.Y(n_4108)
);

AND2x2_ASAP7_75t_SL g4109 ( 
.A(n_3926),
.B(n_3623),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_4029),
.B(n_3852),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_4063),
.B(n_3770),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_SL g4112 ( 
.A(n_4050),
.B(n_3894),
.Y(n_4112)
);

AND2x2_ASAP7_75t_L g4113 ( 
.A(n_3921),
.B(n_3854),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_3904),
.B(n_3770),
.Y(n_4114)
);

AND2x2_ASAP7_75t_L g4115 ( 
.A(n_3934),
.B(n_3623),
.Y(n_4115)
);

OAI221xp5_ASAP7_75t_L g4116 ( 
.A1(n_3936),
.A2(n_3827),
.B1(n_3732),
.B2(n_3777),
.C(n_3766),
.Y(n_4116)
);

NOR2xp33_ASAP7_75t_R g4117 ( 
.A(n_4053),
.B(n_3609),
.Y(n_4117)
);

AND2x2_ASAP7_75t_L g4118 ( 
.A(n_3918),
.B(n_3748),
.Y(n_4118)
);

AOI22xp5_ASAP7_75t_L g4119 ( 
.A1(n_3913),
.A2(n_3892),
.B1(n_3779),
.B2(n_3763),
.Y(n_4119)
);

OAI21xp5_ASAP7_75t_SL g4120 ( 
.A1(n_3899),
.A2(n_3833),
.B(n_3753),
.Y(n_4120)
);

OA21x2_ASAP7_75t_L g4121 ( 
.A1(n_4080),
.A2(n_3817),
.B(n_3741),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_3969),
.B(n_3801),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_3968),
.B(n_3748),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_3914),
.B(n_3748),
.Y(n_4124)
);

NAND3xp33_ASAP7_75t_L g4125 ( 
.A(n_3950),
.B(n_3750),
.C(n_3794),
.Y(n_4125)
);

HB1xp67_ASAP7_75t_L g4126 ( 
.A(n_3979),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_3916),
.B(n_3754),
.Y(n_4127)
);

OAI22xp5_ASAP7_75t_L g4128 ( 
.A1(n_3937),
.A2(n_3638),
.B1(n_3882),
.B2(n_3805),
.Y(n_4128)
);

OAI21xp5_ASAP7_75t_SL g4129 ( 
.A1(n_3927),
.A2(n_3754),
.B(n_3612),
.Y(n_4129)
);

AND2x2_ASAP7_75t_L g4130 ( 
.A(n_4041),
.B(n_3754),
.Y(n_4130)
);

OAI22xp5_ASAP7_75t_L g4131 ( 
.A1(n_3907),
.A2(n_3757),
.B1(n_3717),
.B2(n_3660),
.Y(n_4131)
);

NAND3xp33_ASAP7_75t_L g4132 ( 
.A(n_3948),
.B(n_3930),
.C(n_3958),
.Y(n_4132)
);

AND2x2_ASAP7_75t_L g4133 ( 
.A(n_3979),
.B(n_546),
.Y(n_4133)
);

AND2x2_ASAP7_75t_L g4134 ( 
.A(n_4076),
.B(n_3923),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_3928),
.B(n_548),
.Y(n_4135)
);

AOI21xp33_ASAP7_75t_L g4136 ( 
.A1(n_3920),
.A2(n_3848),
.B(n_548),
.Y(n_4136)
);

NAND3xp33_ASAP7_75t_L g4137 ( 
.A(n_3948),
.B(n_3681),
.C(n_3797),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3962),
.B(n_549),
.Y(n_4138)
);

NOR3xp33_ASAP7_75t_L g4139 ( 
.A(n_3983),
.B(n_3681),
.C(n_3605),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3966),
.B(n_549),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_3989),
.B(n_550),
.Y(n_4141)
);

OAI21xp5_ASAP7_75t_SL g4142 ( 
.A1(n_3909),
.A2(n_3775),
.B(n_550),
.Y(n_4142)
);

OAI21xp5_ASAP7_75t_SL g4143 ( 
.A1(n_4062),
.A2(n_551),
.B(n_552),
.Y(n_4143)
);

HB1xp67_ASAP7_75t_L g4144 ( 
.A(n_4004),
.Y(n_4144)
);

AND2x2_ASAP7_75t_L g4145 ( 
.A(n_3998),
.B(n_551),
.Y(n_4145)
);

AOI221xp5_ASAP7_75t_L g4146 ( 
.A1(n_3945),
.A2(n_552),
.B1(n_553),
.B2(n_554),
.C(n_555),
.Y(n_4146)
);

OAI22xp5_ASAP7_75t_L g4147 ( 
.A1(n_3964),
.A2(n_556),
.B1(n_554),
.B2(n_555),
.Y(n_4147)
);

OAI21xp5_ASAP7_75t_SL g4148 ( 
.A1(n_3932),
.A2(n_557),
.B(n_558),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_4006),
.B(n_559),
.Y(n_4149)
);

NAND3xp33_ASAP7_75t_L g4150 ( 
.A(n_3958),
.B(n_560),
.C(n_561),
.Y(n_4150)
);

NOR3xp33_ASAP7_75t_L g4151 ( 
.A(n_3944),
.B(n_560),
.C(n_561),
.Y(n_4151)
);

NAND3xp33_ASAP7_75t_L g4152 ( 
.A(n_3971),
.B(n_564),
.C(n_565),
.Y(n_4152)
);

OAI21x1_ASAP7_75t_L g4153 ( 
.A1(n_4075),
.A2(n_564),
.B(n_566),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_4010),
.B(n_566),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_4011),
.B(n_567),
.Y(n_4155)
);

AND2x2_ASAP7_75t_L g4156 ( 
.A(n_4030),
.B(n_567),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_4042),
.B(n_569),
.Y(n_4157)
);

NAND3xp33_ASAP7_75t_L g4158 ( 
.A(n_3971),
.B(n_570),
.C(n_571),
.Y(n_4158)
);

NAND3xp33_ASAP7_75t_L g4159 ( 
.A(n_3975),
.B(n_572),
.C(n_573),
.Y(n_4159)
);

NAND4xp25_ASAP7_75t_L g4160 ( 
.A(n_4007),
.B(n_574),
.C(n_572),
.D(n_573),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_SL g4161 ( 
.A(n_4038),
.B(n_575),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_4066),
.B(n_575),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_3995),
.B(n_576),
.Y(n_4163)
);

AND2x2_ASAP7_75t_L g4164 ( 
.A(n_3917),
.B(n_576),
.Y(n_4164)
);

AND2x2_ASAP7_75t_L g4165 ( 
.A(n_3938),
.B(n_3924),
.Y(n_4165)
);

OAI21xp33_ASAP7_75t_SL g4166 ( 
.A1(n_3922),
.A2(n_577),
.B(n_578),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_3942),
.B(n_580),
.Y(n_4167)
);

AOI22xp33_ASAP7_75t_SL g4168 ( 
.A1(n_4081),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.Y(n_4168)
);

INVx2_ASAP7_75t_L g4169 ( 
.A(n_4004),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_3977),
.B(n_581),
.Y(n_4170)
);

OAI21xp5_ASAP7_75t_SL g4171 ( 
.A1(n_3980),
.A2(n_582),
.B(n_583),
.Y(n_4171)
);

NOR2xp33_ASAP7_75t_L g4172 ( 
.A(n_3993),
.B(n_584),
.Y(n_4172)
);

AND2x2_ASAP7_75t_L g4173 ( 
.A(n_3903),
.B(n_585),
.Y(n_4173)
);

AND2x2_ASAP7_75t_L g4174 ( 
.A(n_4081),
.B(n_585),
.Y(n_4174)
);

NAND4xp25_ASAP7_75t_L g4175 ( 
.A(n_4040),
.B(n_587),
.C(n_588),
.D(n_589),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4101),
.Y(n_4176)
);

AND2x2_ASAP7_75t_L g4177 ( 
.A(n_4095),
.B(n_3908),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4104),
.Y(n_4178)
);

AND2x2_ASAP7_75t_L g4179 ( 
.A(n_4087),
.B(n_3925),
.Y(n_4179)
);

NOR3xp33_ASAP7_75t_L g4180 ( 
.A(n_4142),
.B(n_3997),
.C(n_4013),
.Y(n_4180)
);

BUFx3_ASAP7_75t_L g4181 ( 
.A(n_4108),
.Y(n_4181)
);

CKINVDCx5p33_ASAP7_75t_R g4182 ( 
.A(n_4117),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4085),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_4096),
.B(n_3999),
.Y(n_4184)
);

NAND3xp33_ASAP7_75t_L g4185 ( 
.A(n_4120),
.B(n_3978),
.C(n_3975),
.Y(n_4185)
);

NAND3xp33_ASAP7_75t_L g4186 ( 
.A(n_4120),
.B(n_4012),
.C(n_3978),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_L g4187 ( 
.A(n_4093),
.B(n_4001),
.Y(n_4187)
);

OA211x2_ASAP7_75t_L g4188 ( 
.A1(n_4112),
.A2(n_3905),
.B(n_4036),
.C(n_3939),
.Y(n_4188)
);

NAND3xp33_ASAP7_75t_L g4189 ( 
.A(n_4168),
.B(n_4044),
.C(n_4012),
.Y(n_4189)
);

NAND3xp33_ASAP7_75t_L g4190 ( 
.A(n_4174),
.B(n_4046),
.C(n_4044),
.Y(n_4190)
);

OA211x2_ASAP7_75t_L g4191 ( 
.A1(n_4091),
.A2(n_3929),
.B(n_3959),
.C(n_3940),
.Y(n_4191)
);

NAND2x1p5_ASAP7_75t_L g4192 ( 
.A(n_4133),
.B(n_4004),
.Y(n_4192)
);

NAND4xp75_ASAP7_75t_L g4193 ( 
.A(n_4102),
.B(n_4075),
.C(n_4072),
.D(n_4083),
.Y(n_4193)
);

NAND3xp33_ASAP7_75t_L g4194 ( 
.A(n_4132),
.B(n_4098),
.C(n_4088),
.Y(n_4194)
);

AOI22xp5_ASAP7_75t_SL g4195 ( 
.A1(n_4128),
.A2(n_4009),
.B1(n_3902),
.B2(n_3991),
.Y(n_4195)
);

NAND3xp33_ASAP7_75t_L g4196 ( 
.A(n_4142),
.B(n_4049),
.C(n_4046),
.Y(n_4196)
);

AOI22xp33_ASAP7_75t_L g4197 ( 
.A1(n_4151),
.A2(n_3956),
.B1(n_4051),
.B2(n_4049),
.Y(n_4197)
);

AND2x2_ASAP7_75t_L g4198 ( 
.A(n_4113),
.B(n_4004),
.Y(n_4198)
);

HB1xp67_ASAP7_75t_L g4199 ( 
.A(n_4126),
.Y(n_4199)
);

OR2x2_ASAP7_75t_L g4200 ( 
.A(n_4099),
.B(n_4024),
.Y(n_4200)
);

AOI22x1_ASAP7_75t_L g4201 ( 
.A1(n_4092),
.A2(n_3952),
.B1(n_4051),
.B2(n_3901),
.Y(n_4201)
);

AND2x2_ASAP7_75t_L g4202 ( 
.A(n_4115),
.B(n_3919),
.Y(n_4202)
);

INVx5_ASAP7_75t_L g4203 ( 
.A(n_4169),
.Y(n_4203)
);

NAND3xp33_ASAP7_75t_L g4204 ( 
.A(n_4143),
.B(n_4148),
.C(n_4171),
.Y(n_4204)
);

INVx2_ASAP7_75t_SL g4205 ( 
.A(n_4109),
.Y(n_4205)
);

AND2x2_ASAP7_75t_L g4206 ( 
.A(n_4134),
.B(n_4031),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_4118),
.B(n_4058),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4090),
.Y(n_4208)
);

NAND4xp75_ASAP7_75t_L g4209 ( 
.A(n_4136),
.B(n_3967),
.C(n_4067),
.D(n_4060),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_4094),
.B(n_4073),
.Y(n_4210)
);

OAI21xp5_ASAP7_75t_L g4211 ( 
.A1(n_4143),
.A2(n_3986),
.B(n_4039),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_4114),
.B(n_3941),
.Y(n_4212)
);

NAND3xp33_ASAP7_75t_L g4213 ( 
.A(n_4148),
.B(n_3987),
.C(n_3984),
.Y(n_4213)
);

BUFx3_ASAP7_75t_L g4214 ( 
.A(n_4123),
.Y(n_4214)
);

OR2x2_ASAP7_75t_L g4215 ( 
.A(n_4110),
.B(n_4082),
.Y(n_4215)
);

NOR3xp33_ASAP7_75t_L g4216 ( 
.A(n_4137),
.B(n_3974),
.C(n_3972),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_4122),
.B(n_4018),
.Y(n_4217)
);

NAND3xp33_ASAP7_75t_L g4218 ( 
.A(n_4171),
.B(n_4061),
.C(n_4016),
.Y(n_4218)
);

OA211x2_ASAP7_75t_L g4219 ( 
.A1(n_4100),
.A2(n_3960),
.B(n_3953),
.C(n_3981),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4111),
.B(n_3947),
.Y(n_4220)
);

AO21x2_ASAP7_75t_L g4221 ( 
.A1(n_4153),
.A2(n_4161),
.B(n_4124),
.Y(n_4221)
);

INVx2_ASAP7_75t_L g4222 ( 
.A(n_4130),
.Y(n_4222)
);

AO21x2_ASAP7_75t_L g4223 ( 
.A1(n_4162),
.A2(n_3992),
.B(n_4021),
.Y(n_4223)
);

OR2x2_ASAP7_75t_L g4224 ( 
.A(n_4105),
.B(n_4077),
.Y(n_4224)
);

AND2x2_ASAP7_75t_L g4225 ( 
.A(n_4165),
.B(n_4065),
.Y(n_4225)
);

NAND3xp33_ASAP7_75t_L g4226 ( 
.A(n_4116),
.B(n_3946),
.C(n_4014),
.Y(n_4226)
);

AND2x2_ASAP7_75t_L g4227 ( 
.A(n_4144),
.B(n_4103),
.Y(n_4227)
);

AO21x2_ASAP7_75t_L g4228 ( 
.A1(n_4139),
.A2(n_4170),
.B(n_4167),
.Y(n_4228)
);

NOR2xp33_ASAP7_75t_L g4229 ( 
.A(n_4129),
.B(n_3985),
.Y(n_4229)
);

NAND4xp75_ASAP7_75t_L g4230 ( 
.A(n_4119),
.B(n_4017),
.C(n_4003),
.D(n_4045),
.Y(n_4230)
);

NAND3xp33_ASAP7_75t_L g4231 ( 
.A(n_4103),
.B(n_3973),
.C(n_4033),
.Y(n_4231)
);

AO21x2_ASAP7_75t_L g4232 ( 
.A1(n_4173),
.A2(n_4026),
.B(n_3965),
.Y(n_4232)
);

OR2x2_ASAP7_75t_L g4233 ( 
.A(n_4127),
.B(n_4019),
.Y(n_4233)
);

XOR2xp5_ASAP7_75t_L g4234 ( 
.A(n_4131),
.B(n_4079),
.Y(n_4234)
);

NAND4xp75_ASAP7_75t_L g4235 ( 
.A(n_4163),
.B(n_4084),
.C(n_4043),
.D(n_3988),
.Y(n_4235)
);

OR2x2_ASAP7_75t_L g4236 ( 
.A(n_4129),
.B(n_4047),
.Y(n_4236)
);

OA211x2_ASAP7_75t_L g4237 ( 
.A1(n_4097),
.A2(n_3990),
.B(n_3994),
.C(n_4000),
.Y(n_4237)
);

NAND4xp75_ASAP7_75t_L g4238 ( 
.A(n_4145),
.B(n_3963),
.C(n_4015),
.D(n_4078),
.Y(n_4238)
);

HB1xp67_ASAP7_75t_L g4239 ( 
.A(n_4121),
.Y(n_4239)
);

AO21x2_ASAP7_75t_L g4240 ( 
.A1(n_4156),
.A2(n_4057),
.B(n_4034),
.Y(n_4240)
);

AND2x2_ASAP7_75t_L g4241 ( 
.A(n_4121),
.B(n_4022),
.Y(n_4241)
);

AOI21x1_ASAP7_75t_L g4242 ( 
.A1(n_4086),
.A2(n_587),
.B(n_588),
.Y(n_4242)
);

AOI221xp5_ASAP7_75t_L g4243 ( 
.A1(n_4147),
.A2(n_4023),
.B1(n_4020),
.B2(n_4005),
.C(n_4055),
.Y(n_4243)
);

NOR3xp33_ASAP7_75t_L g4244 ( 
.A(n_4089),
.B(n_4054),
.C(n_4052),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4135),
.Y(n_4245)
);

INVx2_ASAP7_75t_SL g4246 ( 
.A(n_4181),
.Y(n_4246)
);

AND2x4_ASAP7_75t_L g4247 ( 
.A(n_4227),
.B(n_4106),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_4176),
.B(n_4164),
.Y(n_4248)
);

AND2x2_ASAP7_75t_L g4249 ( 
.A(n_4214),
.B(n_4138),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_4199),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4176),
.Y(n_4251)
);

XOR2xp5_ASAP7_75t_L g4252 ( 
.A(n_4182),
.B(n_4160),
.Y(n_4252)
);

NAND4xp75_ASAP7_75t_L g4253 ( 
.A(n_4191),
.B(n_4166),
.C(n_4141),
.D(n_4149),
.Y(n_4253)
);

NAND2x1_ASAP7_75t_L g4254 ( 
.A(n_4205),
.B(n_4150),
.Y(n_4254)
);

XNOR2x2_ASAP7_75t_L g4255 ( 
.A(n_4194),
.B(n_4160),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4178),
.Y(n_4256)
);

XOR2x2_ASAP7_75t_L g4257 ( 
.A(n_4204),
.B(n_4152),
.Y(n_4257)
);

XNOR2xp5_ASAP7_75t_L g4258 ( 
.A(n_4234),
.B(n_4175),
.Y(n_4258)
);

AND2x2_ASAP7_75t_L g4259 ( 
.A(n_4198),
.B(n_4140),
.Y(n_4259)
);

NAND4xp75_ASAP7_75t_L g4260 ( 
.A(n_4188),
.B(n_4154),
.C(n_4157),
.D(n_4155),
.Y(n_4260)
);

INVxp67_ASAP7_75t_L g4261 ( 
.A(n_4228),
.Y(n_4261)
);

NAND4xp75_ASAP7_75t_SL g4262 ( 
.A(n_4229),
.B(n_4172),
.C(n_4175),
.D(n_4107),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4178),
.Y(n_4263)
);

NOR2xp33_ASAP7_75t_L g4264 ( 
.A(n_4228),
.B(n_4125),
.Y(n_4264)
);

OR2x2_ASAP7_75t_L g4265 ( 
.A(n_4183),
.B(n_4158),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_4203),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_4208),
.B(n_4146),
.Y(n_4267)
);

XNOR2xp5_ASAP7_75t_L g4268 ( 
.A(n_4195),
.B(n_4159),
.Y(n_4268)
);

NAND4xp25_ASAP7_75t_L g4269 ( 
.A(n_4237),
.B(n_4219),
.C(n_4185),
.D(n_4186),
.Y(n_4269)
);

XOR2x2_ASAP7_75t_L g4270 ( 
.A(n_4196),
.B(n_4056),
.Y(n_4270)
);

XOR2x1_ASAP7_75t_L g4271 ( 
.A(n_4201),
.B(n_4032),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_4222),
.B(n_4035),
.Y(n_4272)
);

NOR2x1_ASAP7_75t_L g4273 ( 
.A(n_4190),
.B(n_4074),
.Y(n_4273)
);

AND2x2_ASAP7_75t_L g4274 ( 
.A(n_4179),
.B(n_4037),
.Y(n_4274)
);

AND2x2_ASAP7_75t_L g4275 ( 
.A(n_4177),
.B(n_4048),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_4210),
.B(n_4064),
.Y(n_4276)
);

XNOR2xp5_ASAP7_75t_L g4277 ( 
.A(n_4206),
.B(n_4059),
.Y(n_4277)
);

AND2x2_ASAP7_75t_L g4278 ( 
.A(n_4202),
.B(n_3954),
.Y(n_4278)
);

NOR3xp33_ASAP7_75t_SL g4279 ( 
.A(n_4226),
.B(n_590),
.C(n_591),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_L g4280 ( 
.A(n_4212),
.B(n_3951),
.Y(n_4280)
);

AND2x2_ASAP7_75t_L g4281 ( 
.A(n_4245),
.B(n_4025),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_SL g4282 ( 
.A(n_4239),
.B(n_4008),
.Y(n_4282)
);

NAND4xp75_ASAP7_75t_L g4283 ( 
.A(n_4241),
.B(n_4071),
.C(n_4070),
.D(n_4069),
.Y(n_4283)
);

INVx1_ASAP7_75t_SL g4284 ( 
.A(n_4203),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4215),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4245),
.B(n_4027),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_4200),
.B(n_4028),
.Y(n_4287)
);

AND2x2_ASAP7_75t_L g4288 ( 
.A(n_4207),
.B(n_3996),
.Y(n_4288)
);

INVx2_ASAP7_75t_SL g4289 ( 
.A(n_4203),
.Y(n_4289)
);

AND2x2_ASAP7_75t_L g4290 ( 
.A(n_4192),
.B(n_3982),
.Y(n_4290)
);

NAND4xp75_ASAP7_75t_L g4291 ( 
.A(n_4225),
.B(n_590),
.C(n_592),
.D(n_593),
.Y(n_4291)
);

INVx1_ASAP7_75t_SL g4292 ( 
.A(n_4236),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4184),
.Y(n_4293)
);

INVxp67_ASAP7_75t_L g4294 ( 
.A(n_4187),
.Y(n_4294)
);

NOR3xp33_ASAP7_75t_L g4295 ( 
.A(n_4242),
.B(n_592),
.C(n_593),
.Y(n_4295)
);

XNOR2x2_ASAP7_75t_L g4296 ( 
.A(n_4193),
.B(n_4189),
.Y(n_4296)
);

INVx1_ASAP7_75t_SL g4297 ( 
.A(n_4233),
.Y(n_4297)
);

OAI22xp5_ASAP7_75t_L g4298 ( 
.A1(n_4197),
.A2(n_594),
.B1(n_595),
.B2(n_596),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4224),
.Y(n_4299)
);

BUFx2_ASAP7_75t_L g4300 ( 
.A(n_4221),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4217),
.Y(n_4301)
);

NAND4xp75_ASAP7_75t_L g4302 ( 
.A(n_4211),
.B(n_594),
.C(n_595),
.D(n_596),
.Y(n_4302)
);

XNOR2xp5_ASAP7_75t_L g4303 ( 
.A(n_4238),
.B(n_597),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_4221),
.B(n_597),
.Y(n_4304)
);

AND2x2_ASAP7_75t_L g4305 ( 
.A(n_4216),
.B(n_598),
.Y(n_4305)
);

NAND4xp75_ASAP7_75t_SL g4306 ( 
.A(n_4180),
.B(n_598),
.C(n_599),
.D(n_600),
.Y(n_4306)
);

XOR2x2_ASAP7_75t_L g4307 ( 
.A(n_4235),
.B(n_600),
.Y(n_4307)
);

XOR2x2_ASAP7_75t_L g4308 ( 
.A(n_4296),
.B(n_4209),
.Y(n_4308)
);

XOR2x2_ASAP7_75t_L g4309 ( 
.A(n_4258),
.B(n_4255),
.Y(n_4309)
);

INVx1_ASAP7_75t_SL g4310 ( 
.A(n_4284),
.Y(n_4310)
);

INVx2_ASAP7_75t_L g4311 ( 
.A(n_4250),
.Y(n_4311)
);

INVx2_ASAP7_75t_L g4312 ( 
.A(n_4251),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4256),
.Y(n_4313)
);

HB1xp67_ASAP7_75t_L g4314 ( 
.A(n_4297),
.Y(n_4314)
);

XOR2x2_ASAP7_75t_L g4315 ( 
.A(n_4268),
.B(n_4213),
.Y(n_4315)
);

XOR2x2_ASAP7_75t_L g4316 ( 
.A(n_4262),
.B(n_4230),
.Y(n_4316)
);

XNOR2xp5_ASAP7_75t_L g4317 ( 
.A(n_4271),
.B(n_4244),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4263),
.Y(n_4318)
);

XNOR2x1_ASAP7_75t_L g4319 ( 
.A(n_4307),
.B(n_4218),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4299),
.Y(n_4320)
);

XOR2x2_ASAP7_75t_L g4321 ( 
.A(n_4252),
.B(n_4231),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4285),
.Y(n_4322)
);

BUFx3_ASAP7_75t_L g4323 ( 
.A(n_4246),
.Y(n_4323)
);

INVx2_ASAP7_75t_L g4324 ( 
.A(n_4284),
.Y(n_4324)
);

INVx1_ASAP7_75t_SL g4325 ( 
.A(n_4289),
.Y(n_4325)
);

INVx2_ASAP7_75t_L g4326 ( 
.A(n_4297),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4265),
.Y(n_4327)
);

XNOR2xp5_ASAP7_75t_L g4328 ( 
.A(n_4269),
.B(n_4220),
.Y(n_4328)
);

INVx2_ASAP7_75t_L g4329 ( 
.A(n_4304),
.Y(n_4329)
);

XNOR2xp5_ASAP7_75t_L g4330 ( 
.A(n_4269),
.B(n_4232),
.Y(n_4330)
);

AND2x2_ASAP7_75t_L g4331 ( 
.A(n_4292),
.B(n_4232),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_4292),
.B(n_4223),
.Y(n_4332)
);

INVxp67_ASAP7_75t_L g4333 ( 
.A(n_4305),
.Y(n_4333)
);

OA22x2_ASAP7_75t_L g4334 ( 
.A1(n_4247),
.A2(n_4240),
.B1(n_4223),
.B2(n_4243),
.Y(n_4334)
);

AND2x2_ASAP7_75t_L g4335 ( 
.A(n_4247),
.B(n_4240),
.Y(n_4335)
);

AND2x2_ASAP7_75t_L g4336 ( 
.A(n_4301),
.B(n_601),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4259),
.B(n_601),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4293),
.Y(n_4338)
);

INVx1_ASAP7_75t_SL g4339 ( 
.A(n_4266),
.Y(n_4339)
);

OAI22x1_ASAP7_75t_L g4340 ( 
.A1(n_4264),
.A2(n_602),
.B1(n_603),
.B2(n_604),
.Y(n_4340)
);

XNOR2x2_ASAP7_75t_L g4341 ( 
.A(n_4257),
.B(n_605),
.Y(n_4341)
);

NOR2xp33_ASAP7_75t_L g4342 ( 
.A(n_4260),
.B(n_605),
.Y(n_4342)
);

OA22x2_ASAP7_75t_L g4343 ( 
.A1(n_4254),
.A2(n_606),
.B1(n_608),
.B2(n_610),
.Y(n_4343)
);

XOR2x2_ASAP7_75t_L g4344 ( 
.A(n_4303),
.B(n_606),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4304),
.Y(n_4345)
);

HB1xp67_ASAP7_75t_L g4346 ( 
.A(n_4261),
.Y(n_4346)
);

INVx1_ASAP7_75t_SL g4347 ( 
.A(n_4249),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_4314),
.Y(n_4348)
);

INVx2_ASAP7_75t_L g4349 ( 
.A(n_4324),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4314),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4326),
.Y(n_4351)
);

AOI22xp5_ASAP7_75t_SL g4352 ( 
.A1(n_4317),
.A2(n_4330),
.B1(n_4323),
.B2(n_4334),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4338),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4320),
.Y(n_4354)
);

INVx1_ASAP7_75t_SL g4355 ( 
.A(n_4323),
.Y(n_4355)
);

INVxp67_ASAP7_75t_L g4356 ( 
.A(n_4342),
.Y(n_4356)
);

OA22x2_ASAP7_75t_L g4357 ( 
.A1(n_4328),
.A2(n_4300),
.B1(n_4277),
.B2(n_4294),
.Y(n_4357)
);

XOR2x2_ASAP7_75t_SL g4358 ( 
.A(n_4309),
.B(n_4298),
.Y(n_4358)
);

XOR2x2_ASAP7_75t_L g4359 ( 
.A(n_4316),
.B(n_4270),
.Y(n_4359)
);

HB1xp67_ASAP7_75t_L g4360 ( 
.A(n_4310),
.Y(n_4360)
);

OA22x2_ASAP7_75t_L g4361 ( 
.A1(n_4335),
.A2(n_4282),
.B1(n_4267),
.B2(n_4298),
.Y(n_4361)
);

INVx2_ASAP7_75t_L g4362 ( 
.A(n_4310),
.Y(n_4362)
);

OA22x2_ASAP7_75t_L g4363 ( 
.A1(n_4331),
.A2(n_4278),
.B1(n_4275),
.B2(n_4274),
.Y(n_4363)
);

OA22x2_ASAP7_75t_L g4364 ( 
.A1(n_4333),
.A2(n_4287),
.B1(n_4276),
.B2(n_4248),
.Y(n_4364)
);

AO22x1_ASAP7_75t_L g4365 ( 
.A1(n_4325),
.A2(n_4273),
.B1(n_4295),
.B2(n_4286),
.Y(n_4365)
);

OA22x2_ASAP7_75t_L g4366 ( 
.A1(n_4333),
.A2(n_4280),
.B1(n_4288),
.B2(n_4281),
.Y(n_4366)
);

AO22x1_ASAP7_75t_L g4367 ( 
.A1(n_4325),
.A2(n_4273),
.B1(n_4290),
.B2(n_4279),
.Y(n_4367)
);

CKINVDCx16_ASAP7_75t_R g4368 ( 
.A(n_4337),
.Y(n_4368)
);

INVx2_ASAP7_75t_SL g4369 ( 
.A(n_4339),
.Y(n_4369)
);

OAI22xp5_ASAP7_75t_L g4370 ( 
.A1(n_4334),
.A2(n_4253),
.B1(n_4283),
.B2(n_4272),
.Y(n_4370)
);

AO22x1_ASAP7_75t_L g4371 ( 
.A1(n_4332),
.A2(n_4306),
.B1(n_4302),
.B2(n_4291),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4313),
.Y(n_4372)
);

INVx2_ASAP7_75t_L g4373 ( 
.A(n_4311),
.Y(n_4373)
);

XNOR2xp5_ASAP7_75t_L g4374 ( 
.A(n_4308),
.B(n_608),
.Y(n_4374)
);

INVxp33_ASAP7_75t_SL g4375 ( 
.A(n_4342),
.Y(n_4375)
);

AOI22xp5_ASAP7_75t_L g4376 ( 
.A1(n_4315),
.A2(n_612),
.B1(n_613),
.B2(n_614),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_4339),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_4312),
.Y(n_4378)
);

XOR2x2_ASAP7_75t_L g4379 ( 
.A(n_4321),
.B(n_615),
.Y(n_4379)
);

XOR2x2_ASAP7_75t_L g4380 ( 
.A(n_4319),
.B(n_615),
.Y(n_4380)
);

AOI22xp5_ASAP7_75t_L g4381 ( 
.A1(n_4343),
.A2(n_617),
.B1(n_618),
.B2(n_619),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4318),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4322),
.Y(n_4383)
);

BUFx2_ASAP7_75t_L g4384 ( 
.A(n_4346),
.Y(n_4384)
);

OA22x2_ASAP7_75t_L g4385 ( 
.A1(n_4327),
.A2(n_617),
.B1(n_619),
.B2(n_620),
.Y(n_4385)
);

OAI22xp5_ASAP7_75t_L g4386 ( 
.A1(n_4347),
.A2(n_621),
.B1(n_622),
.B2(n_623),
.Y(n_4386)
);

XNOR2xp5_ASAP7_75t_L g4387 ( 
.A(n_4344),
.B(n_621),
.Y(n_4387)
);

XNOR2x2_ASAP7_75t_L g4388 ( 
.A(n_4341),
.B(n_623),
.Y(n_4388)
);

AOI22x1_ASAP7_75t_L g4389 ( 
.A1(n_4340),
.A2(n_4346),
.B1(n_4347),
.B2(n_4329),
.Y(n_4389)
);

INVx3_ASAP7_75t_L g4390 ( 
.A(n_4355),
.Y(n_4390)
);

INVxp67_ASAP7_75t_SL g4391 ( 
.A(n_4388),
.Y(n_4391)
);

OR2x2_ASAP7_75t_L g4392 ( 
.A(n_4362),
.B(n_4329),
.Y(n_4392)
);

AOI22xp5_ASAP7_75t_SL g4393 ( 
.A1(n_4366),
.A2(n_4343),
.B1(n_4336),
.B2(n_4345),
.Y(n_4393)
);

HB1xp67_ASAP7_75t_L g4394 ( 
.A(n_4360),
.Y(n_4394)
);

BUFx2_ASAP7_75t_L g4395 ( 
.A(n_4369),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4384),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4384),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4348),
.Y(n_4398)
);

CKINVDCx20_ASAP7_75t_R g4399 ( 
.A(n_4368),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4350),
.Y(n_4400)
);

INVx2_ASAP7_75t_L g4401 ( 
.A(n_4377),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4351),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4349),
.Y(n_4403)
);

HB1xp67_ASAP7_75t_L g4404 ( 
.A(n_4353),
.Y(n_4404)
);

OAI322xp33_ASAP7_75t_L g4405 ( 
.A1(n_4352),
.A2(n_4312),
.A3(n_625),
.B1(n_626),
.B2(n_627),
.C1(n_628),
.C2(n_629),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4354),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4383),
.Y(n_4407)
);

INVx8_ASAP7_75t_L g4408 ( 
.A(n_4385),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4372),
.Y(n_4409)
);

OAI322xp33_ASAP7_75t_L g4410 ( 
.A1(n_4357),
.A2(n_624),
.A3(n_625),
.B1(n_627),
.B2(n_628),
.C1(n_630),
.C2(n_631),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4382),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4378),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4373),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4364),
.Y(n_4414)
);

XOR2x2_ASAP7_75t_L g4415 ( 
.A(n_4358),
.B(n_624),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4361),
.Y(n_4416)
);

HB1xp67_ASAP7_75t_L g4417 ( 
.A(n_4356),
.Y(n_4417)
);

INVxp67_ASAP7_75t_L g4418 ( 
.A(n_4374),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4394),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4390),
.Y(n_4420)
);

NAND4xp75_ASAP7_75t_L g4421 ( 
.A(n_4416),
.B(n_4376),
.C(n_4381),
.D(n_4359),
.Y(n_4421)
);

AOI22xp5_ASAP7_75t_L g4422 ( 
.A1(n_4399),
.A2(n_4370),
.B1(n_4375),
.B2(n_4363),
.Y(n_4422)
);

AOI22xp5_ASAP7_75t_L g4423 ( 
.A1(n_4415),
.A2(n_4367),
.B1(n_4365),
.B2(n_4379),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4390),
.Y(n_4424)
);

OA22x2_ASAP7_75t_L g4425 ( 
.A1(n_4391),
.A2(n_4387),
.B1(n_4389),
.B2(n_4386),
.Y(n_4425)
);

OAI322xp33_ASAP7_75t_L g4426 ( 
.A1(n_4393),
.A2(n_4414),
.A3(n_4396),
.B1(n_4397),
.B2(n_4417),
.C1(n_4418),
.C2(n_4401),
.Y(n_4426)
);

AO22x2_ASAP7_75t_L g4427 ( 
.A1(n_4398),
.A2(n_4380),
.B1(n_4367),
.B2(n_4371),
.Y(n_4427)
);

OAI322xp33_ASAP7_75t_L g4428 ( 
.A1(n_4393),
.A2(n_4371),
.A3(n_632),
.B1(n_633),
.B2(n_634),
.C1(n_635),
.C2(n_636),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_4395),
.Y(n_4429)
);

OAI22xp33_ASAP7_75t_SL g4430 ( 
.A1(n_4400),
.A2(n_631),
.B1(n_632),
.B2(n_634),
.Y(n_4430)
);

INVx1_ASAP7_75t_SL g4431 ( 
.A(n_4392),
.Y(n_4431)
);

OAI22xp5_ASAP7_75t_L g4432 ( 
.A1(n_4408),
.A2(n_635),
.B1(n_636),
.B2(n_637),
.Y(n_4432)
);

OA22x2_ASAP7_75t_L g4433 ( 
.A1(n_4404),
.A2(n_637),
.B1(n_638),
.B2(n_639),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4402),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4403),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4406),
.Y(n_4436)
);

AOI22xp5_ASAP7_75t_SL g4437 ( 
.A1(n_4408),
.A2(n_638),
.B1(n_639),
.B2(n_640),
.Y(n_4437)
);

OAI22xp33_ASAP7_75t_L g4438 ( 
.A1(n_4408),
.A2(n_641),
.B1(n_642),
.B2(n_643),
.Y(n_4438)
);

AO22x2_ASAP7_75t_L g4439 ( 
.A1(n_4407),
.A2(n_644),
.B1(n_645),
.B2(n_647),
.Y(n_4439)
);

OA22x2_ASAP7_75t_L g4440 ( 
.A1(n_4410),
.A2(n_645),
.B1(n_647),
.B2(n_648),
.Y(n_4440)
);

OAI22xp33_ASAP7_75t_L g4441 ( 
.A1(n_4422),
.A2(n_4413),
.B1(n_4412),
.B2(n_4411),
.Y(n_4441)
);

NAND4xp25_ASAP7_75t_L g4442 ( 
.A(n_4423),
.B(n_4405),
.C(n_4409),
.D(n_652),
.Y(n_4442)
);

INVx1_ASAP7_75t_L g4443 ( 
.A(n_4420),
.Y(n_4443)
);

OAI22xp5_ASAP7_75t_L g4444 ( 
.A1(n_4427),
.A2(n_649),
.B1(n_651),
.B2(n_652),
.Y(n_4444)
);

OAI22x1_ASAP7_75t_L g4445 ( 
.A1(n_4429),
.A2(n_649),
.B1(n_654),
.B2(n_655),
.Y(n_4445)
);

AOI221xp5_ASAP7_75t_L g4446 ( 
.A1(n_4426),
.A2(n_655),
.B1(n_656),
.B2(n_659),
.C(n_660),
.Y(n_4446)
);

OAI22x1_ASAP7_75t_L g4447 ( 
.A1(n_4424),
.A2(n_659),
.B1(n_660),
.B2(n_661),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4419),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_4431),
.Y(n_4449)
);

OAI211xp5_ASAP7_75t_L g4450 ( 
.A1(n_4427),
.A2(n_661),
.B(n_663),
.C(n_664),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4439),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_4435),
.Y(n_4452)
);

OAI22xp5_ASAP7_75t_L g4453 ( 
.A1(n_4425),
.A2(n_663),
.B1(n_665),
.B2(n_666),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_4433),
.Y(n_4454)
);

AOI22xp5_ASAP7_75t_L g4455 ( 
.A1(n_4421),
.A2(n_667),
.B1(n_668),
.B2(n_670),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4437),
.Y(n_4456)
);

AOI22xp5_ASAP7_75t_L g4457 ( 
.A1(n_4432),
.A2(n_668),
.B1(n_670),
.B2(n_671),
.Y(n_4457)
);

INVxp67_ASAP7_75t_L g4458 ( 
.A(n_4440),
.Y(n_4458)
);

INVx2_ASAP7_75t_L g4459 ( 
.A(n_4449),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_L g4460 ( 
.A(n_4454),
.B(n_4438),
.Y(n_4460)
);

AOI22xp5_ASAP7_75t_L g4461 ( 
.A1(n_4444),
.A2(n_4434),
.B1(n_4436),
.B2(n_4428),
.Y(n_4461)
);

NOR2x1_ASAP7_75t_L g4462 ( 
.A(n_4450),
.B(n_4430),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4445),
.Y(n_4463)
);

AO22x2_ASAP7_75t_L g4464 ( 
.A1(n_4453),
.A2(n_671),
.B1(n_672),
.B2(n_674),
.Y(n_4464)
);

AOI22xp5_ASAP7_75t_L g4465 ( 
.A1(n_4455),
.A2(n_674),
.B1(n_675),
.B2(n_676),
.Y(n_4465)
);

NOR2x1_ASAP7_75t_L g4466 ( 
.A(n_4442),
.B(n_675),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4458),
.B(n_676),
.Y(n_4467)
);

AOI22xp5_ASAP7_75t_L g4468 ( 
.A1(n_4456),
.A2(n_677),
.B1(n_678),
.B2(n_679),
.Y(n_4468)
);

AOI22xp5_ASAP7_75t_L g4469 ( 
.A1(n_4441),
.A2(n_677),
.B1(n_678),
.B2(n_682),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4447),
.Y(n_4470)
);

AOI22xp5_ASAP7_75t_L g4471 ( 
.A1(n_4446),
.A2(n_682),
.B1(n_683),
.B2(n_684),
.Y(n_4471)
);

INVx1_ASAP7_75t_SL g4472 ( 
.A(n_4459),
.Y(n_4472)
);

BUFx4f_ASAP7_75t_SL g4473 ( 
.A(n_4463),
.Y(n_4473)
);

NOR2x1_ASAP7_75t_L g4474 ( 
.A(n_4467),
.B(n_4451),
.Y(n_4474)
);

NOR2x1_ASAP7_75t_L g4475 ( 
.A(n_4470),
.B(n_4448),
.Y(n_4475)
);

INVx2_ASAP7_75t_L g4476 ( 
.A(n_4464),
.Y(n_4476)
);

INVx2_ASAP7_75t_L g4477 ( 
.A(n_4464),
.Y(n_4477)
);

NOR3xp33_ASAP7_75t_L g4478 ( 
.A(n_4466),
.B(n_4443),
.C(n_4452),
.Y(n_4478)
);

NOR3xp33_ASAP7_75t_SL g4479 ( 
.A(n_4460),
.B(n_4457),
.C(n_684),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4468),
.Y(n_4480)
);

INVx2_ASAP7_75t_L g4481 ( 
.A(n_4462),
.Y(n_4481)
);

AOI22xp5_ASAP7_75t_L g4482 ( 
.A1(n_4461),
.A2(n_683),
.B1(n_685),
.B2(n_686),
.Y(n_4482)
);

NAND4xp25_ASAP7_75t_L g4483 ( 
.A(n_4482),
.B(n_4469),
.C(n_4471),
.D(n_4465),
.Y(n_4483)
);

AOI22xp5_ASAP7_75t_L g4484 ( 
.A1(n_4473),
.A2(n_685),
.B1(n_687),
.B2(n_688),
.Y(n_4484)
);

AOI22xp5_ASAP7_75t_L g4485 ( 
.A1(n_4481),
.A2(n_687),
.B1(n_689),
.B2(n_690),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4475),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4472),
.Y(n_4487)
);

INVx2_ASAP7_75t_L g4488 ( 
.A(n_4476),
.Y(n_4488)
);

AND4x1_ASAP7_75t_L g4489 ( 
.A(n_4479),
.B(n_689),
.C(n_692),
.D(n_693),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4487),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4484),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_4486),
.B(n_4477),
.Y(n_4492)
);

AOI22xp5_ASAP7_75t_L g4493 ( 
.A1(n_4490),
.A2(n_4480),
.B1(n_4483),
.B2(n_4478),
.Y(n_4493)
);

AOI22xp5_ASAP7_75t_L g4494 ( 
.A1(n_4491),
.A2(n_4474),
.B1(n_4488),
.B2(n_4485),
.Y(n_4494)
);

CKINVDCx20_ASAP7_75t_R g4495 ( 
.A(n_4493),
.Y(n_4495)
);

OAI22xp5_ASAP7_75t_L g4496 ( 
.A1(n_4495),
.A2(n_4494),
.B1(n_4492),
.B2(n_4489),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4496),
.Y(n_4497)
);

OAI22xp33_ASAP7_75t_SL g4498 ( 
.A1(n_4497),
.A2(n_692),
.B1(n_693),
.B2(n_694),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4498),
.Y(n_4499)
);

AOI221xp5_ASAP7_75t_L g4500 ( 
.A1(n_4499),
.A2(n_695),
.B1(n_696),
.B2(n_697),
.C(n_699),
.Y(n_4500)
);

AOI211xp5_ASAP7_75t_L g4501 ( 
.A1(n_4500),
.A2(n_695),
.B(n_696),
.C(n_699),
.Y(n_4501)
);


endmodule