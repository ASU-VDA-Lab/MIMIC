module fake_jpeg_14428_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_15),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_3),
.Y(n_17)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_18),
.B(n_9),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_4),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_8),
.B1(n_7),
.B2(n_11),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_23),
.B1(n_19),
.B2(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_18),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_23),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_15),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_32),
.B1(n_20),
.B2(n_24),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_34),
.Y(n_35)
);

OA21x2_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_30),
.B(n_5),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_5),
.Y(n_37)
);


endmodule