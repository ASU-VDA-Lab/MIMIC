module fake_jpeg_7556_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_23),
.B1(n_30),
.B2(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_45),
.Y(n_50)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_0),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_23),
.C(n_30),
.Y(n_59)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NAND2x1_ASAP7_75t_SL g76 ( 
.A(n_46),
.B(n_21),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_41),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_26),
.B1(n_20),
.B2(n_19),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_56),
.B1(n_58),
.B2(n_68),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_25),
.B1(n_34),
.B2(n_32),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_53),
.B(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_20),
.B1(n_35),
.B2(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_20),
.B1(n_19),
.B2(n_18),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_60),
.B(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_23),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_31),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_0),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_36),
.B1(n_34),
.B2(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_70),
.Y(n_98)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_75),
.B1(n_22),
.B2(n_11),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_41),
.B1(n_44),
.B2(n_21),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_87),
.B1(n_92),
.B2(n_109),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_44),
.B1(n_32),
.B2(n_25),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_83),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_81),
.B(n_49),
.Y(n_134)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_84),
.Y(n_139)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_94),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_44),
.B1(n_46),
.B2(n_22),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_48),
.B1(n_56),
.B2(n_71),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_55),
.B1(n_66),
.B2(n_54),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_90),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_46),
.B1(n_22),
.B2(n_17),
.Y(n_92)
);

AO22x2_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_67),
.B1(n_46),
.B2(n_62),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_93),
.A2(n_103),
.B(n_37),
.C(n_9),
.Y(n_144)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_99),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_11),
.Y(n_100)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_15),
.Y(n_119)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_104),
.Y(n_136)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_106),
.Y(n_140)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_60),
.A2(n_22),
.B1(n_37),
.B2(n_11),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_10),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx2_ASAP7_75t_R g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_121),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_74),
.C(n_59),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_143),
.C(n_145),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_119),
.A2(n_122),
.B1(n_126),
.B2(n_109),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_67),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_53),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_112),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_55),
.B1(n_68),
.B2(n_70),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_37),
.B(n_4),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_134),
.B(n_87),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_101),
.Y(n_148)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_90),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_37),
.C(n_70),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_144),
.A2(n_93),
.B1(n_85),
.B2(n_114),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_37),
.C(n_49),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_146),
.A2(n_175),
.B1(n_134),
.B2(n_129),
.Y(n_208)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_153),
.B1(n_168),
.B2(n_144),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_149),
.B(n_154),
.Y(n_210)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_155),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_108),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_115),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_100),
.B(n_115),
.C(n_82),
.D(n_101),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_161),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_159),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_160),
.A2(n_164),
.B(n_165),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_78),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_80),
.C(n_83),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_118),
.Y(n_200)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_167),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_121),
.A2(n_77),
.B(n_99),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_106),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_166),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_113),
.B1(n_49),
.B2(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_174),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_130),
.B(n_105),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_172),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_139),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_94),
.B1(n_86),
.B2(n_104),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_124),
.A2(n_1),
.B(n_4),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_124),
.B(n_133),
.Y(n_187)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_167),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_186),
.B(n_189),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_193),
.B(n_199),
.Y(n_233)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_191),
.B(n_197),
.Y(n_230)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_143),
.B(n_131),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_205),
.B1(n_162),
.B2(n_157),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_178),
.A2(n_131),
.B1(n_129),
.B2(n_119),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_157),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_164),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_201),
.B(n_207),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_137),
.C(n_130),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_208),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_160),
.A2(n_152),
.B(n_176),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_116),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_211),
.C(n_198),
.Y(n_220)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_209),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_153),
.A2(n_116),
.B1(n_146),
.B2(n_165),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_211),
.A2(n_174),
.B1(n_141),
.B2(n_123),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_177),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_220),
.C(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_217),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_195),
.Y(n_239)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_181),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_218),
.B(n_223),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_163),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_221),
.A2(n_225),
.B(n_232),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_150),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_189),
.A2(n_151),
.B1(n_170),
.B2(n_169),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_227),
.A2(n_230),
.B1(n_217),
.B2(n_215),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_229),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_210),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_161),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_179),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_208),
.B1(n_188),
.B2(n_185),
.Y(n_248)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_238),
.B1(n_138),
.B2(n_196),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_123),
.C(n_141),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_195),
.C(n_184),
.Y(n_241)
);

BUFx24_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_244),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_247),
.C(n_255),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_183),
.A3(n_186),
.B1(n_199),
.B2(n_197),
.C1(n_187),
.C2(n_193),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_224),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_213),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_183),
.C(n_205),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_250),
.B1(n_232),
.B2(n_238),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_193),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_257),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_185),
.B1(n_188),
.B2(n_182),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_182),
.C(n_192),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_202),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_202),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_260),
.C(n_4),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_173),
.C(n_90),
.Y(n_260)
);

AO21x1_ASAP7_75t_L g261 ( 
.A1(n_242),
.A2(n_225),
.B(n_234),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_261),
.A2(n_264),
.B(n_276),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_263),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_212),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_214),
.B(n_236),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_224),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_266),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_138),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_245),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_272),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_219),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_219),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_275),
.B(n_7),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_239),
.A2(n_232),
.B1(n_238),
.B2(n_90),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_240),
.C(n_241),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_257),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_280),
.B(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_284),
.C(n_291),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_251),
.B(n_247),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_285),
.A2(n_289),
.B(n_293),
.C(n_277),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g286 ( 
.A(n_264),
.B(n_240),
.CI(n_249),
.CON(n_286),
.SN(n_286)
);

AO22x1_ASAP7_75t_SL g301 ( 
.A1(n_286),
.A2(n_290),
.B1(n_287),
.B2(n_280),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_244),
.B(n_6),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_271),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_7),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_13),
.B(n_14),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_276),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_267),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_300),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_299),
.B(n_303),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_273),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_282),
.B1(n_289),
.B2(n_286),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_302),
.B(n_304),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_285),
.B(n_273),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_274),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_278),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_286),
.Y(n_306)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_306),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_281),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_14),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_284),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_299),
.C(n_295),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_298),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_317),
.C(n_309),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_313),
.A2(n_311),
.B1(n_301),
.B2(n_295),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_316),
.A2(n_320),
.B(n_314),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_5),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_312),
.B(n_310),
.Y(n_321)
);

OAI21x1_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_322),
.B(n_324),
.Y(n_326)
);

OAI321xp33_ASAP7_75t_L g325 ( 
.A1(n_323),
.A2(n_316),
.A3(n_6),
.B1(n_5),
.B2(n_12),
.C(n_8),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_5),
.B(n_8),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_12),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_326),
.Y(n_329)
);


endmodule