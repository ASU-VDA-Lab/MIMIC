module fake_jpeg_2749_n_607 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_607);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_607;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_57),
.B(n_69),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_58),
.B(n_62),
.Y(n_126)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_61),
.B(n_63),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_65),
.B(n_78),
.Y(n_172)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_66),
.Y(n_166)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_67),
.Y(n_128)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_23),
.B(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g155 ( 
.A(n_71),
.Y(n_155)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_20),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_100),
.B(n_40),
.Y(n_120)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_76),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_28),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_80),
.B(n_81),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_21),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_82),
.B(n_87),
.Y(n_175)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_33),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_33),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_25),
.B1(n_49),
.B2(n_47),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_38),
.B(n_0),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_96),
.B(n_98),
.Y(n_171)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_21),
.B(n_2),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_53),
.B(n_2),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_36),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_101),
.B(n_104),
.Y(n_173)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_21),
.B(n_3),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_41),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_110),
.Y(n_176)
);

INVx2_ASAP7_75t_R g108 ( 
.A(n_53),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_111),
.Y(n_130)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_41),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_48),
.B1(n_30),
.B2(n_51),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_118),
.A2(n_123),
.B1(n_124),
.B2(n_129),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_120),
.B(n_56),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_106),
.B1(n_75),
.B2(n_60),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_75),
.A2(n_40),
.B1(n_25),
.B2(n_51),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_141),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_78),
.A2(n_40),
.B1(n_25),
.B2(n_51),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_131),
.A2(n_157),
.B1(n_46),
.B2(n_53),
.Y(n_222)
);

INVx5_ASAP7_75t_SL g133 ( 
.A(n_56),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_133),
.B(n_26),
.Y(n_238)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_57),
.A2(n_22),
.B(n_52),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_81),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_63),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_49),
.B(n_47),
.C(n_37),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_149),
.A2(n_174),
.B(n_26),
.C(n_53),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_54),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_150),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_107),
.A2(n_49),
.B1(n_47),
.B2(n_37),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_152),
.A2(n_160),
.B1(n_162),
.B2(n_164),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_30),
.B1(n_37),
.B2(n_46),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_68),
.A2(n_83),
.B1(n_85),
.B2(n_109),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_79),
.A2(n_30),
.B1(n_50),
.B2(n_31),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_76),
.A2(n_54),
.B1(n_22),
.B2(n_52),
.Y(n_162)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_64),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_88),
.A2(n_54),
.B1(n_22),
.B2(n_52),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_61),
.A2(n_50),
.B1(n_42),
.B2(n_27),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_96),
.A2(n_89),
.B(n_97),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_178),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_172),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_181),
.B(n_183),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_182),
.A2(n_205),
.B1(n_222),
.B2(n_224),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_184),
.Y(n_243)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_185),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_186),
.B(n_195),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_55),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_187),
.B(n_191),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_188),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_175),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_189),
.B(n_199),
.Y(n_251)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_120),
.B(n_59),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_194),
.B(n_202),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_111),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_174),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_196),
.B(n_209),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_136),
.A2(n_94),
.B1(n_93),
.B2(n_92),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_197),
.A2(n_229),
.B(n_134),
.Y(n_272)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_145),
.Y(n_198)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_198),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_126),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_133),
.B(n_67),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_201),
.B(n_208),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_130),
.B(n_29),
.Y(n_202)
);

AO22x1_ASAP7_75t_SL g203 ( 
.A1(n_130),
.A2(n_103),
.B1(n_91),
.B2(n_86),
.Y(n_203)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_203),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_130),
.B(n_50),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_204),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_135),
.A2(n_84),
.B1(n_77),
.B2(n_74),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

INVx3_ASAP7_75t_SL g266 ( 
.A(n_206),
.Y(n_266)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_207),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_121),
.B(n_166),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_140),
.B(n_42),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_121),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_210),
.B(n_211),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_166),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_150),
.B(n_42),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_212),
.B(n_213),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_150),
.B(n_31),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_122),
.A2(n_27),
.B(n_29),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_214),
.B(n_227),
.C(n_236),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_143),
.B(n_72),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_215),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_157),
.A2(n_70),
.B1(n_46),
.B2(n_53),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_216),
.A2(n_241),
.B1(n_161),
.B2(n_137),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_144),
.Y(n_217)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_143),
.A2(n_46),
.B1(n_73),
.B2(n_26),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g250 ( 
.A1(n_219),
.A2(n_169),
.A3(n_167),
.B1(n_147),
.B2(n_155),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_128),
.B(n_71),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_220),
.B(n_231),
.Y(n_289)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_221),
.Y(n_286)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_119),
.Y(n_223)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_113),
.A2(n_139),
.B1(n_138),
.B2(n_137),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_142),
.Y(n_225)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_158),
.B(n_177),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_159),
.Y(n_228)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_230),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_112),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_128),
.B(n_3),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_232),
.B(n_233),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_147),
.B(n_3),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_132),
.Y(n_234)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_235),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_122),
.A2(n_53),
.B(n_26),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_112),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_237),
.B(n_4),
.Y(n_296)
);

NAND2x1_ASAP7_75t_SL g278 ( 
.A(n_238),
.B(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_158),
.Y(n_239)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_177),
.B(n_4),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_113),
.A2(n_53),
.B1(n_32),
.B2(n_6),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_125),
.Y(n_242)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_182),
.A2(n_125),
.B1(n_151),
.B2(n_155),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_244),
.A2(n_231),
.B1(n_192),
.B2(n_219),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_196),
.A2(n_114),
.B1(n_139),
.B2(n_163),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_246),
.A2(n_248),
.B1(n_262),
.B2(n_263),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_195),
.A2(n_200),
.B1(n_191),
.B2(n_179),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_250),
.B(n_272),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_193),
.A2(n_151),
.B1(n_132),
.B2(n_117),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_253),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_206),
.Y(n_255)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_190),
.Y(n_256)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_256),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_184),
.Y(n_257)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_257),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_222),
.A2(n_229),
.B1(n_226),
.B2(n_193),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_187),
.A2(n_114),
.B1(n_161),
.B2(n_138),
.Y(n_263)
);

NOR3xp33_ASAP7_75t_SL g267 ( 
.A(n_178),
.B(n_117),
.C(n_142),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_267),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_194),
.B(n_169),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_270),
.B(n_238),
.C(n_204),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_218),
.A2(n_197),
.B1(n_194),
.B2(n_209),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_273),
.A2(n_293),
.B1(n_294),
.B2(n_202),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_227),
.A2(n_134),
.B1(n_116),
.B2(n_32),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_275),
.A2(n_279),
.B1(n_211),
.B2(n_237),
.Y(n_322)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_207),
.Y(n_290)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_290),
.Y(n_333)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_242),
.Y(n_292)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_292),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_218),
.A2(n_116),
.B1(n_32),
.B2(n_6),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_203),
.A2(n_32),
.B1(n_5),
.B2(n_6),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_296),
.Y(n_324)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_185),
.Y(n_299)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_299),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_236),
.B(n_238),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_300),
.A2(n_302),
.B(n_316),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_247),
.B(n_268),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_301),
.B(n_305),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_272),
.A2(n_278),
.B(n_268),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_264),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_304),
.B(n_320),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_247),
.B(n_248),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_284),
.Y(n_307)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_307),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_251),
.B(n_186),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g377 ( 
.A(n_310),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_265),
.B(n_181),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_311),
.B(n_317),
.Y(n_360)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_252),
.Y(n_312)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_312),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_315),
.A2(n_192),
.B1(n_259),
.B2(n_258),
.Y(n_379)
);

A2O1A1O1Ixp25_ASAP7_75t_L g316 ( 
.A1(n_285),
.A2(n_212),
.B(n_213),
.C(n_204),
.D(n_202),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_254),
.B(n_199),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_269),
.A2(n_224),
.B1(n_205),
.B2(n_203),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_318),
.A2(n_339),
.B1(n_352),
.B2(n_249),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_319),
.B(n_351),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_289),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_240),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_321),
.B(n_326),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_322),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_254),
.B(n_230),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_325),
.B(n_335),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_285),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_260),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_329),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_295),
.B(n_240),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_328),
.B(n_332),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_287),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_284),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_227),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_277),
.C(n_290),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_271),
.B(n_214),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_278),
.Y(n_335)
);

INVx13_ASAP7_75t_L g337 ( 
.A(n_245),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_337),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_278),
.A2(n_219),
.B(n_239),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_338),
.A2(n_215),
.B(n_282),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_269),
.A2(n_262),
.B1(n_273),
.B2(n_246),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_287),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_340),
.B(n_344),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_271),
.B(n_203),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_341),
.B(n_347),
.Y(n_372)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_261),
.Y(n_342)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_342),
.Y(n_367)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_261),
.Y(n_343)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_343),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_299),
.Y(n_344)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_345),
.Y(n_371)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_274),
.Y(n_346)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_346),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_270),
.B(n_210),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_281),
.B(n_234),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_348),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_297),
.B(n_219),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_349),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_274),
.B(n_198),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_350),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_221),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_249),
.A2(n_241),
.B1(n_192),
.B2(n_184),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_313),
.A2(n_243),
.B1(n_252),
.B2(n_281),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_357),
.A2(n_392),
.B1(n_329),
.B2(n_344),
.Y(n_411)
);

OR2x6_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_294),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_359),
.B(n_217),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_362),
.A2(n_373),
.B1(n_385),
.B2(n_391),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_300),
.A2(n_250),
.B(n_243),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_365),
.A2(n_308),
.B(n_32),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_382),
.C(n_383),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_339),
.A2(n_263),
.B1(n_267),
.B2(n_277),
.Y(n_373)
);

AO22x1_ASAP7_75t_SL g374 ( 
.A1(n_306),
.A2(n_292),
.B1(n_282),
.B2(n_215),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_376),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_375),
.Y(n_400)
);

OAI32xp33_ASAP7_75t_L g376 ( 
.A1(n_305),
.A2(n_228),
.A3(n_235),
.B1(n_286),
.B2(n_283),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_379),
.A2(n_318),
.B1(n_352),
.B2(n_340),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_326),
.B(n_298),
.C(n_288),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_301),
.B(n_331),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_309),
.A2(n_298),
.B1(n_288),
.B2(n_286),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_302),
.A2(n_266),
.B(n_258),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_386),
.A2(n_338),
.B(n_349),
.Y(n_413)
);

OAI32xp33_ASAP7_75t_L g389 ( 
.A1(n_306),
.A2(n_283),
.A3(n_276),
.B1(n_259),
.B2(n_266),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_393),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_309),
.A2(n_276),
.B1(n_223),
.B2(n_180),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_313),
.A2(n_245),
.B1(n_255),
.B2(n_180),
.Y(n_392)
);

OAI32xp33_ASAP7_75t_L g393 ( 
.A1(n_306),
.A2(n_217),
.A3(n_225),
.B1(n_8),
.B2(n_10),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_394),
.Y(n_401)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_395),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_311),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_399),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_341),
.A2(n_217),
.B1(n_32),
.B2(n_8),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_397),
.A2(n_308),
.B1(n_337),
.B2(n_8),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_317),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_378),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_404),
.B(n_412),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_304),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g457 ( 
.A(n_405),
.Y(n_457)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_367),
.Y(n_407)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_407),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_327),
.Y(n_408)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_408),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_435),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_411),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_369),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_413),
.A2(n_425),
.B(n_432),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_356),
.B(n_320),
.Y(n_414)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_414),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_396),
.B(n_347),
.Y(n_415)
);

OAI21xp33_ASAP7_75t_SL g462 ( 
.A1(n_415),
.A2(n_426),
.B(n_431),
.Y(n_462)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_367),
.Y(n_417)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_417),
.Y(n_469)
);

NAND3xp33_ASAP7_75t_L g418 ( 
.A(n_360),
.B(n_328),
.C(n_324),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_418),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_381),
.B(n_319),
.C(n_351),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_421),
.C(n_427),
.Y(n_446)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_389),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_420),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_381),
.B(n_321),
.C(n_332),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_370),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_423),
.B(n_424),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_346),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_361),
.A2(n_316),
.B(n_303),
.Y(n_425)
);

AOI322xp5_ASAP7_75t_L g426 ( 
.A1(n_384),
.A2(n_315),
.A3(n_343),
.B1(n_342),
.B2(n_324),
.C1(n_334),
.C2(n_314),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_383),
.B(n_314),
.C(n_334),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_307),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_428),
.Y(n_444)
);

CKINVDCx14_ASAP7_75t_R g429 ( 
.A(n_353),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_429),
.A2(n_430),
.B1(n_433),
.B2(n_436),
.Y(n_448)
);

OAI21xp33_ASAP7_75t_L g430 ( 
.A1(n_368),
.A2(n_307),
.B(n_330),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_361),
.A2(n_336),
.B(n_323),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_371),
.A2(n_336),
.B1(n_323),
.B2(n_312),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_363),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_434),
.Y(n_468)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_370),
.Y(n_435)
);

NOR2x1_ASAP7_75t_R g437 ( 
.A(n_368),
.B(n_337),
.Y(n_437)
);

OAI21xp33_ASAP7_75t_SL g473 ( 
.A1(n_437),
.A2(n_359),
.B(n_376),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_438),
.A2(n_375),
.B(n_386),
.Y(n_460)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_380),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_439),
.A2(n_359),
.B1(n_390),
.B2(n_397),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_420),
.A2(n_365),
.B1(n_371),
.B2(n_372),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_441),
.A2(n_445),
.B1(n_463),
.B2(n_472),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_387),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_443),
.B(n_449),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_416),
.A2(n_398),
.B1(n_354),
.B2(n_384),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_402),
.B(n_387),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_419),
.B(n_382),
.C(n_366),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_451),
.C(n_454),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_398),
.C(n_364),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_421),
.B(n_355),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_404),
.A2(n_422),
.B1(n_416),
.B2(n_362),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_459),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_460),
.A2(n_461),
.B(n_413),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_400),
.A2(n_354),
.B(n_393),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_409),
.A2(n_379),
.B1(n_359),
.B2(n_374),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_425),
.B(n_374),
.C(n_395),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_465),
.B(n_466),
.C(n_471),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_415),
.B(n_373),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_422),
.A2(n_359),
.B1(n_391),
.B2(n_358),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_470),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_400),
.B(n_394),
.C(n_380),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_409),
.A2(n_359),
.B1(n_358),
.B2(n_385),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_473),
.B(n_403),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_437),
.B(n_369),
.C(n_363),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_474),
.B(n_431),
.C(n_438),
.Y(n_495)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_475),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_447),
.B(n_424),
.Y(n_476)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_476),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_412),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_479),
.B(n_485),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_457),
.B(n_428),
.Y(n_482)
);

CKINVDCx14_ASAP7_75t_R g508 ( 
.A(n_482),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_454),
.B(n_451),
.Y(n_483)
);

MAJx2_ASAP7_75t_L g514 ( 
.A(n_483),
.B(n_492),
.C(n_465),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_458),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_458),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_486),
.B(n_489),
.Y(n_521)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_453),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_487),
.B(n_488),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_432),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_469),
.Y(n_489)
);

CKINVDCx14_ASAP7_75t_R g513 ( 
.A(n_490),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_460),
.A2(n_431),
.B(n_406),
.Y(n_491)
);

NAND4xp25_ASAP7_75t_L g507 ( 
.A(n_491),
.B(n_500),
.C(n_461),
.D(n_479),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_443),
.B(n_449),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_444),
.B(n_435),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_493),
.B(n_497),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_474),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_456),
.B(n_439),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_496),
.A2(n_498),
.B1(n_499),
.B2(n_506),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_468),
.B(n_407),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_445),
.A2(n_406),
.B1(n_410),
.B2(n_417),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_452),
.A2(n_423),
.B1(n_403),
.B2(n_401),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_452),
.B(n_469),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_501),
.B(n_504),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_467),
.A2(n_401),
.B1(n_436),
.B2(n_390),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_502),
.A2(n_448),
.B1(n_472),
.B2(n_463),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_453),
.B(n_5),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_503),
.B(n_18),
.Y(n_522)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_455),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_442),
.B(n_7),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_507),
.A2(n_499),
.B(n_493),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_478),
.B(n_450),
.C(n_446),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_509),
.B(n_511),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_510),
.A2(n_520),
.B1(n_500),
.B2(n_476),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_478),
.B(n_446),
.C(n_471),
.Y(n_511)
);

XNOR2x1_ASAP7_75t_L g533 ( 
.A(n_514),
.B(n_516),
.Y(n_533)
);

AOI32xp33_ASAP7_75t_L g517 ( 
.A1(n_505),
.A2(n_440),
.A3(n_462),
.B1(n_442),
.B2(n_441),
.Y(n_517)
);

OAI211xp5_ASAP7_75t_L g552 ( 
.A1(n_517),
.A2(n_523),
.B(n_15),
.C(n_17),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_492),
.B(n_494),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_518),
.B(n_532),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_481),
.B(n_452),
.C(n_466),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_519),
.B(n_531),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_480),
.A2(n_440),
.B1(n_467),
.B2(n_11),
.Y(n_520)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_522),
.Y(n_535)
);

A2O1A1O1Ixp25_ASAP7_75t_L g523 ( 
.A1(n_485),
.A2(n_7),
.B(n_10),
.C(n_12),
.D(n_13),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_477),
.A2(n_7),
.B1(n_10),
.B2(n_12),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_526),
.A2(n_17),
.B1(n_18),
.B2(n_513),
.Y(n_553)
);

INVx11_ASAP7_75t_L g528 ( 
.A(n_496),
.Y(n_528)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_528),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_497),
.Y(n_529)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_529),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_481),
.B(n_18),
.C(n_15),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_494),
.B(n_14),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_534),
.A2(n_542),
.B1(n_548),
.B2(n_510),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_511),
.B(n_483),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_537),
.B(n_532),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_509),
.B(n_495),
.C(n_484),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_538),
.B(n_539),
.Y(n_558)
);

A2O1A1Ixp33_ASAP7_75t_SL g539 ( 
.A1(n_515),
.A2(n_484),
.B(n_491),
.C(n_502),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_519),
.B(n_490),
.C(n_501),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_540),
.B(n_547),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_524),
.A2(n_477),
.B1(n_486),
.B2(n_498),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_525),
.Y(n_543)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_543),
.Y(n_555)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_525),
.Y(n_546)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_546),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_506),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_516),
.B(n_489),
.C(n_504),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_549),
.B(n_551),
.C(n_512),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_518),
.B(n_15),
.C(n_16),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_552),
.B(n_523),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_553),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_545),
.B(n_531),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_554),
.B(n_566),
.Y(n_579)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_556),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_535),
.B(n_549),
.Y(n_557)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_557),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_SL g559 ( 
.A(n_533),
.B(n_514),
.Y(n_559)
);

MAJx2_ASAP7_75t_L g578 ( 
.A(n_559),
.B(n_570),
.C(n_533),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_563),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_562),
.A2(n_520),
.B1(n_521),
.B2(n_527),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_540),
.B(n_508),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_565),
.A2(n_567),
.B(n_568),
.Y(n_572)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_536),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_550),
.B(n_529),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_548),
.A2(n_515),
.B(n_512),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_538),
.B(n_521),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_541),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_571),
.B(n_527),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_561),
.B(n_542),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_573),
.Y(n_587)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_575),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_558),
.A2(n_507),
.B(n_539),
.Y(n_577)
);

MAJx2_ASAP7_75t_L g588 ( 
.A(n_577),
.B(n_578),
.C(n_560),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_580),
.B(n_581),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_570),
.B(n_537),
.C(n_563),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_569),
.B(n_544),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_582),
.B(n_564),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_555),
.A2(n_539),
.B1(n_526),
.B2(n_528),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_584),
.B(n_585),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_559),
.B(n_544),
.C(n_539),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_588),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_583),
.B(n_556),
.C(n_551),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_591),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_581),
.B(n_564),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g598 ( 
.A(n_592),
.B(n_594),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_574),
.B(n_576),
.C(n_572),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_590),
.B(n_574),
.C(n_579),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_595),
.A2(n_587),
.B(n_591),
.Y(n_601)
);

AOI321xp33_ASAP7_75t_L g596 ( 
.A1(n_586),
.A2(n_577),
.A3(n_578),
.B1(n_588),
.B2(n_582),
.C(n_593),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_596),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_601),
.B(n_602),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_598),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_600),
.A2(n_597),
.B(n_599),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_603),
.B(n_587),
.C(n_584),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_605),
.B(n_604),
.C(n_573),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_606),
.B(n_585),
.Y(n_607)
);


endmodule