module fake_jpeg_13595_n_614 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_614);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_614;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_63),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_27),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_65),
.B(n_84),
.Y(n_134)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_32),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_67),
.B(n_95),
.Y(n_206)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_75),
.Y(n_131)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_71),
.Y(n_190)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_79),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_80),
.Y(n_171)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_17),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_85),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_26),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_86),
.B(n_101),
.Y(n_164)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_20),
.B(n_17),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_93),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_20),
.B(n_16),
.Y(n_93)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_94),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_23),
.B(n_16),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

BUFx10_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_97),
.Y(n_183)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_100),
.Y(n_200)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_103),
.Y(n_203)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_23),
.B(n_16),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_114),
.Y(n_147)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_21),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_25),
.B(n_15),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_115),
.Y(n_174)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_34),
.Y(n_112)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_19),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_25),
.B(n_14),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_116),
.B(n_117),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_42),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_118),
.B(n_120),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_29),
.B(n_0),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_119),
.B(n_49),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_55),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_122),
.Y(n_184)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_21),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_21),
.B(n_2),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_129),
.B(n_163),
.C(n_12),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_135),
.B(n_139),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_97),
.A2(n_57),
.B1(n_21),
.B2(n_43),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_137),
.A2(n_161),
.B(n_182),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_59),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_L g143 ( 
.A1(n_69),
.A2(n_57),
.B1(n_43),
.B2(n_40),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_143),
.A2(n_159),
.B1(n_210),
.B2(n_152),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_66),
.B(n_59),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_145),
.B(n_29),
.Y(n_221)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_150),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_81),
.B(n_46),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_151),
.B(n_180),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_62),
.A2(n_43),
.B1(n_40),
.B2(n_30),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_105),
.A2(n_21),
.B1(n_40),
.B2(n_30),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_30),
.C(n_52),
.Y(n_163)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_64),
.Y(n_172)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_172),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_79),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_176),
.B(n_177),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_79),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_87),
.B(n_52),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_181),
.B(n_193),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_110),
.A2(n_58),
.B1(n_49),
.B2(n_48),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_48),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_187),
.B(n_198),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_124),
.A2(n_58),
.B1(n_46),
.B2(n_36),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_188),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_94),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_72),
.B(n_36),
.Y(n_198)
);

INVx6_ASAP7_75t_SL g199 ( 
.A(n_85),
.Y(n_199)
);

CKINVDCx11_ASAP7_75t_R g222 ( 
.A(n_199),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_113),
.B(n_33),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_201),
.B(n_208),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_102),
.B(n_35),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_204),
.B(n_12),
.Y(n_262)
);

INVx6_ASAP7_75t_SL g205 ( 
.A(n_74),
.Y(n_205)
);

BUFx12f_ASAP7_75t_SL g237 ( 
.A(n_205),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_78),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_207),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_80),
.B(n_33),
.Y(n_208)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_88),
.Y(n_209)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_211),
.B(n_212),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_127),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_213),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_164),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_214),
.B(n_230),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_159),
.A2(n_126),
.B1(n_111),
.B2(n_108),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_L g308 ( 
.A1(n_216),
.A2(n_239),
.B1(n_278),
.B2(n_179),
.Y(n_308)
);

AO22x1_ASAP7_75t_SL g218 ( 
.A1(n_142),
.A2(n_91),
.B1(n_89),
.B2(n_35),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_218),
.B(n_220),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_147),
.B(n_140),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_221),
.B(n_263),
.Y(n_284)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_223),
.Y(n_302)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_128),
.Y(n_224)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_131),
.B(n_1),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_225),
.B(n_233),
.Y(n_312)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_132),
.Y(n_226)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_226),
.Y(n_318)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_227),
.Y(n_309)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_149),
.Y(n_228)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

BUFx8_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

BUFx24_ASAP7_75t_L g293 ( 
.A(n_229),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_197),
.Y(n_230)
);

INVx13_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

INVx13_ASAP7_75t_L g305 ( 
.A(n_231),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_1),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_145),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_236),
.A2(n_248),
.B1(n_160),
.B2(n_162),
.Y(n_327)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_153),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_238),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_143),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_239)
);

INVx11_ASAP7_75t_L g240 ( 
.A(n_133),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_241),
.Y(n_310)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_243),
.Y(n_311)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_144),
.Y(n_244)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_244),
.Y(n_320)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_157),
.Y(n_245)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_245),
.Y(n_288)
);

BUFx8_ASAP7_75t_L g247 ( 
.A(n_173),
.Y(n_247)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_247),
.Y(n_340)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_200),
.Y(n_250)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_183),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_251),
.Y(n_319)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_148),
.Y(n_252)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_183),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_254),
.A2(n_281),
.B1(n_282),
.B2(n_130),
.Y(n_287)
);

CKINVDCx6p67_ASAP7_75t_R g255 ( 
.A(n_173),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_255),
.Y(n_314)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_127),
.Y(n_256)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_256),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_136),
.Y(n_257)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_257),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_139),
.A2(n_9),
.B(n_11),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_258),
.B(n_259),
.Y(n_313)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_148),
.Y(n_260)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_155),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_261),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_267),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_174),
.B(n_14),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_134),
.B(n_14),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_264),
.B(n_266),
.Y(n_324)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_175),
.Y(n_265)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_265),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_156),
.B(n_190),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_175),
.B(n_139),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_175),
.B(n_188),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_273),
.Y(n_303)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_166),
.Y(n_269)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_269),
.Y(n_315)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_194),
.Y(n_271)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_271),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_L g272 ( 
.A1(n_161),
.A2(n_137),
.B1(n_182),
.B2(n_202),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_272),
.A2(n_210),
.B1(n_186),
.B2(n_152),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_135),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_155),
.Y(n_274)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_274),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_191),
.B(n_168),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_279),
.Y(n_304)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_277),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_191),
.B(n_170),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_169),
.Y(n_280)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_280),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_138),
.A2(n_158),
.B1(n_146),
.B2(n_165),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_138),
.A2(n_209),
.B1(n_172),
.B2(n_130),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_150),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_166),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_287),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_251),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_295),
.B(n_316),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_297),
.A2(n_327),
.B1(n_232),
.B2(n_234),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_185),
.B1(n_186),
.B2(n_136),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_301),
.A2(n_307),
.B1(n_337),
.B2(n_256),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_246),
.B(n_185),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_325),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_218),
.A2(n_179),
.B1(n_178),
.B2(n_160),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_308),
.A2(n_280),
.B1(n_213),
.B2(n_257),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_251),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_317),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_251),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_321),
.B(n_222),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_242),
.B(n_235),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_220),
.B(n_141),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_335),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_217),
.B(n_141),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_217),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_272),
.A2(n_162),
.B1(n_171),
.B2(n_178),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_334),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_259),
.B(n_154),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_217),
.A2(n_154),
.B1(n_171),
.B2(n_218),
.Y(n_337)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_341),
.Y(n_385)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_291),
.Y(n_343)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_344),
.Y(n_402)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_345),
.Y(n_399)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_300),
.Y(n_347)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_347),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_348),
.Y(n_401)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_322),
.Y(n_349)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_349),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_350),
.A2(n_364),
.B1(n_378),
.B2(n_382),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_351),
.Y(n_410)
);

INVx13_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_352),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_325),
.B(n_219),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_353),
.B(n_356),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_244),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_366),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_324),
.B(n_215),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_326),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_365),
.Y(n_393)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_313),
.A2(n_276),
.B1(n_258),
.B2(n_243),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_359),
.A2(n_380),
.B(n_384),
.Y(n_397)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_360),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_361),
.B(n_362),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_293),
.Y(n_362)
);

INVx13_ASAP7_75t_L g363 ( 
.A(n_293),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_363),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_286),
.B(n_237),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_296),
.B(n_271),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_284),
.B(n_237),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_367),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_308),
.A2(n_276),
.B1(n_253),
.B2(n_277),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_369),
.B(n_371),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_223),
.C(n_227),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_332),
.C(n_329),
.Y(n_390)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_328),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_328),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_373),
.Y(n_395)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_336),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_339),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_375),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_376),
.A2(n_292),
.B1(n_332),
.B2(n_319),
.Y(n_387)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_336),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_379),
.Y(n_388)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_311),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_288),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_312),
.B(n_255),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_288),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_383),
.A2(n_340),
.B(n_294),
.Y(n_392)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_289),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_387),
.A2(n_405),
.B(n_369),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_390),
.B(n_398),
.C(n_412),
.Y(n_437)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_392),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_350),
.A2(n_292),
.B1(n_306),
.B2(n_313),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_396),
.A2(n_407),
.B1(n_411),
.B2(n_384),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_346),
.B(n_313),
.C(n_303),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_359),
.A2(n_337),
.B(n_297),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_368),
.A2(n_304),
.B(n_327),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_406),
.A2(n_352),
.B(n_363),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_381),
.A2(n_289),
.B1(n_290),
.B2(n_311),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_381),
.A2(n_346),
.B1(n_354),
.B2(n_342),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_370),
.B(n_298),
.C(n_318),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_342),
.B(n_299),
.C(n_315),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_420),
.C(n_329),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_351),
.B(n_290),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_416),
.B(n_419),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_351),
.B(n_339),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_355),
.B(n_315),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_357),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_422),
.B(n_423),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_383),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_395),
.Y(n_424)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_424),
.Y(n_464)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_395),
.Y(n_425)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_425),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_374),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_426),
.B(n_432),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_438),
.Y(n_456)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_428),
.Y(n_485)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_385),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_431),
.Y(n_461)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_386),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_393),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_374),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_433),
.B(n_443),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_388),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_434),
.B(n_436),
.Y(n_471)
);

CKINVDCx10_ASAP7_75t_R g435 ( 
.A(n_394),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_435),
.Y(n_473)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_386),
.Y(n_436)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_400),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_439),
.A2(n_396),
.B1(n_408),
.B2(n_420),
.Y(n_466)
);

AND2x6_ASAP7_75t_L g440 ( 
.A(n_397),
.B(n_368),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_440),
.A2(n_445),
.B(n_447),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_404),
.A2(n_364),
.B1(n_382),
.B2(n_379),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_442),
.A2(n_451),
.B1(n_454),
.B2(n_428),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_338),
.Y(n_443)
);

INVx13_ASAP7_75t_L g444 ( 
.A(n_394),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_444),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_411),
.A2(n_362),
.B(n_338),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_389),
.B(n_341),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_446),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_389),
.B(n_417),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_449),
.Y(n_468)
);

AO22x1_ASAP7_75t_SL g449 ( 
.A1(n_405),
.A2(n_347),
.B1(n_358),
.B2(n_343),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_377),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_450),
.B(n_455),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_391),
.A2(n_373),
.B1(n_372),
.B2(n_371),
.Y(n_451)
);

MAJx2_ASAP7_75t_L g475 ( 
.A(n_452),
.B(n_416),
.C(n_419),
.Y(n_475)
);

INVx13_ASAP7_75t_L g453 ( 
.A(n_404),
.Y(n_453)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_453),
.Y(n_467)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_400),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_454),
.B(n_408),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g455 ( 
.A(n_397),
.B(n_398),
.Y(n_455)
);

AO22x1_ASAP7_75t_L g458 ( 
.A1(n_449),
.A2(n_410),
.B1(n_391),
.B2(n_406),
.Y(n_458)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_458),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_390),
.C(n_410),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_459),
.B(n_480),
.C(n_486),
.Y(n_492)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_462),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_450),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_463),
.B(n_470),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_437),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_465),
.B(n_476),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_466),
.A2(n_481),
.B1(n_451),
.B2(n_445),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_447),
.A2(n_388),
.B(n_392),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_469),
.Y(n_494)
);

NOR3xp33_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_401),
.C(n_387),
.Y(n_470)
);

MAJx2_ASAP7_75t_L g514 ( 
.A(n_475),
.B(n_320),
.C(n_274),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_441),
.B(n_401),
.Y(n_476)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_479),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_425),
.C(n_424),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_439),
.A2(n_409),
.B1(n_399),
.B2(n_414),
.Y(n_481)
);

OA21x2_ASAP7_75t_L g483 ( 
.A1(n_449),
.A2(n_407),
.B(n_399),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_483),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_446),
.B(n_414),
.C(n_403),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_448),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_502),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_471),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_489),
.B(n_495),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_483),
.A2(n_429),
.B1(n_434),
.B2(n_427),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_490),
.A2(n_493),
.B1(n_499),
.B2(n_503),
.Y(n_524)
);

CKINVDCx14_ASAP7_75t_R g491 ( 
.A(n_472),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_491),
.B(n_500),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_483),
.A2(n_429),
.B1(n_432),
.B2(n_440),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_460),
.B(n_435),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_459),
.B(n_476),
.C(n_475),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_504),
.C(n_462),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_456),
.A2(n_430),
.B1(n_436),
.B2(n_438),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_474),
.B(n_431),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_501),
.A2(n_478),
.B1(n_457),
.B2(n_469),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_344),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_456),
.A2(n_402),
.B1(n_453),
.B2(n_403),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_402),
.C(n_360),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_462),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_506),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_456),
.A2(n_453),
.B1(n_345),
.B2(n_378),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_509),
.A2(n_511),
.B1(n_467),
.B2(n_473),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_466),
.B(n_349),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_510),
.B(n_485),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_464),
.A2(n_333),
.B1(n_330),
.B2(n_323),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_477),
.A2(n_330),
.B1(n_323),
.B2(n_333),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_512),
.B(n_481),
.Y(n_515)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_471),
.Y(n_513)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_513),
.Y(n_522)
);

XNOR2x1_ASAP7_75t_SL g530 ( 
.A(n_514),
.B(n_458),
.Y(n_530)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_515),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_516),
.B(n_530),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_484),
.C(n_464),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_519),
.B(n_523),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_494),
.A2(n_468),
.B(n_484),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_492),
.B(n_508),
.C(n_487),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_525),
.B(n_531),
.C(n_514),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_526),
.A2(n_497),
.B1(n_498),
.B2(n_493),
.Y(n_545)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_499),
.Y(n_527)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_527),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_505),
.B(n_461),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_528),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_488),
.A2(n_478),
.B1(n_461),
.B2(n_467),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_529),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_508),
.B(n_485),
.C(n_473),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_532),
.B(n_533),
.Y(n_548)
);

XOR2x1_ASAP7_75t_L g533 ( 
.A(n_490),
.B(n_458),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_534),
.A2(n_294),
.B1(n_249),
.B2(n_232),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_494),
.A2(n_482),
.B(n_444),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_535),
.B(n_536),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_502),
.B(n_482),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_503),
.Y(n_537)
);

AOI31xp33_ASAP7_75t_L g544 ( 
.A1(n_537),
.A2(n_538),
.A3(n_497),
.B(n_507),
.Y(n_544)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_511),
.Y(n_538)
);

BUFx12_ASAP7_75t_L g539 ( 
.A(n_535),
.Y(n_539)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_539),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_SL g540 ( 
.A(n_519),
.B(n_496),
.C(n_504),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_540),
.B(n_520),
.Y(n_558)
);

BUFx12_ASAP7_75t_L g541 ( 
.A(n_531),
.Y(n_541)
);

CKINVDCx14_ASAP7_75t_R g573 ( 
.A(n_541),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_543),
.B(n_556),
.Y(n_559)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_544),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_545),
.A2(n_522),
.B1(n_534),
.B2(n_521),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_517),
.A2(n_509),
.B(n_510),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_546),
.B(n_549),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_516),
.B(n_309),
.C(n_302),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_554),
.B(n_557),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_525),
.B(n_520),
.C(n_536),
.Y(n_556)
);

NOR3xp33_ASAP7_75t_SL g557 ( 
.A(n_522),
.B(n_255),
.C(n_305),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_558),
.B(n_541),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_542),
.B(n_521),
.Y(n_563)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_563),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_556),
.B(n_532),
.C(n_524),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_564),
.B(n_566),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_555),
.A2(n_518),
.B(n_528),
.Y(n_565)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_565),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_543),
.B(n_549),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_550),
.B(n_551),
.C(n_548),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_567),
.B(n_569),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_550),
.B(n_524),
.C(n_527),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_553),
.A2(n_526),
.B(n_523),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_570),
.B(n_557),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_548),
.B(n_533),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_571),
.B(n_572),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_564),
.B(n_551),
.C(n_547),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_574),
.B(n_581),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_561),
.A2(n_552),
.B1(n_545),
.B2(n_538),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_576),
.B(n_579),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_559),
.B(n_541),
.Y(n_580)
);

NAND3xp33_ASAP7_75t_L g587 ( 
.A(n_580),
.B(n_584),
.C(n_568),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_573),
.A2(n_515),
.B1(n_530),
.B2(n_539),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_583),
.Y(n_591)
);

NOR2x1_ASAP7_75t_L g584 ( 
.A(n_560),
.B(n_539),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_569),
.B(n_554),
.C(n_309),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_585),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_587),
.B(n_592),
.Y(n_601)
);

XOR2x2_ASAP7_75t_L g592 ( 
.A(n_582),
.B(n_567),
.Y(n_592)
);

AOI32xp33_ASAP7_75t_L g593 ( 
.A1(n_575),
.A2(n_563),
.A3(n_570),
.B1(n_560),
.B2(n_562),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_593),
.A2(n_585),
.B1(n_574),
.B2(n_584),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_578),
.A2(n_571),
.B1(n_562),
.B2(n_572),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_594),
.B(n_596),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_577),
.B(n_228),
.C(n_302),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_595),
.B(n_586),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g596 ( 
.A(n_581),
.B(n_305),
.C(n_255),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_597),
.B(n_598),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_590),
.B(n_586),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_599),
.B(n_600),
.Y(n_604)
);

AOI322xp5_ASAP7_75t_L g600 ( 
.A1(n_588),
.A2(n_576),
.A3(n_583),
.B1(n_240),
.B2(n_249),
.C1(n_283),
.C2(n_231),
.Y(n_600)
);

AOI322xp5_ASAP7_75t_L g603 ( 
.A1(n_588),
.A2(n_310),
.A3(n_320),
.B1(n_234),
.B2(n_241),
.C1(n_270),
.C2(n_265),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_603),
.B(n_270),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_605),
.A2(n_606),
.B(n_601),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_602),
.B(n_589),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_608),
.B(n_609),
.C(n_591),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_607),
.A2(n_604),
.B(n_602),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_610),
.A2(n_269),
.B1(n_310),
.B2(n_247),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_611),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_612),
.B(n_247),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_613),
.B(n_229),
.C(n_293),
.Y(n_614)
);


endmodule