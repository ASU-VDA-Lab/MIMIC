module fake_jpeg_26724_n_324 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_36),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_17),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_48),
.Y(n_112)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_52),
.B(n_53),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_18),
.Y(n_53)
);

AO22x1_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_20),
.B1(n_31),
.B2(n_24),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_24),
.B(n_31),
.C(n_32),
.Y(n_89)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_74),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_23),
.B1(n_20),
.B2(n_29),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_70),
.B1(n_76),
.B2(n_31),
.Y(n_106)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_75),
.B(n_33),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_23),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_68),
.Y(n_110)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_26),
.B1(n_22),
.B2(n_36),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_34),
.B1(n_18),
.B2(n_33),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_39),
.B(n_34),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_26),
.B1(n_22),
.B2(n_29),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_40),
.B(n_35),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_26),
.B1(n_24),
.B2(n_33),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_47),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_77),
.A2(n_81),
.B(n_89),
.Y(n_123)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_79),
.B(n_84),
.Y(n_139)
);

AND2x4_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_43),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_48),
.A2(n_32),
.B1(n_35),
.B2(n_34),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_83),
.A2(n_86),
.B1(n_97),
.B2(n_102),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_88),
.Y(n_147)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_90),
.B(n_91),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_53),
.C(n_71),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_96),
.C(n_49),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_94),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_47),
.C(n_44),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_19),
.B1(n_25),
.B2(n_27),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_72),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_56),
.B1(n_64),
.B2(n_54),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_57),
.B1(n_65),
.B2(n_44),
.Y(n_119)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_28),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_101),
.B(n_17),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_35),
.B1(n_28),
.B2(n_30),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_107),
.Y(n_124)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_66),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_105),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_19),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_74),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_55),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_69),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_17),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_51),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_67),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_30),
.B1(n_67),
.B2(n_51),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_49),
.B(n_61),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_117),
.A2(n_128),
.B(n_115),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_121),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_99),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_120),
.A2(n_125),
.B1(n_126),
.B2(n_95),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_30),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_122),
.B(n_92),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_65),
.B1(n_19),
.B2(n_25),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_77),
.A2(n_27),
.B1(n_19),
.B2(n_25),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_69),
.B1(n_27),
.B2(n_25),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_103),
.B1(n_107),
.B2(n_109),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_10),
.B1(n_12),
.B2(n_11),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_69),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_143),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_81),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_85),
.A2(n_0),
.B(n_1),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_89),
.B(n_91),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_8),
.B1(n_9),
.B2(n_16),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_27),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_0),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_99),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_168),
.B1(n_134),
.B2(n_126),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_77),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_155),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_152),
.A2(n_140),
.B(n_119),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_79),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_156),
.B(n_166),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_157),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_84),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_160),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_101),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_161),
.B(n_121),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_86),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_174),
.Y(n_201)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_81),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_164),
.A2(n_167),
.B(n_172),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_165),
.A2(n_136),
.B1(n_143),
.B2(n_120),
.Y(n_199)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_96),
.B1(n_99),
.B2(n_116),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_112),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_170),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_88),
.Y(n_170)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_177),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_78),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_175),
.A2(n_178),
.B(n_180),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_104),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_123),
.A2(n_114),
.B(n_78),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_181),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_87),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_87),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_180),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_191),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

NOR2x1p5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_133),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_197),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_154),
.B1(n_151),
.B2(n_153),
.Y(n_216)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_176),
.B(n_162),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_195),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_153),
.Y(n_225)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_120),
.B1(n_136),
.B2(n_119),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_198),
.A2(n_210),
.B1(n_165),
.B2(n_179),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_172),
.B1(n_154),
.B2(n_166),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_157),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_149),
.B(n_138),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_212),
.Y(n_222)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_146),
.C(n_147),
.Y(n_207)
);

NAND3xp33_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_7),
.C(n_15),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_119),
.B1(n_129),
.B2(n_95),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_213),
.A2(n_199),
.B1(n_185),
.B2(n_198),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_195),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_203),
.B(n_155),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_215),
.B(n_189),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g239 ( 
.A1(n_216),
.A2(n_217),
.B(n_227),
.C(n_193),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_158),
.B(n_171),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_149),
.C(n_202),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_221),
.C(n_229),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_164),
.C(n_161),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_225),
.B(n_230),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_191),
.A2(n_158),
.B(n_180),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_159),
.B1(n_175),
.B2(n_152),
.Y(n_228)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_186),
.C(n_209),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_160),
.Y(n_230)
);

A2O1A1O1Ixp25_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_128),
.B(n_146),
.C(n_67),
.D(n_88),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_212),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_132),
.C(n_82),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_184),
.C(n_195),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_80),
.B1(n_82),
.B2(n_132),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_238),
.B(n_12),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_258),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_242),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_223),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_241),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_220),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_201),
.B(n_229),
.C(n_224),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_201),
.B(n_189),
.C(n_226),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_188),
.Y(n_244)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

OAI22x1_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_236),
.B1(n_217),
.B2(n_227),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_246),
.A2(n_248),
.B1(n_253),
.B2(n_254),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_187),
.B1(n_205),
.B2(n_182),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_250),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_220),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_218),
.B1(n_182),
.B2(n_204),
.Y(n_277)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_255),
.A2(n_228),
.B1(n_210),
.B2(n_213),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_222),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_183),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_258),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_262),
.B(n_272),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_221),
.C(n_219),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_268),
.C(n_269),
.Y(n_279)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_225),
.C(n_222),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_230),
.C(n_211),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_273),
.C(n_274),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_192),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_192),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_218),
.C(n_233),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_243),
.C(n_239),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_80),
.C(n_1),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_259),
.B1(n_255),
.B2(n_253),
.Y(n_280)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_275),
.A2(n_246),
.B(n_259),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_289),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_283),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_263),
.A2(n_239),
.B(n_256),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_239),
.Y(n_286)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_261),
.A2(n_265),
.B(n_266),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_290),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_266),
.A2(n_0),
.B(n_1),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_2),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_286),
.A2(n_270),
.B1(n_264),
.B2(n_269),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_292),
.A2(n_293),
.B1(n_279),
.B2(n_6),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_285),
.A2(n_271),
.B1(n_268),
.B2(n_4),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_108),
.C(n_8),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_300),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_108),
.C(n_9),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_291),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_297),
.A2(n_287),
.B(n_288),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_296),
.A2(n_278),
.B(n_283),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_281),
.B(n_289),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_279),
.B1(n_282),
.B2(n_12),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_293),
.A3(n_294),
.B1(n_300),
.B2(n_295),
.C1(n_301),
.C2(n_292),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_309),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_294),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_315),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_6),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_312),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_6),
.A3(n_14),
.B1(n_15),
.B2(n_5),
.C1(n_2),
.C2(n_3),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_306),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_313),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_320),
.C(n_318),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_317),
.A2(n_311),
.B1(n_309),
.B2(n_302),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_312),
.B1(n_14),
.B2(n_5),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_4),
.Y(n_324)
);


endmodule