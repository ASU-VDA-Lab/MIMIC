module fake_jpeg_18141_n_57 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_57);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

AOI22x1_ASAP7_75t_L g38 ( 
.A1(n_20),
.A2(n_34),
.B1(n_32),
.B2(n_25),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_35),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_23),
.A2(n_17),
.B1(n_29),
.B2(n_27),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_21),
.B1(n_18),
.B2(n_24),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_45),
.B1(n_39),
.B2(n_42),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.C(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_47),
.B(n_38),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_43),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_53),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_41),
.B(n_37),
.Y(n_56)
);

AO21x1_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_36),
.B(n_40),
.Y(n_57)
);


endmodule