module fake_jpeg_8387_n_182 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_182);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_52),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_47),
.B(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_22),
.B1(n_30),
.B2(n_29),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_29),
.B1(n_37),
.B2(n_32),
.Y(n_68)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_29),
.B1(n_15),
.B2(n_26),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_26),
.B1(n_27),
.B2(n_19),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_16),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_39),
.Y(n_66)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_62),
.Y(n_82)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_35),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_39),
.B(n_40),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_70),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_73),
.B1(n_78),
.B2(n_83),
.Y(n_87)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_75),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_61),
.B(n_58),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_80),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_32),
.B1(n_33),
.B2(n_51),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_76),
.B1(n_50),
.B2(n_51),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_35),
.B(n_38),
.C(n_39),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_16),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_33),
.B1(n_25),
.B2(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_40),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_25),
.B1(n_28),
.B2(n_24),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_80),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_93),
.Y(n_103)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_59),
.A3(n_23),
.B1(n_17),
.B2(n_31),
.Y(n_85)
);

AO22x1_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_96),
.B1(n_49),
.B2(n_23),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_11),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_79),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_94),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_66),
.C(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_64),
.B(n_69),
.Y(n_94)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_54),
.Y(n_101)
);

NOR2xp67_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_65),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_43),
.B1(n_63),
.B2(n_52),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_70),
.B1(n_62),
.B2(n_49),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_119),
.B1(n_120),
.B2(n_92),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_65),
.B(n_75),
.C(n_73),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_109),
.B(n_114),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_108),
.C(n_87),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_98),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_77),
.C(n_82),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_43),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_0),
.B(n_1),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_115),
.B(n_116),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_118),
.B(n_90),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_117),
.B(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_86),
.Y(n_127)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_100),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_131),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_117),
.B(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_87),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_136),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_17),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_103),
.B(n_17),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_0),
.Y(n_146)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_141),
.Y(n_156)
);

INVxp33_ASAP7_75t_SL g140 ( 
.A(n_132),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

OAI321xp33_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_109),
.A3(n_105),
.B1(n_119),
.B2(n_24),
.C(n_21),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_146),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_122),
.B1(n_105),
.B2(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_139),
.A2(n_135),
.B1(n_128),
.B2(n_24),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_142),
.B1(n_141),
.B2(n_148),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_23),
.C(n_21),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_158),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_9),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_143),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_160),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_7),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_6),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_149),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_159),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_2),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_160),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_171),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_163),
.A2(n_157),
.B1(n_154),
.B2(n_156),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_5),
.B1(n_162),
.B2(n_168),
.Y(n_177)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_158),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_167),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_173),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_155),
.C(n_4),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_173),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_178),
.A2(n_179),
.B(n_174),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_175),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g182 ( 
.A(n_181),
.Y(n_182)
);


endmodule