module fake_jpeg_31395_n_64 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_64);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_64;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx3_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_8),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_16),
.A2(n_18),
.B1(n_2),
.B2(n_4),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_1),
.Y(n_30)
);

NOR3xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_21),
.C(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_26),
.B1(n_5),
.B2(n_6),
.Y(n_39)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_23),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_41),
.B1(n_27),
.B2(n_35),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_24),
.B1(n_22),
.B2(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_7),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_22),
.Y(n_49)
);

OA21x2_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_41),
.B(n_38),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_39),
.B(n_10),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

OAI322xp33_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_9),
.A3(n_13),
.B1(n_15),
.B2(n_19),
.C1(n_46),
.C2(n_50),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_50),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_54),
.C(n_55),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_62),
.B(n_58),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_54),
.C(n_53),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_60),
.B(n_9),
.Y(n_64)
);


endmodule