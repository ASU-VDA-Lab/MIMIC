module fake_jpeg_6686_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_37),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_0),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_43),
.B(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_36),
.B1(n_38),
.B2(n_33),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_21),
.B1(n_23),
.B2(n_18),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_52),
.B1(n_26),
.B2(n_28),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_20),
.B1(n_22),
.B2(n_19),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_53),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_17),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_29),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_20),
.B1(n_24),
.B2(n_27),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_71),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_82),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_58),
.B(n_51),
.C(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_79),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_54),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_56),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_36),
.B1(n_32),
.B2(n_33),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_85),
.B1(n_61),
.B2(n_46),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_38),
.B1(n_27),
.B2(n_28),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_31),
.B1(n_56),
.B2(n_57),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_31),
.B1(n_27),
.B2(n_29),
.Y(n_101)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_79),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_40),
.B1(n_35),
.B2(n_34),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_40),
.B1(n_31),
.B2(n_28),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_49),
.B1(n_40),
.B2(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_103),
.Y(n_118)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_45),
.Y(n_91)
);

NOR2x1_ASAP7_75t_SL g121 ( 
.A(n_91),
.B(n_85),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_92),
.A2(n_99),
.B1(n_89),
.B2(n_109),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_93),
.A2(n_66),
.B1(n_59),
.B2(n_3),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_46),
.B1(n_40),
.B2(n_49),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_101),
.B1(n_105),
.B2(n_70),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_98),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_24),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_71),
.B1(n_81),
.B2(n_78),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_34),
.C(n_57),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_104),
.C(n_68),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_110),
.B1(n_70),
.B2(n_82),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_34),
.C(n_57),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_59),
.B1(n_56),
.B2(n_24),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_66),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_79),
.B(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_73),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_112),
.B(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_116),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_123),
.B1(n_131),
.B2(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_85),
.B1(n_67),
.B2(n_75),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_125),
.B1(n_127),
.B2(n_93),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_85),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_121),
.A2(n_134),
.B(n_97),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_91),
.B(n_80),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_135),
.Y(n_145)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_103),
.C(n_109),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_82),
.B1(n_83),
.B2(n_75),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_68),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_106),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_130),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_59),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_1),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_150),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_107),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_143),
.B(n_117),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_107),
.B(n_88),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_159),
.B(n_117),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_96),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_153),
.C(n_157),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_111),
.B1(n_101),
.B2(n_105),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_148),
.A2(n_131),
.B1(n_122),
.B2(n_112),
.Y(n_169)
);

BUFx12_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_152),
.Y(n_161)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_111),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_123),
.B(n_106),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_134),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_135),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_4),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_116),
.A2(n_109),
.B1(n_97),
.B2(n_3),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_120),
.B1(n_124),
.B2(n_128),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_164),
.B(n_168),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_139),
.B1(n_145),
.B2(n_152),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_133),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_173),
.Y(n_183)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_171),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_159),
.A2(n_129),
.B(n_119),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_177),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_129),
.B(n_114),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_128),
.B1(n_134),
.B2(n_119),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_179),
.B1(n_181),
.B2(n_140),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_178),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_97),
.B1(n_2),
.B2(n_4),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_1),
.C(n_2),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_156),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_179)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_136),
.B1(n_139),
.B2(n_151),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_182),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_187),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_161),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_195),
.B1(n_200),
.B2(n_201),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_196),
.B(n_199),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_157),
.B1(n_155),
.B2(n_138),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_145),
.Y(n_197)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_176),
.A2(n_136),
.B1(n_143),
.B2(n_154),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_140),
.B1(n_182),
.B2(n_169),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_165),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_205),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_170),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_170),
.C(n_173),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_215),
.C(n_217),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_184),
.A2(n_164),
.B1(n_167),
.B2(n_168),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_211),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_184),
.A2(n_174),
.B1(n_160),
.B2(n_179),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_214),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_190),
.A2(n_143),
.B1(n_181),
.B2(n_175),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_178),
.C(n_150),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_149),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_150),
.C(n_149),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_215),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_150),
.B1(n_6),
.B2(n_5),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_194),
.B1(n_191),
.B2(n_197),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_209),
.B(n_185),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_200),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_208),
.B(n_188),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_217),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_187),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_207),
.A2(n_199),
.B1(n_210),
.B2(n_189),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_233),
.B(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_230),
.A2(n_232),
.B(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_213),
.B(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_191),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_192),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_238),
.B(n_239),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_206),
.C(n_203),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_236),
.C(n_225),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_237),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_242),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_219),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_222),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_243),
.A2(n_211),
.B1(n_221),
.B2(n_187),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_235),
.B1(n_205),
.B2(n_240),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_223),
.B1(n_229),
.B2(n_212),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_247),
.A2(n_251),
.B1(n_7),
.B2(n_10),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_14),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_249),
.A2(n_6),
.B(n_7),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_253),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_244),
.A2(n_214),
.B1(n_225),
.B2(n_8),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_252),
.A2(n_236),
.B(n_245),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_256),
.B(n_257),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_259),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_254),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_247),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_260),
.B(n_252),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g263 ( 
.A(n_261),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_262),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_261),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_12),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_264),
.A2(n_10),
.B(n_11),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_265),
.C(n_263),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_12),
.B1(n_13),
.B2(n_271),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_13),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_13),
.Y(n_274)
);


endmodule