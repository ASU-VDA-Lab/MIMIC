module fake_jpeg_9504_n_276 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_31),
.B1(n_29),
.B2(n_21),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_50),
.B1(n_52),
.B2(n_55),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_31),
.B1(n_29),
.B2(n_21),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_51),
.B1(n_64),
.B2(n_32),
.Y(n_70)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_31),
.B1(n_24),
.B2(n_29),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_22),
.B1(n_30),
.B2(n_26),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_24),
.B1(n_17),
.B2(n_20),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_28),
.B1(n_33),
.B2(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_28),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_23),
.B(n_33),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_19),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_22),
.B1(n_30),
.B2(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_68),
.B(n_70),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_75),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_88),
.Y(n_102)
);

NOR2x1_ASAP7_75t_R g74 ( 
.A(n_48),
.B(n_34),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_5),
.C(n_16),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_25),
.B1(n_23),
.B2(n_55),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_82),
.B1(n_96),
.B2(n_100),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_78),
.Y(n_116)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_18),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_83),
.Y(n_117)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_80),
.Y(n_128)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_44),
.A2(n_46),
.B1(n_52),
.B2(n_53),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_87),
.Y(n_126)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_49),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_98),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_34),
.B1(n_9),
.B2(n_10),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_92),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_34),
.B1(n_9),
.B2(n_10),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_34),
.B1(n_10),
.B2(n_12),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_49),
.B(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_19),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_95),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_53),
.A2(n_19),
.B1(n_8),
.B2(n_12),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_45),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_45),
.A2(n_19),
.B(n_1),
.C(n_2),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_47),
.A2(n_19),
.B1(n_7),
.B2(n_8),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_47),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_5),
.B1(n_7),
.B2(n_16),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_88),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_112),
.C(n_96),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_6),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_106),
.Y(n_141)
);

AOI32xp33_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_6),
.A3(n_14),
.B1(n_13),
.B2(n_8),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_76),
.C(n_5),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_0),
.C(n_1),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_0),
.B(n_1),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_99),
.B(n_94),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_127),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_122),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_87),
.B1(n_100),
.B2(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_71),
.Y(n_132)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_80),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_134),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_80),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_157),
.B(n_102),
.Y(n_175)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_154),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_158),
.B(n_102),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_144),
.Y(n_165)
);

OAI21x1_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_110),
.B(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_73),
.B(n_97),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_145),
.A2(n_155),
.B(n_156),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_115),
.A2(n_70),
.B1(n_81),
.B2(n_72),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_105),
.B1(n_121),
.B2(n_119),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_112),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_83),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_150),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_98),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_65),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_85),
.Y(n_153)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_85),
.B(n_77),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_104),
.A2(n_0),
.B(n_3),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_3),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_72),
.B(n_67),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_146),
.B1(n_154),
.B2(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_171),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_105),
.B1(n_106),
.B2(n_125),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_168),
.A2(n_179),
.B1(n_134),
.B2(n_131),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_185),
.B1(n_131),
.B2(n_132),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_180),
.C(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_175),
.B(n_177),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_145),
.C(n_153),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_184),
.C(n_182),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_125),
.B(n_114),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_130),
.A2(n_121),
.B1(n_124),
.B2(n_67),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_77),
.C(n_158),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_135),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_144),
.C(n_136),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_141),
.A2(n_130),
.B1(n_143),
.B2(n_142),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_133),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_193),
.C(n_207),
.Y(n_216)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_202),
.B1(n_203),
.B2(n_164),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_191),
.B(n_200),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_150),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_192),
.B(n_196),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_135),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_152),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_173),
.B(n_156),
.CI(n_157),
.CON(n_198),
.SN(n_198)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_199),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_157),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_170),
.B(n_157),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_SL g201 ( 
.A1(n_185),
.A2(n_151),
.A3(n_139),
.B1(n_147),
.B2(n_155),
.C1(n_138),
.C2(n_154),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_201),
.B(n_165),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_160),
.A2(n_139),
.B1(n_155),
.B2(n_151),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_146),
.C(n_154),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_206),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_175),
.B(n_177),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_194),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_212),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_164),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_184),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_215),
.C(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_218),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_162),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_217),
.A2(n_222),
.B1(n_197),
.B2(n_202),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_195),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_190),
.Y(n_220)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g221 ( 
.A(n_204),
.B(n_163),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_178),
.B(n_159),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_163),
.B1(n_171),
.B2(n_166),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_200),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_205),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_231),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_213),
.B(n_197),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_239),
.C(n_213),
.Y(n_240)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_209),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_210),
.B(n_219),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_188),
.B1(n_198),
.B2(n_186),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_214),
.B1(n_221),
.B2(n_223),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_165),
.C(n_198),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_241),
.C(n_244),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_215),
.C(n_216),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_211),
.C(n_221),
.Y(n_244)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_238),
.B(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_230),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_224),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_250),
.B(n_178),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_234),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_256),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_253),
.B(n_257),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_254),
.A2(n_244),
.B(n_240),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_233),
.B1(n_228),
.B2(n_209),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_254),
.B(n_247),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_258),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_252),
.A2(n_249),
.B1(n_236),
.B2(n_243),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_262),
.C(n_263),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_241),
.B(n_234),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_252),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_255),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_245),
.C(n_226),
.Y(n_271)
);

AOI31xp33_ASAP7_75t_L g270 ( 
.A1(n_267),
.A2(n_262),
.A3(n_253),
.B(n_245),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_270),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_268),
.B(n_269),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_274),
.A2(n_273),
.B(n_265),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_275),
.Y(n_276)
);


endmodule