module fake_jpeg_29498_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_25),
.B(n_39),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_0),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

HAxp5_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_69),
.CON(n_80),
.SN(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_1),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_19),
.C(n_42),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_55),
.B(n_57),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_59),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_60),
.B1(n_57),
.B2(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_73),
.B1(n_18),
.B2(n_40),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_49),
.B1(n_51),
.B2(n_54),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_51),
.B(n_56),
.C(n_53),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_47),
.B1(n_48),
.B2(n_44),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_2),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g81 ( 
.A(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_43),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_83),
.B(n_87),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_10),
.B(n_38),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_92),
.B1(n_72),
.B2(n_8),
.Y(n_100)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_91),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_103)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_4),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_5),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_27),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_6),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_99),
.Y(n_101)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_6),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_103),
.B1(n_111),
.B2(n_113),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_22),
.C(n_36),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_109),
.C(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_106),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_11),
.C(n_12),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_31),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_118),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_35),
.B1(n_100),
.B2(n_113),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_121),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_114),
.C(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_123),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_112),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_126),
.B(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_127),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_126),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_130),
.A2(n_131),
.B(n_119),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_136),
.Y(n_138)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_137),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_130),
.C(n_133),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_128),
.B1(n_122),
.B2(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);


endmodule