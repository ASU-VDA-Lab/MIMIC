module fake_jpeg_7749_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_155;
wire n_207;
wire n_31;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_28),
.B1(n_18),
.B2(n_30),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_40),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_48),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_21),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_24),
.B1(n_38),
.B2(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_55),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_57),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_16),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_24),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_33),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_65),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_64),
.B1(n_66),
.B2(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_32),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_36),
.A2(n_17),
.B1(n_29),
.B2(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_24),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_73),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_54),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_79),
.B(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_83),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_81),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_0),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_0),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_44),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_44),
.A2(n_41),
.B1(n_22),
.B2(n_20),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_88),
.B1(n_43),
.B2(n_66),
.Y(n_101)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_50),
.B1(n_49),
.B2(n_60),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_86),
.B(n_58),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_89),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_41),
.B1(n_22),
.B2(n_20),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_26),
.B(n_17),
.C(n_29),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_94),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_43),
.B1(n_53),
.B2(n_56),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_97),
.B1(n_83),
.B2(n_84),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_113),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_62),
.B1(n_51),
.B2(n_64),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_104),
.B(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_101),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_102),
.B(n_90),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_53),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_110),
.B1(n_87),
.B2(n_73),
.Y(n_134)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_108),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_78),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_71),
.B(n_34),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_68),
.C(n_69),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_50),
.B1(n_49),
.B2(n_60),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_74),
.B(n_63),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_55),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_68),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_117),
.Y(n_149)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_70),
.Y(n_120)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx2_ASAP7_75t_R g121 ( 
.A(n_102),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_82),
.B(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_128),
.B1(n_133),
.B2(n_138),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_86),
.B1(n_104),
.B2(n_111),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_77),
.Y(n_130)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_80),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_139),
.B1(n_112),
.B2(n_110),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_111),
.C(n_69),
.Y(n_142)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_100),
.B(n_80),
.Y(n_139)
);

OAI21x1_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_131),
.B(n_99),
.Y(n_154)
);

CKINVDCx12_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_145),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_146),
.C(n_159),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_129),
.B(n_135),
.Y(n_183)
);

CKINVDCx12_ASAP7_75t_R g145 ( 
.A(n_121),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_115),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_95),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_147),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_97),
.A3(n_95),
.B1(n_101),
.B2(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_157),
.B1(n_152),
.B2(n_159),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_144),
.Y(n_176)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_156),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_104),
.B1(n_111),
.B2(n_108),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_114),
.C(n_57),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_114),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_137),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_114),
.C(n_11),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_162),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_88),
.B1(n_52),
.B2(n_60),
.Y(n_163)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_123),
.B1(n_122),
.B2(n_117),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_168),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_175),
.C(n_177),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_137),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_176),
.B(n_179),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_118),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_144),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_160),
.B(n_126),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_140),
.B1(n_125),
.B2(n_126),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_134),
.B(n_129),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_157),
.B1(n_151),
.B2(n_143),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_148),
.A2(n_125),
.B1(n_116),
.B2(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_125),
.B1(n_132),
.B2(n_120),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_139),
.B1(n_129),
.B2(n_105),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_34),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_65),
.C(n_46),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_149),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_201),
.B(n_202),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_143),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_187),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_156),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_203),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_153),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_204),
.B(n_206),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_155),
.C(n_166),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_210),
.C(n_214),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_155),
.C(n_46),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_164),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_212),
.A2(n_213),
.B1(n_173),
.B2(n_178),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_94),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_107),
.C(n_34),
.Y(n_214)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_182),
.B1(n_184),
.B2(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_211),
.A2(n_182),
.B1(n_183),
.B2(n_169),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_220),
.B(n_226),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_175),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_222),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_177),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_191),
.B1(n_105),
.B2(n_107),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_227),
.B1(n_203),
.B2(n_194),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_170),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_87),
.B1(n_25),
.B2(n_27),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_37),
.C(n_34),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_230),
.C(n_231),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_37),
.C(n_23),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_23),
.C(n_73),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_211),
.A2(n_25),
.B1(n_27),
.B2(n_73),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_232),
.A2(n_192),
.B1(n_205),
.B2(n_27),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_22),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_239),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_217),
.A2(n_198),
.B1(n_206),
.B2(n_212),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_224),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_207),
.B1(n_218),
.B2(n_198),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_247),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_233),
.B(n_193),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_224),
.C(n_226),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_207),
.C(n_201),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_251),
.C(n_31),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_202),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_232),
.B(n_9),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_248),
.B(n_14),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_23),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_250),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_54),
.C(n_23),
.Y(n_251)
);

AO221x1_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_234),
.B1(n_233),
.B2(n_230),
.C(n_229),
.Y(n_252)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_265),
.Y(n_277)
);

AO21x1_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_260),
.B(n_262),
.Y(n_276)
);

AOI322xp5_ASAP7_75t_SL g255 ( 
.A1(n_237),
.A2(n_234),
.A3(n_9),
.B1(n_10),
.B2(n_14),
.C1(n_13),
.C2(n_8),
.Y(n_255)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_2),
.C(n_3),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_31),
.C(n_8),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_240),
.C(n_245),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_2),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_SL g262 ( 
.A1(n_249),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_236),
.B(n_13),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_263),
.B(n_264),
.Y(n_269)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_10),
.B(n_9),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_1),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_269),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_241),
.B1(n_238),
.B2(n_240),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_267),
.A3(n_276),
.B1(n_266),
.B2(n_277),
.C1(n_274),
.C2(n_262),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_270),
.B(n_272),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_243),
.B(n_251),
.Y(n_271)
);

NOR3xp33_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_273),
.C(n_262),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_23),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_3),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_244),
.C(n_31),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_244),
.C(n_268),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_285),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_280),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_255),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_281),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_4),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_286),
.C(n_4),
.Y(n_292)
);

INVx11_ASAP7_75t_L g285 ( 
.A(n_276),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_3),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_4),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_291),
.B(n_292),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_4),
.B(n_5),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_279),
.B(n_6),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_5),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_291),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_295),
.A2(n_297),
.B(n_287),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_283),
.B(n_286),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_298),
.A2(n_299),
.B1(n_288),
.B2(n_296),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_6),
.C(n_7),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_301),
.B(n_6),
.Y(n_302)
);


endmodule