module fake_aes_2677_n_1568 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_374, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_376, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_377, n_343, n_127, n_291, n_170, n_356, n_281, n_341, n_58, n_122, n_187, n_375, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1568);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_374;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_376;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_377;
input n_343;
input n_127;
input n_291;
input n_170;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_375;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1568;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1533;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_1563;
wire n_824;
wire n_793;
wire n_753;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_1557;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1432;
wire n_1315;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_688;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_606;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_386;
wire n_659;
wire n_432;
wire n_1329;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_401;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_1275;
wire n_955;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1389;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_600;
wire n_1531;
wire n_1548;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_210), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_175), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_231), .Y(n_380) );
INVxp67_ASAP7_75t_L g381 ( .A(n_57), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_160), .B(n_208), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_16), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_320), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_44), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_175), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_337), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_352), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_336), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_90), .Y(n_390) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_242), .B(n_34), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_372), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_274), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_123), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_269), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_324), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_123), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_311), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_303), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_17), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_260), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_136), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_275), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_246), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_226), .Y(n_405) );
INVxp33_ASAP7_75t_SL g406 ( .A(n_218), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_180), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_111), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_101), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_166), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_188), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_157), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_66), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_293), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_209), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_193), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_80), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_130), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_159), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_69), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_318), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_328), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_27), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_207), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_224), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_249), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_304), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_358), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_179), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_370), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_96), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_78), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_168), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_368), .Y(n_434) );
INVxp33_ASAP7_75t_SL g435 ( .A(n_5), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_202), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_200), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_333), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_143), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_84), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_189), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_79), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g443 ( .A(n_230), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_16), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_20), .Y(n_445) );
INVx4_ASAP7_75t_R g446 ( .A(n_302), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_38), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_184), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_10), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_119), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_355), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_340), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_237), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_288), .Y(n_454) );
INVxp67_ASAP7_75t_L g455 ( .A(n_96), .Y(n_455) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_92), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_213), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_362), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_28), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_74), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_332), .B(n_72), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_285), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_204), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_326), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_1), .Y(n_465) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_363), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_113), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_334), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_11), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_143), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_192), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_298), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_35), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_206), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_196), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_270), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_82), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_371), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_166), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_297), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_162), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_69), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_151), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_290), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_150), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_27), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_193), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_177), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_339), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_28), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_20), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_103), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_140), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_137), .Y(n_494) );
BUFx5_ASAP7_75t_L g495 ( .A(n_281), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_21), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_278), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_65), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_29), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_145), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_261), .Y(n_501) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_283), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_147), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_50), .Y(n_504) );
CKINVDCx14_ASAP7_75t_R g505 ( .A(n_118), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_159), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_313), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_235), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_105), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_51), .Y(n_510) );
INVx1_ASAP7_75t_SL g511 ( .A(n_146), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_7), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_219), .Y(n_513) );
INVx3_ASAP7_75t_L g514 ( .A(n_366), .Y(n_514) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_369), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_239), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_54), .Y(n_517) );
INVxp67_ASAP7_75t_SL g518 ( .A(n_68), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_296), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_300), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_268), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_364), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_264), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_250), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_365), .Y(n_525) );
NOR2xp67_ASAP7_75t_L g526 ( .A(n_199), .B(n_321), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_287), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_43), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_148), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_104), .Y(n_530) );
INVxp67_ASAP7_75t_SL g531 ( .A(n_15), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_198), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_203), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_178), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_280), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_106), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_350), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_116), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_1), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_117), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_146), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_314), .Y(n_542) );
BUFx3_ASAP7_75t_L g543 ( .A(n_54), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_9), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_227), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_73), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_168), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_323), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_291), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_158), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_216), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_9), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_221), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_252), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_26), .Y(n_555) );
INVxp33_ASAP7_75t_L g556 ( .A(n_187), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_282), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_108), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_154), .Y(n_559) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_129), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_46), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_40), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_197), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_346), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_91), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_105), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_121), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_93), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_243), .Y(n_569) );
INVxp67_ASAP7_75t_L g570 ( .A(n_110), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_465), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_514), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_556), .B(n_0), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_405), .B(n_0), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_480), .B(n_2), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_514), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_465), .B(n_2), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_505), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_514), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_465), .B(n_3), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_556), .B(n_4), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_400), .Y(n_582) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_436), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_505), .Y(n_584) );
BUFx8_ASAP7_75t_L g585 ( .A(n_382), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_495), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_495), .Y(n_587) );
AND2x6_ASAP7_75t_L g588 ( .A(n_382), .B(n_201), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_458), .B(n_6), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_495), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_495), .Y(n_591) );
CKINVDCx11_ASAP7_75t_R g592 ( .A(n_390), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_495), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_534), .A2(n_8), .B1(n_6), .B2(n_7), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_450), .Y(n_595) );
AND2x2_ASAP7_75t_SL g596 ( .A(n_382), .B(n_205), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_495), .Y(n_597) );
INVx4_ASAP7_75t_L g598 ( .A(n_462), .Y(n_598) );
OAI22xp5_ASAP7_75t_SL g599 ( .A1(n_390), .A2(n_11), .B1(n_8), .B2(n_10), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_436), .Y(n_600) );
BUFx3_ASAP7_75t_L g601 ( .A(n_462), .Y(n_601) );
CKINVDCx6p67_ASAP7_75t_R g602 ( .A(n_443), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_458), .B(n_12), .Y(n_603) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_436), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_436), .B(n_12), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_440), .B(n_13), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_491), .Y(n_607) );
INVx3_ASAP7_75t_L g608 ( .A(n_402), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_466), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_571), .B(n_415), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_602), .B(n_472), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_573), .B(n_479), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_573), .A2(n_504), .B1(n_386), .B2(n_408), .Y(n_613) );
BUFx4f_ASAP7_75t_L g614 ( .A(n_588), .Y(n_614) );
OR2x6_ASAP7_75t_L g615 ( .A(n_578), .B(n_418), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_573), .A2(n_410), .B1(n_411), .B2(n_407), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_581), .B(n_517), .Y(n_617) );
INVx3_ASAP7_75t_L g618 ( .A(n_589), .Y(n_618) );
NAND2xp33_ASAP7_75t_SL g619 ( .A(n_584), .B(n_497), .Y(n_619) );
OR2x6_ASAP7_75t_L g620 ( .A(n_578), .B(n_544), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_571), .B(n_484), .Y(n_621) );
INVx4_ASAP7_75t_SL g622 ( .A(n_588), .Y(n_622) );
AND2x2_ASAP7_75t_SL g623 ( .A(n_596), .B(n_533), .Y(n_623) );
OAI22xp33_ASAP7_75t_L g624 ( .A1(n_602), .A2(n_379), .B1(n_397), .B2(n_394), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_585), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_608), .B(n_392), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_585), .B(n_378), .Y(n_627) );
INVx4_ASAP7_75t_L g628 ( .A(n_588), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_586), .Y(n_629) );
INVx2_ASAP7_75t_SL g630 ( .A(n_585), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_583), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_583), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_586), .Y(n_633) );
INVx4_ASAP7_75t_L g634 ( .A(n_588), .Y(n_634) );
AND2x6_ASAP7_75t_L g635 ( .A(n_589), .B(n_380), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_581), .A2(n_423), .B1(n_429), .B2(n_417), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_585), .B(n_378), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_583), .Y(n_638) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_583), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_587), .Y(n_640) );
AND2x6_ASAP7_75t_L g641 ( .A(n_589), .B(n_384), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_585), .B(n_404), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_583), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_587), .Y(n_644) );
CKINVDCx14_ASAP7_75t_R g645 ( .A(n_602), .Y(n_645) );
AND2x6_ASAP7_75t_L g646 ( .A(n_589), .B(n_387), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_623), .A2(n_596), .B1(n_612), .B2(n_617), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_623), .A2(n_596), .B1(n_588), .B2(n_589), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_612), .B(n_581), .Y(n_649) );
BUFx3_ASAP7_75t_L g650 ( .A(n_625), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_617), .B(n_606), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_610), .B(n_606), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_618), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_623), .A2(n_588), .B1(n_606), .B2(n_603), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_618), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_626), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_610), .B(n_574), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_621), .B(n_574), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_621), .B(n_575), .Y(n_659) );
INVx5_ASAP7_75t_L g660 ( .A(n_635), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_635), .A2(n_588), .B1(n_435), .B2(n_608), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_635), .B(n_575), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_626), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_635), .B(n_601), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g665 ( .A(n_645), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_635), .B(n_601), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_618), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_619), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_611), .Y(n_669) );
OR2x6_ASAP7_75t_L g670 ( .A(n_615), .B(n_599), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_624), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_635), .B(n_641), .Y(n_672) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_625), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_618), .Y(n_674) );
INVx2_ASAP7_75t_SL g675 ( .A(n_641), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_613), .A2(n_457), .B1(n_557), .B2(n_497), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_627), .B(n_637), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_641), .A2(n_588), .B1(n_435), .B2(n_608), .Y(n_678) );
INVx8_ASAP7_75t_L g679 ( .A(n_641), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_642), .B(n_577), .Y(n_680) );
NAND2xp33_ASAP7_75t_SL g681 ( .A(n_630), .B(n_457), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_615), .Y(n_682) );
NAND2x1p5_ASAP7_75t_L g683 ( .A(n_630), .B(n_614), .Y(n_683) );
O2A1O1Ixp5_ASAP7_75t_L g684 ( .A1(n_614), .A2(n_598), .B(n_605), .C(n_580), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_629), .Y(n_685) );
AND2x4_ASAP7_75t_L g686 ( .A(n_630), .B(n_641), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_641), .B(n_598), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_641), .A2(n_588), .B1(n_557), .B2(n_599), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_628), .B(n_590), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_628), .B(n_590), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_646), .B(n_577), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_646), .B(n_580), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_646), .B(n_608), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_646), .A2(n_406), .B1(n_475), .B2(n_402), .Y(n_694) );
OAI21xp5_ASAP7_75t_L g695 ( .A1(n_629), .A2(n_591), .B(n_590), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_633), .Y(n_696) );
A2O1A1Ixp33_ASAP7_75t_SL g697 ( .A1(n_633), .A2(n_461), .B(n_593), .C(n_591), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_616), .B(n_394), .C(n_379), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_636), .B(n_414), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_615), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_640), .Y(n_701) );
O2A1O1Ixp5_ASAP7_75t_L g702 ( .A1(n_614), .A2(n_576), .B(n_579), .C(n_572), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g703 ( .A(n_615), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_640), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_644), .Y(n_705) );
AND2x6_ASAP7_75t_SL g706 ( .A(n_615), .B(n_592), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_634), .B(n_451), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_622), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_622), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_634), .B(n_451), .Y(n_710) );
OR2x6_ASAP7_75t_L g711 ( .A(n_620), .B(n_594), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_634), .B(n_463), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_620), .A2(n_412), .B1(n_416), .B2(n_397), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_622), .B(n_463), .Y(n_714) );
INVx2_ASAP7_75t_SL g715 ( .A(n_620), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_622), .B(n_464), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_620), .B(n_412), .Y(n_717) );
BUFx3_ASAP7_75t_L g718 ( .A(n_665), .Y(n_718) );
INVx2_ASAP7_75t_SL g719 ( .A(n_658), .Y(n_719) );
O2A1O1Ixp33_ASAP7_75t_L g720 ( .A1(n_649), .A2(n_620), .B(n_594), .C(n_455), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_656), .Y(n_721) );
OAI22xp5_ASAP7_75t_SL g722 ( .A1(n_700), .A2(n_409), .B1(n_433), .B2(n_413), .Y(n_722) );
INVx1_ASAP7_75t_SL g723 ( .A(n_663), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_685), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_648), .A2(n_413), .B1(n_433), .B2(n_409), .Y(n_725) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_650), .Y(n_726) );
INVx3_ASAP7_75t_L g727 ( .A(n_679), .Y(n_727) );
BUFx6f_ASAP7_75t_L g728 ( .A(n_650), .Y(n_728) );
BUFx2_ASAP7_75t_L g729 ( .A(n_681), .Y(n_729) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_679), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_690), .A2(n_597), .B(n_576), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_647), .A2(n_448), .B1(n_541), .B2(n_510), .Y(n_732) );
AND2x4_ASAP7_75t_L g733 ( .A(n_715), .B(n_456), .Y(n_733) );
BUFx2_ASAP7_75t_SL g734 ( .A(n_700), .Y(n_734) );
INVxp67_ASAP7_75t_L g735 ( .A(n_657), .Y(n_735) );
NOR2xp33_ASAP7_75t_SL g736 ( .A(n_679), .B(n_448), .Y(n_736) );
NOR2xp33_ASAP7_75t_SL g737 ( .A(n_679), .B(n_510), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_659), .B(n_652), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_669), .B(n_540), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_651), .B(n_540), .Y(n_740) );
O2A1O1Ixp33_ASAP7_75t_L g741 ( .A1(n_671), .A2(n_536), .B(n_562), .C(n_381), .Y(n_741) );
O2A1O1Ixp33_ASAP7_75t_L g742 ( .A1(n_699), .A2(n_570), .B(n_531), .C(n_518), .Y(n_742) );
O2A1O1Ixp33_ASAP7_75t_L g743 ( .A1(n_697), .A2(n_431), .B(n_441), .C(n_439), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_717), .B(n_541), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_698), .B(n_547), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_704), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_654), .A2(n_688), .B1(n_662), .B2(n_691), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_692), .A2(n_550), .B1(n_555), .B2(n_547), .Y(n_748) );
NOR2xp33_ASAP7_75t_SL g749 ( .A(n_660), .B(n_464), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_682), .A2(n_555), .B1(n_558), .B2(n_550), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_706), .Y(n_751) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_673), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_653), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_713), .A2(n_561), .B1(n_566), .B2(n_558), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_703), .B(n_561), .Y(n_755) );
AO32x1_ASAP7_75t_L g756 ( .A1(n_697), .A2(n_609), .A3(n_600), .B1(n_396), .B2(n_399), .Y(n_756) );
BUFx2_ASAP7_75t_L g757 ( .A(n_676), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_704), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_711), .B(n_566), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_670), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_711), .A2(n_567), .B1(n_385), .B2(n_420), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_661), .A2(n_567), .B1(n_525), .B2(n_527), .Y(n_762) );
NOR3xp33_ASAP7_75t_SL g763 ( .A(n_670), .B(n_432), .C(n_419), .Y(n_763) );
INVx2_ASAP7_75t_SL g764 ( .A(n_711), .Y(n_764) );
A2O1A1Ixp33_ASAP7_75t_L g765 ( .A1(n_680), .A2(n_543), .B(n_445), .C(n_449), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_705), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_653), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_680), .B(n_442), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_670), .B(n_383), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_677), .A2(n_469), .B1(n_477), .B2(n_471), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_705), .B(n_444), .Y(n_771) );
BUFx2_ASAP7_75t_L g772 ( .A(n_668), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_653), .Y(n_773) );
NOR3xp33_ASAP7_75t_SL g774 ( .A(n_677), .B(n_492), .C(n_487), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_694), .B(n_493), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_668), .B(n_511), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_667), .Y(n_777) );
INVx3_ASAP7_75t_L g778 ( .A(n_686), .Y(n_778) );
NAND2x1p5_ASAP7_75t_L g779 ( .A(n_660), .B(n_582), .Y(n_779) );
A2O1A1Ixp33_ASAP7_75t_L g780 ( .A1(n_696), .A2(n_459), .B(n_460), .C(n_447), .Y(n_780) );
A2O1A1Ixp33_ASAP7_75t_L g781 ( .A1(n_701), .A2(n_470), .B(n_473), .C(n_467), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_678), .B(n_512), .Y(n_782) );
A2O1A1Ixp33_ASAP7_75t_L g783 ( .A1(n_702), .A2(n_482), .B(n_483), .C(n_481), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_655), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_687), .A2(n_632), .B(n_631), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_660), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_655), .A2(n_638), .B(n_632), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_674), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_686), .B(n_496), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_674), .A2(n_643), .B(n_638), .Y(n_790) );
INVx1_ASAP7_75t_SL g791 ( .A(n_660), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_672), .A2(n_525), .B1(n_527), .B2(n_522), .Y(n_792) );
O2A1O1Ixp33_ASAP7_75t_L g793 ( .A1(n_693), .A2(n_486), .B(n_488), .C(n_485), .Y(n_793) );
BUFx6f_ASAP7_75t_L g794 ( .A(n_673), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_675), .A2(n_542), .B1(n_545), .B2(n_522), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_684), .Y(n_796) );
BUFx6f_ASAP7_75t_L g797 ( .A(n_673), .Y(n_797) );
NAND2xp5_ASAP7_75t_SL g798 ( .A(n_686), .B(n_542), .Y(n_798) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_664), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_707), .B(n_499), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_710), .B(n_500), .Y(n_801) );
AOI21x1_ASAP7_75t_L g802 ( .A1(n_666), .A2(n_643), .B(n_526), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_712), .A2(n_395), .B(n_388), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_683), .A2(n_553), .B1(n_554), .B2(n_545), .Y(n_804) );
NAND2xp5_ASAP7_75t_SL g805 ( .A(n_673), .B(n_553), .Y(n_805) );
BUFx3_ASAP7_75t_L g806 ( .A(n_708), .Y(n_806) );
A2O1A1Ixp33_ASAP7_75t_L g807 ( .A1(n_695), .A2(n_494), .B(n_498), .C(n_490), .Y(n_807) );
NOR3xp33_ASAP7_75t_L g808 ( .A(n_714), .B(n_509), .C(n_506), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_716), .B(n_503), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_709), .Y(n_810) );
INVx3_ASAP7_75t_L g811 ( .A(n_683), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_689), .A2(n_403), .B(n_401), .Y(n_812) );
OAI21xp33_ASAP7_75t_L g813 ( .A1(n_657), .A2(n_529), .B(n_528), .Y(n_813) );
O2A1O1Ixp33_ASAP7_75t_L g814 ( .A1(n_649), .A2(n_530), .B(n_538), .C(n_532), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_648), .A2(n_554), .B1(n_539), .B2(n_546), .Y(n_815) );
INVxp33_ASAP7_75t_SL g816 ( .A(n_676), .Y(n_816) );
O2A1O1Ixp33_ASAP7_75t_SL g817 ( .A1(n_697), .A2(n_425), .B(n_427), .C(n_424), .Y(n_817) );
INVx4_ASAP7_75t_L g818 ( .A(n_679), .Y(n_818) );
NAND2x1_ASAP7_75t_SL g819 ( .A(n_713), .B(n_391), .Y(n_819) );
O2A1O1Ixp33_ASAP7_75t_L g820 ( .A1(n_649), .A2(n_552), .B(n_565), .C(n_559), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_656), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_648), .A2(n_568), .B1(n_563), .B2(n_491), .Y(n_822) );
NOR2xp33_ASAP7_75t_R g823 ( .A(n_681), .B(n_389), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_647), .A2(n_428), .B1(n_434), .B2(n_430), .Y(n_824) );
OAI21xp5_ASAP7_75t_L g825 ( .A1(n_702), .A2(n_438), .B(n_437), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_656), .Y(n_826) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_665), .Y(n_827) );
AOI22xp33_ASAP7_75t_SL g828 ( .A1(n_816), .A2(n_563), .B1(n_560), .B2(n_595), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_757), .A2(n_560), .B1(n_454), .B2(n_474), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_719), .B(n_607), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_735), .B(n_607), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_723), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_738), .A2(n_489), .B(n_452), .Y(n_833) );
NAND4xp25_ASAP7_75t_SL g834 ( .A(n_720), .B(n_398), .C(n_426), .D(n_422), .Y(n_834) );
OAI21xp5_ASAP7_75t_L g835 ( .A1(n_825), .A2(n_508), .B(n_501), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_721), .B(n_560), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_744), .B(n_560), .Y(n_837) );
AO21x1_ASAP7_75t_L g838 ( .A1(n_743), .A2(n_523), .B(n_520), .Y(n_838) );
AO32x2_ASAP7_75t_L g839 ( .A1(n_822), .A2(n_604), .A3(n_609), .B1(n_600), .B2(n_446), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_759), .A2(n_535), .B1(n_537), .B2(n_524), .Y(n_840) );
INVx6_ASAP7_75t_SL g841 ( .A(n_733), .Y(n_841) );
A2O1A1Ixp33_ASAP7_75t_L g842 ( .A1(n_803), .A2(n_569), .B(n_564), .C(n_421), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_732), .A2(n_548), .B1(n_549), .B2(n_393), .Y(n_843) );
INVx2_ASAP7_75t_SL g844 ( .A(n_718), .Y(n_844) );
A2O1A1Ixp33_ASAP7_75t_L g845 ( .A1(n_793), .A2(n_549), .B(n_551), .C(n_548), .Y(n_845) );
OAI21xp5_ASAP7_75t_L g846 ( .A1(n_783), .A2(n_551), .B(n_600), .Y(n_846) );
OR2x2_ASAP7_75t_L g847 ( .A(n_725), .B(n_13), .Y(n_847) );
OAI21xp5_ASAP7_75t_L g848 ( .A1(n_825), .A2(n_609), .B(n_453), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_821), .B(n_468), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_736), .A2(n_476), .B1(n_507), .B2(n_478), .Y(n_850) );
NOR2xp33_ASAP7_75t_SL g851 ( .A(n_736), .B(n_513), .Y(n_851) );
A2O1A1Ixp33_ASAP7_75t_L g852 ( .A1(n_826), .A2(n_502), .B(n_515), .C(n_466), .Y(n_852) );
A2O1A1Ixp33_ASAP7_75t_L g853 ( .A1(n_814), .A2(n_502), .B(n_515), .C(n_466), .Y(n_853) );
AO31x2_ASAP7_75t_L g854 ( .A1(n_796), .A2(n_604), .A3(n_515), .B(n_516), .Y(n_854) );
BUFx2_ASAP7_75t_L g855 ( .A(n_823), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_724), .Y(n_856) );
AOI21xp33_ASAP7_75t_L g857 ( .A1(n_739), .A2(n_519), .B(n_515), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_764), .B(n_14), .Y(n_858) );
AOI21xp5_ASAP7_75t_L g859 ( .A1(n_785), .A2(n_639), .B(n_516), .Y(n_859) );
O2A1O1Ixp33_ASAP7_75t_L g860 ( .A1(n_765), .A2(n_17), .B(n_14), .C(n_15), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_771), .B(n_18), .Y(n_861) );
AOI221xp5_ASAP7_75t_L g862 ( .A1(n_741), .A2(n_521), .B1(n_516), .B2(n_502), .C(n_604), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_737), .A2(n_521), .B1(n_516), .B2(n_604), .Y(n_863) );
BUFx2_ASAP7_75t_SL g864 ( .A(n_818), .Y(n_864) );
AO21x2_ASAP7_75t_L g865 ( .A1(n_817), .A2(n_604), .B(n_639), .Y(n_865) );
BUFx4f_ASAP7_75t_SL g866 ( .A(n_772), .Y(n_866) );
OR2x2_ASAP7_75t_L g867 ( .A(n_722), .B(n_18), .Y(n_867) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_760), .B(n_19), .Y(n_868) );
A2O1A1Ixp33_ASAP7_75t_L g869 ( .A1(n_820), .A2(n_604), .B(n_639), .C(n_22), .Y(n_869) );
NAND3x1_ASAP7_75t_L g870 ( .A(n_769), .B(n_19), .C(n_21), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_824), .A2(n_25), .B1(n_23), .B2(n_24), .Y(n_871) );
A2O1A1Ixp33_ASAP7_75t_L g872 ( .A1(n_809), .A2(n_29), .B(n_23), .C(n_26), .Y(n_872) );
A2O1A1Ixp33_ASAP7_75t_L g873 ( .A1(n_800), .A2(n_32), .B(n_30), .C(n_31), .Y(n_873) );
O2A1O1Ixp33_ASAP7_75t_SL g874 ( .A1(n_807), .A2(n_212), .B(n_214), .C(n_211), .Y(n_874) );
INVx3_ASAP7_75t_L g875 ( .A(n_730), .Y(n_875) );
AOI21xp5_ASAP7_75t_L g876 ( .A1(n_746), .A2(n_217), .B(n_215), .Y(n_876) );
NAND2xp5_ASAP7_75t_SL g877 ( .A(n_737), .B(n_32), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_758), .Y(n_878) );
OAI21x1_ASAP7_75t_L g879 ( .A1(n_787), .A2(n_222), .B(n_220), .Y(n_879) );
BUFx2_ASAP7_75t_L g880 ( .A(n_776), .Y(n_880) );
OAI21x1_ASAP7_75t_L g881 ( .A1(n_790), .A2(n_225), .B(n_223), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_766), .Y(n_882) );
A2O1A1Ixp33_ASAP7_75t_L g883 ( .A1(n_801), .A2(n_35), .B(n_33), .C(n_34), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_777), .Y(n_884) );
INVx1_ASAP7_75t_SL g885 ( .A(n_734), .Y(n_885) );
INVx6_ASAP7_75t_L g886 ( .A(n_733), .Y(n_886) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_827), .Y(n_887) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_750), .Y(n_888) );
OR2x2_ASAP7_75t_L g889 ( .A(n_754), .B(n_36), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_782), .B(n_36), .Y(n_890) );
AOI21xp5_ASAP7_75t_L g891 ( .A1(n_731), .A2(n_229), .B(n_228), .Y(n_891) );
AO32x2_ASAP7_75t_L g892 ( .A1(n_815), .A2(n_39), .A3(n_37), .B1(n_38), .B2(n_40), .Y(n_892) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_804), .Y(n_893) );
O2A1O1Ixp33_ASAP7_75t_SL g894 ( .A1(n_780), .A2(n_233), .B(n_234), .C(n_232), .Y(n_894) );
BUFx3_ASAP7_75t_L g895 ( .A(n_751), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_740), .Y(n_896) );
INVx1_ASAP7_75t_SL g897 ( .A(n_779), .Y(n_897) );
A2O1A1Ixp33_ASAP7_75t_L g898 ( .A1(n_742), .A2(n_41), .B(n_37), .C(n_39), .Y(n_898) );
AO31x2_ASAP7_75t_L g899 ( .A1(n_747), .A2(n_43), .A3(n_41), .B(n_42), .Y(n_899) );
BUFx10_ASAP7_75t_L g900 ( .A(n_755), .Y(n_900) );
INVx3_ASAP7_75t_L g901 ( .A(n_730), .Y(n_901) );
AO31x2_ASAP7_75t_L g902 ( .A1(n_781), .A2(n_45), .A3(n_42), .B(n_44), .Y(n_902) );
INVx2_ASAP7_75t_L g903 ( .A(n_784), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_788), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_753), .Y(n_905) );
OR2x2_ASAP7_75t_L g906 ( .A(n_748), .B(n_45), .Y(n_906) );
BUFx2_ASAP7_75t_L g907 ( .A(n_729), .Y(n_907) );
AO31x2_ASAP7_75t_L g908 ( .A1(n_756), .A2(n_48), .A3(n_46), .B(n_47), .Y(n_908) );
NOR2xp33_ASAP7_75t_L g909 ( .A(n_761), .B(n_47), .Y(n_909) );
CKINVDCx5p33_ASAP7_75t_R g910 ( .A(n_763), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_768), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_767), .Y(n_912) );
BUFx6f_ASAP7_75t_L g913 ( .A(n_730), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_813), .B(n_48), .Y(n_914) );
AO31x2_ASAP7_75t_L g915 ( .A1(n_756), .A2(n_51), .A3(n_49), .B(n_50), .Y(n_915) );
INVx2_ASAP7_75t_SL g916 ( .A(n_819), .Y(n_916) );
CKINVDCx6p67_ASAP7_75t_R g917 ( .A(n_798), .Y(n_917) );
INVxp67_ASAP7_75t_SL g918 ( .A(n_726), .Y(n_918) );
OAI21xp5_ASAP7_75t_L g919 ( .A1(n_812), .A2(n_49), .B(n_52), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_799), .A2(n_55), .B1(n_52), .B2(n_53), .Y(n_920) );
A2O1A1Ixp33_ASAP7_75t_L g921 ( .A1(n_745), .A2(n_56), .B(n_53), .C(n_55), .Y(n_921) );
O2A1O1Ixp33_ASAP7_75t_L g922 ( .A1(n_775), .A2(n_58), .B(n_56), .C(n_57), .Y(n_922) );
O2A1O1Ixp33_ASAP7_75t_SL g923 ( .A1(n_805), .A2(n_238), .B(n_240), .C(n_236), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_778), .A2(n_60), .B1(n_58), .B2(n_59), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_774), .B(n_60), .Y(n_925) );
BUFx3_ASAP7_75t_L g926 ( .A(n_779), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_773), .Y(n_927) );
O2A1O1Ixp33_ASAP7_75t_SL g928 ( .A1(n_791), .A2(n_244), .B(n_245), .C(n_241), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_778), .A2(n_63), .B1(n_61), .B2(n_62), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_762), .Y(n_930) );
OA21x2_ASAP7_75t_L g931 ( .A1(n_810), .A2(n_248), .B(n_247), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_789), .Y(n_932) );
BUFx3_ASAP7_75t_L g933 ( .A(n_811), .Y(n_933) );
NOR2xp33_ASAP7_75t_SL g934 ( .A(n_749), .B(n_251), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_808), .Y(n_935) );
A2O1A1Ixp33_ASAP7_75t_L g936 ( .A1(n_811), .A2(n_63), .B(n_61), .C(n_62), .Y(n_936) );
NAND2x1p5_ASAP7_75t_L g937 ( .A(n_727), .B(n_64), .Y(n_937) );
NOR2xp33_ASAP7_75t_L g938 ( .A(n_770), .B(n_64), .Y(n_938) );
OR2x2_ASAP7_75t_L g939 ( .A(n_795), .B(n_65), .Y(n_939) );
OAI21x1_ASAP7_75t_SL g940 ( .A1(n_792), .A2(n_66), .B(n_67), .Y(n_940) );
AOI21xp5_ASAP7_75t_L g941 ( .A1(n_749), .A2(n_254), .B(n_253), .Y(n_941) );
AOI21xp5_ASAP7_75t_L g942 ( .A1(n_752), .A2(n_256), .B(n_255), .Y(n_942) );
AOI21xp5_ASAP7_75t_L g943 ( .A1(n_752), .A2(n_258), .B(n_257), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_806), .Y(n_944) );
BUFx2_ASAP7_75t_L g945 ( .A(n_786), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_791), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_727), .A2(n_70), .B1(n_67), .B2(n_68), .Y(n_947) );
BUFx2_ASAP7_75t_SL g948 ( .A(n_726), .Y(n_948) );
A2O1A1Ixp33_ASAP7_75t_L g949 ( .A1(n_726), .A2(n_72), .B(n_70), .C(n_71), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_728), .Y(n_950) );
AO31x2_ASAP7_75t_L g951 ( .A1(n_752), .A2(n_74), .A3(n_71), .B(n_73), .Y(n_951) );
INVx3_ASAP7_75t_L g952 ( .A(n_728), .Y(n_952) );
O2A1O1Ixp33_ASAP7_75t_L g953 ( .A1(n_794), .A2(n_77), .B(n_75), .C(n_76), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_794), .B(n_79), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_797), .B(n_80), .Y(n_955) );
CKINVDCx11_ASAP7_75t_R g956 ( .A(n_797), .Y(n_956) );
AOI221xp5_ASAP7_75t_L g957 ( .A1(n_735), .A2(n_81), .B1(n_82), .B2(n_83), .C(n_84), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_719), .Y(n_958) );
OAI21xp5_ASAP7_75t_L g959 ( .A1(n_825), .A2(n_262), .B(n_259), .Y(n_959) );
OAI21xp5_ASAP7_75t_L g960 ( .A1(n_825), .A2(n_265), .B(n_263), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_719), .B(n_81), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g962 ( .A1(n_723), .A2(n_86), .B1(n_83), .B2(n_85), .Y(n_962) );
AOI21xp33_ASAP7_75t_L g963 ( .A1(n_739), .A2(n_85), .B(n_86), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_723), .Y(n_964) );
AOI21xp5_ASAP7_75t_L g965 ( .A1(n_738), .A2(n_267), .B(n_266), .Y(n_965) );
AOI22xp5_ASAP7_75t_L g966 ( .A1(n_723), .A2(n_89), .B1(n_87), .B2(n_88), .Y(n_966) );
NAND2x1p5_ASAP7_75t_L g967 ( .A(n_723), .B(n_87), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_735), .A2(n_88), .B1(n_89), .B2(n_91), .C(n_93), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g969 ( .A(n_816), .B(n_94), .Y(n_969) );
AOI21xp5_ASAP7_75t_L g970 ( .A1(n_738), .A2(n_272), .B(n_271), .Y(n_970) );
OAI21x1_ASAP7_75t_L g971 ( .A1(n_802), .A2(n_276), .B(n_273), .Y(n_971) );
AOI21xp5_ASAP7_75t_L g972 ( .A1(n_859), .A2(n_279), .B(n_277), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_884), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_967), .A2(n_95), .B1(n_97), .B2(n_98), .Y(n_974) );
OR2x6_ASAP7_75t_L g975 ( .A(n_864), .B(n_97), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_830), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_969), .A2(n_99), .B1(n_100), .B2(n_101), .Y(n_977) );
OAI21xp5_ASAP7_75t_L g978 ( .A1(n_835), .A2(n_99), .B(n_100), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_896), .B(n_102), .Y(n_979) );
OR2x2_ASAP7_75t_L g980 ( .A(n_880), .B(n_103), .Y(n_980) );
INVx3_ASAP7_75t_L g981 ( .A(n_926), .Y(n_981) );
AOI222xp33_ASAP7_75t_L g982 ( .A1(n_911), .A2(n_104), .B1(n_106), .B2(n_107), .C1(n_108), .C2(n_109), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_832), .Y(n_983) );
AOI21xp5_ASAP7_75t_L g984 ( .A1(n_934), .A2(n_286), .B(n_284), .Y(n_984) );
BUFx2_ASAP7_75t_L g985 ( .A(n_887), .Y(n_985) );
OAI221xp5_ASAP7_75t_L g986 ( .A1(n_840), .A2(n_107), .B1(n_109), .B2(n_110), .C(n_111), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_888), .B(n_112), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_964), .Y(n_988) );
A2O1A1Ixp33_ASAP7_75t_L g989 ( .A1(n_860), .A2(n_114), .B(n_115), .C(n_117), .Y(n_989) );
AOI21xp33_ASAP7_75t_SL g990 ( .A1(n_910), .A2(n_115), .B(n_118), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_831), .B(n_119), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_861), .B(n_120), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_932), .B(n_120), .Y(n_993) );
AOI21xp33_ASAP7_75t_L g994 ( .A1(n_890), .A2(n_121), .B(n_122), .Y(n_994) );
AOI21xp5_ASAP7_75t_L g995 ( .A1(n_934), .A2(n_292), .B(n_289), .Y(n_995) );
AOI21xp5_ASAP7_75t_L g996 ( .A1(n_848), .A2(n_295), .B(n_294), .Y(n_996) );
OAI21xp5_ASAP7_75t_L g997 ( .A1(n_848), .A2(n_122), .B(n_124), .Y(n_997) );
NAND2xp5_ASAP7_75t_SL g998 ( .A(n_851), .B(n_124), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_961), .Y(n_999) );
INVx5_ASAP7_75t_L g1000 ( .A(n_913), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_958), .Y(n_1001) );
NAND2x1p5_ASAP7_75t_L g1002 ( .A(n_897), .B(n_125), .Y(n_1002) );
OAI21x1_ASAP7_75t_L g1003 ( .A1(n_971), .A2(n_301), .B(n_299), .Y(n_1003) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_967), .A2(n_125), .B1(n_126), .B2(n_127), .Y(n_1004) );
OA21x2_ASAP7_75t_L g1005 ( .A1(n_959), .A2(n_306), .B(n_305), .Y(n_1005) );
OA21x2_ASAP7_75t_L g1006 ( .A1(n_960), .A2(n_308), .B(n_307), .Y(n_1006) );
INVx1_ASAP7_75t_SL g1007 ( .A(n_897), .Y(n_1007) );
NAND3xp33_ASAP7_75t_L g1008 ( .A(n_869), .B(n_853), .C(n_873), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_843), .B(n_126), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_834), .A2(n_127), .B1(n_128), .B2(n_129), .Y(n_1010) );
AO21x2_ASAP7_75t_L g1011 ( .A1(n_865), .A2(n_309), .B(n_377), .Y(n_1011) );
AO21x2_ASAP7_75t_L g1012 ( .A1(n_865), .A2(n_376), .B(n_375), .Y(n_1012) );
INVx2_ASAP7_75t_L g1013 ( .A(n_856), .Y(n_1013) );
OAI22xp33_ASAP7_75t_L g1014 ( .A1(n_851), .A2(n_128), .B1(n_130), .B2(n_131), .Y(n_1014) );
BUFx3_ASAP7_75t_L g1015 ( .A(n_956), .Y(n_1015) );
OAI22x1_ASAP7_75t_L g1016 ( .A1(n_966), .A2(n_132), .B1(n_133), .B2(n_134), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_893), .B(n_134), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_837), .Y(n_1018) );
BUFx8_ASAP7_75t_L g1019 ( .A(n_855), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_836), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_904), .Y(n_1021) );
OA21x2_ASAP7_75t_L g1022 ( .A1(n_852), .A2(n_310), .B(n_373), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_878), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_863), .A2(n_135), .B1(n_136), .B2(n_137), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_882), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_903), .Y(n_1026) );
INVx3_ASAP7_75t_L g1027 ( .A(n_913), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_847), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_889), .Y(n_1029) );
AND2x4_ASAP7_75t_L g1030 ( .A(n_933), .B(n_138), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_920), .Y(n_1031) );
AOI21xp5_ASAP7_75t_L g1032 ( .A1(n_874), .A2(n_833), .B(n_894), .Y(n_1032) );
OAI21xp5_ASAP7_75t_L g1033 ( .A1(n_846), .A2(n_138), .B(n_139), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_902), .Y(n_1034) );
INVx4_ASAP7_75t_L g1035 ( .A(n_913), .Y(n_1035) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_886), .B(n_139), .Y(n_1036) );
HB1xp67_ASAP7_75t_L g1037 ( .A(n_937), .Y(n_1037) );
BUFx12f_ASAP7_75t_L g1038 ( .A(n_844), .Y(n_1038) );
AOI21x1_ASAP7_75t_L g1039 ( .A1(n_931), .A2(n_374), .B(n_367), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_927), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_909), .A2(n_141), .B1(n_142), .B2(n_144), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_935), .B(n_141), .Y(n_1042) );
INVx8_ASAP7_75t_L g1043 ( .A(n_875), .Y(n_1043) );
O2A1O1Ixp33_ASAP7_75t_L g1044 ( .A1(n_898), .A2(n_142), .B(n_144), .C(n_145), .Y(n_1044) );
INVx3_ASAP7_75t_L g1045 ( .A(n_875), .Y(n_1045) );
INVx4_ASAP7_75t_L g1046 ( .A(n_866), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_930), .B(n_148), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_966), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_938), .B(n_149), .Y(n_1049) );
OAI21xp5_ASAP7_75t_L g1050 ( .A1(n_846), .A2(n_845), .B(n_842), .Y(n_1050) );
AOI21xp5_ASAP7_75t_L g1051 ( .A1(n_928), .A2(n_312), .B(n_360), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_937), .Y(n_1052) );
BUFx8_ASAP7_75t_L g1053 ( .A(n_895), .Y(n_1053) );
CKINVDCx12_ASAP7_75t_R g1054 ( .A(n_867), .Y(n_1054) );
OA21x2_ASAP7_75t_L g1055 ( .A1(n_879), .A2(n_361), .B(n_359), .Y(n_1055) );
NOR2xp33_ASAP7_75t_L g1056 ( .A(n_886), .B(n_149), .Y(n_1056) );
AOI222xp33_ASAP7_75t_L g1057 ( .A1(n_957), .A2(n_150), .B1(n_151), .B2(n_152), .C1(n_153), .C2(n_154), .Y(n_1057) );
OA21x2_ASAP7_75t_L g1058 ( .A1(n_881), .A2(n_315), .B(n_357), .Y(n_1058) );
AOI21xp5_ASAP7_75t_L g1059 ( .A1(n_891), .A2(n_970), .B(n_965), .Y(n_1059) );
INVx3_ASAP7_75t_SL g1060 ( .A(n_885), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_828), .A2(n_152), .B1(n_153), .B2(n_155), .Y(n_1061) );
BUFx8_ASAP7_75t_SL g1062 ( .A(n_945), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_885), .B(n_155), .Y(n_1063) );
AO31x2_ASAP7_75t_L g1064 ( .A1(n_838), .A2(n_914), .A3(n_921), .B(n_883), .Y(n_1064) );
AOI21x1_ASAP7_75t_SL g1065 ( .A1(n_925), .A2(n_156), .B(n_158), .Y(n_1065) );
A2O1A1Ixp33_ASAP7_75t_L g1066 ( .A1(n_922), .A2(n_156), .B(n_160), .C(n_161), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_906), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_924), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_841), .A2(n_162), .B1(n_163), .B2(n_164), .Y(n_1069) );
CKINVDCx11_ASAP7_75t_R g1070 ( .A(n_900), .Y(n_1070) );
OAI221xp5_ASAP7_75t_L g1071 ( .A1(n_916), .A2(n_163), .B1(n_164), .B2(n_165), .C(n_167), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_900), .B(n_165), .Y(n_1072) );
OAI222xp33_ASAP7_75t_L g1073 ( .A1(n_962), .A2(n_167), .B1(n_169), .B2(n_170), .C1(n_171), .C2(n_172), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_841), .A2(n_169), .B1(n_170), .B2(n_171), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_907), .B(n_172), .Y(n_1075) );
INVx2_ASAP7_75t_L g1076 ( .A(n_905), .Y(n_1076) );
A2O1A1Ixp33_ASAP7_75t_L g1077 ( .A1(n_862), .A2(n_173), .B(n_174), .C(n_176), .Y(n_1077) );
AOI221xp5_ASAP7_75t_L g1078 ( .A1(n_963), .A2(n_173), .B1(n_174), .B2(n_176), .C(n_177), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_917), .B(n_178), .Y(n_1079) );
INVxp67_ASAP7_75t_L g1080 ( .A(n_868), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_850), .B(n_179), .Y(n_1081) );
NOR2xp33_ASAP7_75t_L g1082 ( .A(n_944), .B(n_180), .Y(n_1082) );
CKINVDCx5p33_ASAP7_75t_R g1083 ( .A(n_948), .Y(n_1083) );
AOI222xp33_ASAP7_75t_L g1084 ( .A1(n_968), .A2(n_181), .B1(n_182), .B2(n_183), .C1(n_184), .C2(n_185), .Y(n_1084) );
NOR2xp33_ASAP7_75t_L g1085 ( .A(n_849), .B(n_181), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_863), .A2(n_182), .B1(n_183), .B2(n_185), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_892), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_871), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_829), .B(n_186), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_899), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_850), .B(n_186), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_858), .B(n_187), .Y(n_1092) );
BUFx3_ASAP7_75t_L g1093 ( .A(n_901), .Y(n_1093) );
OA21x2_ASAP7_75t_L g1094 ( .A1(n_919), .A2(n_331), .B(n_356), .Y(n_1094) );
BUFx2_ASAP7_75t_L g1095 ( .A(n_946), .Y(n_1095) );
AOI21xp5_ASAP7_75t_L g1096 ( .A1(n_955), .A2(n_330), .B(n_354), .Y(n_1096) );
NAND3xp33_ASAP7_75t_L g1097 ( .A(n_872), .B(n_188), .C(n_189), .Y(n_1097) );
AOI22xp33_ASAP7_75t_SL g1098 ( .A1(n_940), .A2(n_190), .B1(n_191), .B2(n_192), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_939), .B(n_190), .Y(n_1099) );
AOI21xp5_ASAP7_75t_L g1100 ( .A1(n_923), .A2(n_335), .B(n_353), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_899), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_899), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_929), .B(n_191), .Y(n_1103) );
INVx2_ASAP7_75t_L g1104 ( .A(n_912), .Y(n_1104) );
INVx1_ASAP7_75t_SL g1105 ( .A(n_952), .Y(n_1105) );
OAI22xp33_ASAP7_75t_L g1106 ( .A1(n_877), .A2(n_194), .B1(n_195), .B2(n_196), .Y(n_1106) );
AOI21xp5_ASAP7_75t_L g1107 ( .A1(n_876), .A2(n_338), .B(n_351), .Y(n_1107) );
OAI221xp5_ASAP7_75t_L g1108 ( .A1(n_857), .A2(n_194), .B1(n_195), .B2(n_197), .C(n_198), .Y(n_1108) );
AND2x4_ASAP7_75t_L g1109 ( .A(n_901), .B(n_952), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_870), .Y(n_1110) );
AOI21xp33_ASAP7_75t_L g1111 ( .A1(n_953), .A2(n_316), .B(n_317), .Y(n_1111) );
AOI21xp5_ASAP7_75t_L g1112 ( .A1(n_931), .A2(n_319), .B(n_322), .Y(n_1112) );
AOI21xp5_ASAP7_75t_L g1113 ( .A1(n_941), .A2(n_325), .B(n_327), .Y(n_1113) );
AOI21xp5_ASAP7_75t_L g1114 ( .A1(n_918), .A2(n_329), .B(n_341), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_936), .Y(n_1115) );
OAI21xp5_ASAP7_75t_L g1116 ( .A1(n_954), .A2(n_943), .B(n_942), .Y(n_1116) );
AO21x2_ASAP7_75t_L g1117 ( .A1(n_949), .A2(n_342), .B(n_343), .Y(n_1117) );
INVx2_ASAP7_75t_L g1118 ( .A(n_950), .Y(n_1118) );
OR2x6_ASAP7_75t_L g1119 ( .A(n_947), .B(n_344), .Y(n_1119) );
AOI21xp5_ASAP7_75t_L g1120 ( .A1(n_839), .A2(n_345), .B(n_347), .Y(n_1120) );
CKINVDCx20_ASAP7_75t_R g1121 ( .A(n_1062), .Y(n_1121) );
OAI221xp5_ASAP7_75t_L g1122 ( .A1(n_1080), .A2(n_951), .B1(n_839), .B2(n_908), .C(n_915), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1029), .B(n_975), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_973), .Y(n_1124) );
AOI33xp33_ASAP7_75t_L g1125 ( .A1(n_1067), .A2(n_951), .A3(n_915), .B1(n_908), .B2(n_839), .B3(n_854), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1013), .B(n_908), .Y(n_1126) );
INVx2_ASAP7_75t_L g1127 ( .A(n_983), .Y(n_1127) );
INVx2_ASAP7_75t_L g1128 ( .A(n_988), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1021), .Y(n_1129) );
NOR2xp33_ASAP7_75t_L g1130 ( .A(n_1028), .B(n_348), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_976), .B(n_915), .Y(n_1131) );
OAI21xp5_ASAP7_75t_L g1132 ( .A1(n_1008), .A2(n_854), .B(n_349), .Y(n_1132) );
HB1xp67_ASAP7_75t_L g1133 ( .A(n_1007), .Y(n_1133) );
INVx4_ASAP7_75t_L g1134 ( .A(n_1000), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1040), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1023), .B(n_1025), .Y(n_1136) );
AOI22xp5_ASAP7_75t_L g1137 ( .A1(n_1054), .A2(n_975), .B1(n_1081), .B2(n_1091), .Y(n_1137) );
BUFx6f_ASAP7_75t_L g1138 ( .A(n_1000), .Y(n_1138) );
BUFx2_ASAP7_75t_L g1139 ( .A(n_1083), .Y(n_1139) );
INVx3_ASAP7_75t_L g1140 ( .A(n_1000), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1026), .Y(n_1141) );
OA21x2_ASAP7_75t_L g1142 ( .A1(n_1101), .A2(n_1102), .B(n_1034), .Y(n_1142) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_980), .B(n_1060), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1076), .B(n_1104), .Y(n_1144) );
OR2x2_ASAP7_75t_L g1145 ( .A(n_975), .B(n_1047), .Y(n_1145) );
OR2x6_ASAP7_75t_L g1146 ( .A(n_1002), .B(n_1119), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_981), .B(n_1095), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1088), .B(n_978), .Y(n_1148) );
OA21x2_ASAP7_75t_L g1149 ( .A1(n_1087), .A2(n_1120), .B(n_1032), .Y(n_1149) );
OR2x6_ASAP7_75t_L g1150 ( .A(n_1002), .B(n_1119), .Y(n_1150) );
OA21x2_ASAP7_75t_L g1151 ( .A1(n_1112), .A2(n_1059), .B(n_1050), .Y(n_1151) );
OR2x6_ASAP7_75t_L g1152 ( .A(n_1119), .B(n_1037), .Y(n_1152) );
BUFx6f_ASAP7_75t_L g1153 ( .A(n_1035), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1001), .Y(n_1154) );
OAI222xp33_ASAP7_75t_L g1155 ( .A1(n_974), .A2(n_1004), .B1(n_1024), .B2(n_1086), .C1(n_1110), .C2(n_1071), .Y(n_1155) );
AND2x4_ASAP7_75t_L g1156 ( .A(n_1052), .B(n_1007), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1031), .B(n_1099), .Y(n_1157) );
OR2x2_ASAP7_75t_L g1158 ( .A(n_1075), .B(n_1030), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_979), .Y(n_1159) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1055), .Y(n_1160) );
INVx1_ASAP7_75t_SL g1161 ( .A(n_1070), .Y(n_1161) );
OR2x6_ASAP7_75t_L g1162 ( .A(n_974), .B(n_1004), .Y(n_1162) );
BUFx3_ASAP7_75t_L g1163 ( .A(n_1038), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_999), .B(n_992), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_993), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1082), .Y(n_1166) );
AND2x4_ASAP7_75t_L g1167 ( .A(n_1035), .B(n_1109), .Y(n_1167) );
BUFx6f_ASAP7_75t_L g1168 ( .A(n_1027), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1063), .Y(n_1169) );
HB1xp67_ASAP7_75t_L g1170 ( .A(n_1105), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1042), .Y(n_1171) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1055), .Y(n_1172) );
INVx2_ASAP7_75t_L g1173 ( .A(n_1058), .Y(n_1173) );
INVx2_ASAP7_75t_L g1174 ( .A(n_1058), .Y(n_1174) );
CKINVDCx8_ASAP7_75t_R g1175 ( .A(n_985), .Y(n_1175) );
BUFx3_ASAP7_75t_L g1176 ( .A(n_1043), .Y(n_1176) );
OA21x2_ASAP7_75t_L g1177 ( .A1(n_1050), .A2(n_1051), .B(n_1116), .Y(n_1177) );
INVx2_ASAP7_75t_SL g1178 ( .A(n_1043), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1030), .B(n_982), .Y(n_1179) );
OA21x2_ASAP7_75t_L g1180 ( .A1(n_1116), .A2(n_1008), .B(n_1003), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_987), .Y(n_1181) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1094), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_991), .B(n_1017), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1118), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1185 ( .A(n_1072), .B(n_1049), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_978), .B(n_1033), .Y(n_1186) );
AO21x2_ASAP7_75t_L g1187 ( .A1(n_997), .A2(n_1111), .B(n_1048), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_1085), .B(n_1068), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1016), .Y(n_1189) );
OR2x6_ASAP7_75t_L g1190 ( .A(n_1033), .B(n_1043), .Y(n_1190) );
BUFx2_ASAP7_75t_L g1191 ( .A(n_1019), .Y(n_1191) );
NOR2xp33_ASAP7_75t_L g1192 ( .A(n_1046), .B(n_1092), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1036), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1115), .B(n_1018), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1094), .Y(n_1195) );
INVx1_ASAP7_75t_SL g1196 ( .A(n_1015), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1057), .B(n_1084), .Y(n_1197) );
INVx3_ASAP7_75t_L g1198 ( .A(n_1027), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1056), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1057), .B(n_1084), .Y(n_1200) );
OA21x2_ASAP7_75t_L g1201 ( .A1(n_1100), .A2(n_1097), .B(n_996), .Y(n_1201) );
OR2x2_ASAP7_75t_L g1202 ( .A(n_1093), .B(n_1079), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1103), .B(n_1109), .Y(n_1203) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1011), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1045), .B(n_1064), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1045), .B(n_1064), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_986), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1009), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1046), .B(n_994), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1064), .B(n_1086), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1041), .B(n_1010), .Y(n_1211) );
OAI321xp33_ASAP7_75t_L g1212 ( .A1(n_1024), .A2(n_1014), .A3(n_1097), .B1(n_1108), .B2(n_1106), .C(n_977), .Y(n_1212) );
INVx2_ASAP7_75t_L g1213 ( .A(n_1012), .Y(n_1213) );
OR2x6_ASAP7_75t_L g1214 ( .A(n_984), .B(n_995), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1089), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_1061), .A2(n_1098), .B1(n_1069), .B2(n_1074), .Y(n_1216) );
OAI21xp5_ASAP7_75t_L g1217 ( .A1(n_989), .A2(n_1066), .B(n_1077), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_998), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_994), .B(n_1105), .Y(n_1219) );
INVxp67_ASAP7_75t_L g1220 ( .A(n_1019), .Y(n_1220) );
OR2x6_ASAP7_75t_L g1221 ( .A(n_1020), .B(n_1044), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1078), .Y(n_1222) );
HB1xp67_ASAP7_75t_L g1223 ( .A(n_1117), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_990), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1005), .B(n_1006), .Y(n_1225) );
BUFx2_ASAP7_75t_L g1226 ( .A(n_1053), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1053), .Y(n_1227) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1022), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1005), .B(n_1006), .Y(n_1229) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1022), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1096), .B(n_1114), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_972), .B(n_1113), .Y(n_1232) );
INVx3_ASAP7_75t_L g1233 ( .A(n_1065), .Y(n_1233) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1073), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1107), .B(n_980), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1013), .B(n_1023), .Y(n_1236) );
BUFx2_ASAP7_75t_L g1237 ( .A(n_1083), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_1088), .A2(n_670), .B1(n_816), .B2(n_711), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_973), .Y(n_1239) );
INVx3_ASAP7_75t_L g1240 ( .A(n_1000), .Y(n_1240) );
OR2x6_ASAP7_75t_L g1241 ( .A(n_975), .B(n_967), .Y(n_1241) );
AOI21x1_ASAP7_75t_L g1242 ( .A1(n_1039), .A2(n_1101), .B(n_1090), .Y(n_1242) );
INVxp67_ASAP7_75t_SL g1243 ( .A(n_1037), .Y(n_1243) );
OAI222xp33_ASAP7_75t_L g1244 ( .A1(n_975), .A2(n_670), .B1(n_967), .B2(n_1004), .C1(n_974), .C2(n_1002), .Y(n_1244) );
INVx2_ASAP7_75t_SL g1245 ( .A(n_1000), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_973), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_973), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_973), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1013), .B(n_1023), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_973), .Y(n_1250) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1142), .Y(n_1251) );
AND2x4_ASAP7_75t_L g1252 ( .A(n_1205), .B(n_1206), .Y(n_1252) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1142), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1210), .B(n_1205), .Y(n_1254) );
HB1xp67_ASAP7_75t_L g1255 ( .A(n_1133), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1210), .B(n_1206), .Y(n_1256) );
INVx3_ASAP7_75t_L g1257 ( .A(n_1152), .Y(n_1257) );
INVx1_ASAP7_75t_SL g1258 ( .A(n_1139), .Y(n_1258) );
HB1xp67_ASAP7_75t_L g1259 ( .A(n_1133), .Y(n_1259) );
BUFx2_ASAP7_75t_L g1260 ( .A(n_1152), .Y(n_1260) );
BUFx2_ASAP7_75t_L g1261 ( .A(n_1152), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1126), .B(n_1136), .Y(n_1262) );
NOR2xp33_ASAP7_75t_L g1263 ( .A(n_1145), .B(n_1192), .Y(n_1263) );
NAND4xp25_ASAP7_75t_L g1264 ( .A(n_1188), .B(n_1137), .C(n_1238), .D(n_1179), .Y(n_1264) );
AND2x4_ASAP7_75t_L g1265 ( .A(n_1152), .B(n_1126), .Y(n_1265) );
AND2x4_ASAP7_75t_L g1266 ( .A(n_1146), .B(n_1150), .Y(n_1266) );
INVxp67_ASAP7_75t_L g1267 ( .A(n_1237), .Y(n_1267) );
INVx1_ASAP7_75t_SL g1268 ( .A(n_1191), .Y(n_1268) );
INVx4_ASAP7_75t_L g1269 ( .A(n_1146), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1131), .Y(n_1270) );
INVx3_ASAP7_75t_L g1271 ( .A(n_1146), .Y(n_1271) );
INVxp67_ASAP7_75t_L g1272 ( .A(n_1143), .Y(n_1272) );
AND2x4_ASAP7_75t_L g1273 ( .A(n_1146), .B(n_1150), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1274 ( .A(n_1162), .B(n_1157), .Y(n_1274) );
BUFx3_ASAP7_75t_L g1275 ( .A(n_1176), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1236), .B(n_1249), .Y(n_1276) );
BUFx3_ASAP7_75t_L g1277 ( .A(n_1176), .Y(n_1277) );
INVx4_ASAP7_75t_R g1278 ( .A(n_1163), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1136), .B(n_1148), .Y(n_1279) );
OR2x6_ASAP7_75t_L g1280 ( .A(n_1150), .B(n_1162), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1148), .B(n_1236), .Y(n_1281) );
BUFx3_ASAP7_75t_L g1282 ( .A(n_1138), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1249), .B(n_1144), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1242), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1200), .B(n_1124), .Y(n_1285) );
INVx2_ASAP7_75t_L g1286 ( .A(n_1127), .Y(n_1286) );
OAI211xp5_ASAP7_75t_SL g1287 ( .A1(n_1166), .A2(n_1164), .B(n_1175), .C(n_1185), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1128), .B(n_1194), .Y(n_1288) );
INVxp67_ASAP7_75t_L g1289 ( .A(n_1243), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_1170), .B(n_1150), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1194), .Y(n_1291) );
AND2x4_ASAP7_75t_L g1292 ( .A(n_1190), .B(n_1156), .Y(n_1292) );
BUFx3_ASAP7_75t_L g1293 ( .A(n_1138), .Y(n_1293) );
OR2x2_ASAP7_75t_L g1294 ( .A(n_1170), .B(n_1189), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1135), .B(n_1129), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1125), .Y(n_1296) );
AND2x4_ASAP7_75t_L g1297 ( .A(n_1190), .B(n_1156), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1125), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1239), .B(n_1246), .Y(n_1299) );
AND2x4_ASAP7_75t_L g1300 ( .A(n_1190), .B(n_1156), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1169), .B(n_1181), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1154), .Y(n_1302) );
OAI221xp5_ASAP7_75t_L g1303 ( .A1(n_1238), .A2(n_1197), .B1(n_1224), .B2(n_1209), .C(n_1193), .Y(n_1303) );
NAND2xp33_ASAP7_75t_R g1304 ( .A(n_1226), .B(n_1241), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1247), .B(n_1248), .Y(n_1305) );
BUFx2_ASAP7_75t_L g1306 ( .A(n_1241), .Y(n_1306) );
INVx4_ASAP7_75t_L g1307 ( .A(n_1241), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1250), .B(n_1141), .Y(n_1308) );
AND2x4_ASAP7_75t_L g1309 ( .A(n_1190), .B(n_1219), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1184), .B(n_1219), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1186), .B(n_1203), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1186), .B(n_1203), .Y(n_1312) );
OR2x2_ASAP7_75t_L g1313 ( .A(n_1147), .B(n_1158), .Y(n_1313) );
NAND4xp25_ASAP7_75t_L g1314 ( .A(n_1200), .B(n_1123), .C(n_1199), .D(n_1192), .Y(n_1314) );
AND2x4_ASAP7_75t_L g1315 ( .A(n_1241), .B(n_1153), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1180), .B(n_1171), .Y(n_1316) );
INVx4_ASAP7_75t_L g1317 ( .A(n_1138), .Y(n_1317) );
INVx3_ASAP7_75t_L g1318 ( .A(n_1153), .Y(n_1318) );
AND2x4_ASAP7_75t_L g1319 ( .A(n_1153), .B(n_1167), .Y(n_1319) );
AND2x4_ASAP7_75t_L g1320 ( .A(n_1153), .B(n_1167), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1159), .B(n_1165), .Y(n_1321) );
HB1xp67_ASAP7_75t_L g1322 ( .A(n_1245), .Y(n_1322) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_1207), .A2(n_1234), .B1(n_1216), .B2(n_1211), .Y(n_1323) );
HB1xp67_ASAP7_75t_L g1324 ( .A(n_1245), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1180), .B(n_1234), .Y(n_1325) );
HB1xp67_ASAP7_75t_L g1326 ( .A(n_1138), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1183), .B(n_1215), .Y(n_1327) );
CKINVDCx10_ASAP7_75t_R g1328 ( .A(n_1121), .Y(n_1328) );
OR2x2_ASAP7_75t_L g1329 ( .A(n_1202), .B(n_1208), .Y(n_1329) );
OAI221xp5_ASAP7_75t_L g1330 ( .A1(n_1222), .A2(n_1217), .B1(n_1235), .B2(n_1175), .C(n_1221), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1187), .B(n_1177), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1177), .B(n_1151), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1130), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1177), .B(n_1151), .Y(n_1334) );
AOI22xp33_ASAP7_75t_L g1335 ( .A1(n_1221), .A2(n_1130), .B1(n_1218), .B2(n_1233), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1140), .Y(n_1336) );
AND2x2_ASAP7_75t_SL g1337 ( .A(n_1244), .B(n_1134), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1299), .Y(n_1338) );
INVx3_ASAP7_75t_SL g1339 ( .A(n_1275), .Y(n_1339) );
NOR2x1_ASAP7_75t_L g1340 ( .A(n_1275), .B(n_1277), .Y(n_1340) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_1283), .B(n_1167), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1342 ( .A(n_1279), .B(n_1196), .Y(n_1342) );
AND2x4_ASAP7_75t_L g1343 ( .A(n_1252), .B(n_1223), .Y(n_1343) );
AND2x4_ASAP7_75t_SL g1344 ( .A(n_1307), .B(n_1134), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1305), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1308), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1254), .B(n_1223), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1308), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1283), .B(n_1227), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1254), .B(n_1213), .Y(n_1350) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1251), .Y(n_1351) );
NOR2xp33_ASAP7_75t_L g1352 ( .A(n_1264), .B(n_1155), .Y(n_1352) );
OR2x2_ASAP7_75t_L g1353 ( .A(n_1279), .B(n_1161), .Y(n_1353) );
NOR2x1_ASAP7_75t_L g1354 ( .A(n_1277), .B(n_1121), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1256), .B(n_1204), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1291), .B(n_1140), .Y(n_1356) );
OR2x2_ASAP7_75t_L g1357 ( .A(n_1281), .B(n_1240), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1256), .B(n_1213), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1302), .Y(n_1359) );
INVx2_ASAP7_75t_L g1360 ( .A(n_1251), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1262), .B(n_1204), .Y(n_1361) );
NAND2x1p5_ASAP7_75t_L g1362 ( .A(n_1317), .B(n_1134), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1262), .B(n_1149), .Y(n_1363) );
NAND2xp5_ASAP7_75t_L g1364 ( .A(n_1291), .B(n_1240), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1295), .Y(n_1365) );
OR2x2_ASAP7_75t_L g1366 ( .A(n_1313), .B(n_1198), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1311), .B(n_1149), .Y(n_1367) );
NOR2x1_ASAP7_75t_L g1368 ( .A(n_1317), .B(n_1163), .Y(n_1368) );
NOR2x1_ASAP7_75t_L g1369 ( .A(n_1317), .B(n_1233), .Y(n_1369) );
NOR2xp67_ASAP7_75t_L g1370 ( .A(n_1314), .B(n_1220), .Y(n_1370) );
INVx1_ASAP7_75t_SL g1371 ( .A(n_1268), .Y(n_1371) );
OR2x2_ASAP7_75t_L g1372 ( .A(n_1313), .B(n_1198), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1312), .B(n_1198), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1252), .B(n_1195), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1252), .B(n_1195), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1310), .B(n_1182), .Y(n_1376) );
NOR3xp33_ASAP7_75t_SL g1377 ( .A(n_1304), .B(n_1212), .C(n_1122), .Y(n_1377) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1295), .Y(n_1378) );
OR2x2_ASAP7_75t_L g1379 ( .A(n_1276), .B(n_1178), .Y(n_1379) );
NAND2xp5_ASAP7_75t_L g1380 ( .A(n_1288), .B(n_1221), .Y(n_1380) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1288), .B(n_1221), .Y(n_1381) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1301), .Y(n_1382) );
AND2x4_ASAP7_75t_SL g1383 ( .A(n_1307), .B(n_1168), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1301), .Y(n_1384) );
INVxp67_ASAP7_75t_SL g1385 ( .A(n_1253), .Y(n_1385) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1316), .B(n_1225), .Y(n_1386) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1294), .Y(n_1387) );
BUFx3_ASAP7_75t_L g1388 ( .A(n_1282), .Y(n_1388) );
NAND2xp5_ASAP7_75t_L g1389 ( .A(n_1285), .B(n_1178), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1294), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1329), .Y(n_1391) );
OR2x2_ASAP7_75t_L g1392 ( .A(n_1274), .B(n_1168), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1316), .B(n_1225), .Y(n_1393) );
HB1xp67_ASAP7_75t_L g1394 ( .A(n_1255), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1325), .B(n_1173), .Y(n_1395) );
NAND5xp2_ASAP7_75t_L g1396 ( .A(n_1330), .B(n_1323), .C(n_1335), .D(n_1303), .E(n_1306), .Y(n_1396) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1329), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1325), .B(n_1173), .Y(n_1398) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1259), .Y(n_1399) );
OR2x2_ASAP7_75t_L g1400 ( .A(n_1274), .B(n_1168), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1309), .B(n_1172), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1309), .B(n_1172), .Y(n_1402) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1321), .Y(n_1403) );
OR2x2_ASAP7_75t_L g1404 ( .A(n_1289), .B(n_1228), .Y(n_1404) );
HB1xp67_ASAP7_75t_L g1405 ( .A(n_1286), .Y(n_1405) );
INVx1_ASAP7_75t_SL g1406 ( .A(n_1258), .Y(n_1406) );
OR2x2_ASAP7_75t_L g1407 ( .A(n_1272), .B(n_1230), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1309), .B(n_1160), .Y(n_1408) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1265), .B(n_1174), .Y(n_1409) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1322), .Y(n_1410) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1324), .Y(n_1411) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_1265), .B(n_1174), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1265), .B(n_1229), .Y(n_1413) );
NAND2x1_ASAP7_75t_SL g1414 ( .A(n_1266), .B(n_1231), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_1386), .B(n_1280), .Y(n_1415) );
NAND2xp5_ASAP7_75t_SL g1416 ( .A(n_1370), .B(n_1337), .Y(n_1416) );
INVx2_ASAP7_75t_SL g1417 ( .A(n_1339), .Y(n_1417) );
INVxp67_ASAP7_75t_L g1418 ( .A(n_1394), .Y(n_1418) );
OR2x2_ASAP7_75t_L g1419 ( .A(n_1357), .B(n_1290), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1386), .B(n_1280), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1373), .B(n_1280), .Y(n_1421) );
NOR2xp33_ASAP7_75t_L g1422 ( .A(n_1352), .B(n_1396), .Y(n_1422) );
NAND2xp5_ASAP7_75t_L g1423 ( .A(n_1338), .B(n_1327), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1342), .B(n_1413), .Y(n_1424) );
INVx2_ASAP7_75t_SL g1425 ( .A(n_1339), .Y(n_1425) );
NOR2xp33_ASAP7_75t_L g1426 ( .A(n_1352), .B(n_1287), .Y(n_1426) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1351), .Y(n_1427) );
AND3x2_ASAP7_75t_L g1428 ( .A(n_1410), .B(n_1306), .C(n_1260), .Y(n_1428) );
INVx2_ASAP7_75t_L g1429 ( .A(n_1351), .Y(n_1429) );
INVx2_ASAP7_75t_L g1430 ( .A(n_1360), .Y(n_1430) );
BUFx2_ASAP7_75t_L g1431 ( .A(n_1340), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1359), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1393), .B(n_1280), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1413), .B(n_1263), .Y(n_1434) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1391), .B(n_1270), .Y(n_1435) );
INVx4_ASAP7_75t_L g1436 ( .A(n_1344), .Y(n_1436) );
INVx2_ASAP7_75t_SL g1437 ( .A(n_1388), .Y(n_1437) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1387), .Y(n_1438) );
AND2x4_ASAP7_75t_L g1439 ( .A(n_1343), .B(n_1266), .Y(n_1439) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_1345), .B(n_1296), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1397), .B(n_1266), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1393), .B(n_1298), .Y(n_1442) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1390), .Y(n_1443) );
AOI22xp5_ASAP7_75t_L g1444 ( .A1(n_1377), .A2(n_1273), .B1(n_1269), .B2(n_1307), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1399), .Y(n_1445) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1382), .Y(n_1446) );
OR2x2_ASAP7_75t_L g1447 ( .A(n_1346), .B(n_1273), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1348), .B(n_1333), .Y(n_1448) );
OR2x2_ASAP7_75t_L g1449 ( .A(n_1384), .B(n_1273), .Y(n_1449) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1365), .Y(n_1450) );
OR2x2_ASAP7_75t_L g1451 ( .A(n_1378), .B(n_1292), .Y(n_1451) );
OR2x2_ASAP7_75t_L g1452 ( .A(n_1341), .B(n_1292), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1350), .B(n_1332), .Y(n_1453) );
OR2x2_ASAP7_75t_L g1454 ( .A(n_1407), .B(n_1292), .Y(n_1454) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1353), .B(n_1297), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1403), .B(n_1271), .Y(n_1456) );
OR2x2_ASAP7_75t_L g1457 ( .A(n_1366), .B(n_1297), .Y(n_1457) );
OR2x2_ASAP7_75t_L g1458 ( .A(n_1372), .B(n_1297), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1411), .B(n_1300), .Y(n_1459) );
NAND2x1p5_ASAP7_75t_L g1460 ( .A(n_1368), .B(n_1269), .Y(n_1460) );
INVxp67_ASAP7_75t_SL g1461 ( .A(n_1405), .Y(n_1461) );
OR2x2_ASAP7_75t_L g1462 ( .A(n_1349), .B(n_1361), .Y(n_1462) );
NAND2xp5_ASAP7_75t_L g1463 ( .A(n_1356), .B(n_1271), .Y(n_1463) );
INVx1_ASAP7_75t_SL g1464 ( .A(n_1371), .Y(n_1464) );
INVx2_ASAP7_75t_SL g1465 ( .A(n_1388), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1466 ( .A(n_1364), .B(n_1271), .Y(n_1466) );
OR2x2_ASAP7_75t_L g1467 ( .A(n_1361), .B(n_1300), .Y(n_1467) );
OAI21xp33_ASAP7_75t_L g1468 ( .A1(n_1422), .A2(n_1377), .B(n_1414), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1424), .B(n_1347), .Y(n_1469) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1432), .Y(n_1470) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1442), .B(n_1363), .Y(n_1471) );
NAND2xp5_ASAP7_75t_SL g1472 ( .A(n_1436), .B(n_1354), .Y(n_1472) );
NAND2xp5_ASAP7_75t_L g1473 ( .A(n_1442), .B(n_1363), .Y(n_1473) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_1422), .A2(n_1389), .B1(n_1269), .B2(n_1379), .Y(n_1474) );
NAND2xp5_ASAP7_75t_SL g1475 ( .A(n_1436), .B(n_1406), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1453), .B(n_1367), .Y(n_1476) );
NAND2xp5_ASAP7_75t_L g1477 ( .A(n_1440), .B(n_1347), .Y(n_1477) );
NAND2xp33_ASAP7_75t_L g1478 ( .A(n_1417), .B(n_1362), .Y(n_1478) );
INVx2_ASAP7_75t_SL g1479 ( .A(n_1417), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1453), .B(n_1350), .Y(n_1480) );
HB1xp67_ASAP7_75t_L g1481 ( .A(n_1418), .Y(n_1481) );
OR2x2_ASAP7_75t_L g1482 ( .A(n_1462), .B(n_1355), .Y(n_1482) );
OAI21xp5_ASAP7_75t_L g1483 ( .A1(n_1426), .A2(n_1267), .B(n_1362), .Y(n_1483) );
AOI22xp5_ASAP7_75t_L g1484 ( .A1(n_1426), .A2(n_1380), .B1(n_1381), .B2(n_1343), .Y(n_1484) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1415), .B(n_1358), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1486 ( .A(n_1415), .B(n_1358), .Y(n_1486) );
INVx2_ASAP7_75t_L g1487 ( .A(n_1427), .Y(n_1487) );
AOI21xp33_ASAP7_75t_SL g1488 ( .A1(n_1425), .A2(n_1278), .B(n_1328), .Y(n_1488) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1450), .B(n_1376), .Y(n_1489) );
NAND2xp5_ASAP7_75t_L g1490 ( .A(n_1438), .B(n_1395), .Y(n_1490) );
AOI22xp33_ASAP7_75t_L g1491 ( .A1(n_1416), .A2(n_1260), .B1(n_1261), .B2(n_1300), .Y(n_1491) );
NAND2xp5_ASAP7_75t_L g1492 ( .A(n_1443), .B(n_1395), .Y(n_1492) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1445), .Y(n_1493) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1435), .Y(n_1494) );
OR2x6_ASAP7_75t_L g1495 ( .A(n_1436), .B(n_1261), .Y(n_1495) );
NAND2xp5_ASAP7_75t_L g1496 ( .A(n_1446), .B(n_1398), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1497 ( .A(n_1419), .B(n_1404), .Y(n_1497) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1448), .Y(n_1498) );
NAND2xp5_ASAP7_75t_L g1499 ( .A(n_1498), .B(n_1434), .Y(n_1499) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1481), .Y(n_1500) );
NOR2xp33_ASAP7_75t_L g1501 ( .A(n_1468), .B(n_1464), .Y(n_1501) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1470), .Y(n_1502) );
O2A1O1Ixp33_ASAP7_75t_L g1503 ( .A1(n_1488), .A2(n_1431), .B(n_1423), .C(n_1456), .Y(n_1503) );
AOI22xp5_ASAP7_75t_L g1504 ( .A1(n_1475), .A2(n_1420), .B1(n_1433), .B2(n_1459), .Y(n_1504) );
OR2x2_ASAP7_75t_L g1505 ( .A(n_1482), .B(n_1461), .Y(n_1505) );
AOI22xp33_ASAP7_75t_L g1506 ( .A1(n_1474), .A2(n_1441), .B1(n_1343), .B2(n_1433), .Y(n_1506) );
INVx2_ASAP7_75t_L g1507 ( .A(n_1487), .Y(n_1507) );
NAND2xp5_ASAP7_75t_L g1508 ( .A(n_1480), .B(n_1455), .Y(n_1508) );
NOR2xp33_ASAP7_75t_L g1509 ( .A(n_1479), .B(n_1452), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1476), .B(n_1374), .Y(n_1510) );
OR2x2_ASAP7_75t_L g1511 ( .A(n_1471), .B(n_1467), .Y(n_1511) );
AOI22xp5_ASAP7_75t_L g1512 ( .A1(n_1484), .A2(n_1444), .B1(n_1439), .B2(n_1421), .Y(n_1512) );
NAND2xp5_ASAP7_75t_L g1513 ( .A(n_1480), .B(n_1437), .Y(n_1513) );
AOI21xp33_ASAP7_75t_L g1514 ( .A1(n_1483), .A2(n_1437), .B(n_1465), .Y(n_1514) );
OAI21xp5_ASAP7_75t_L g1515 ( .A1(n_1472), .A2(n_1460), .B(n_1465), .Y(n_1515) );
NAND2xp5_ASAP7_75t_L g1516 ( .A(n_1477), .B(n_1451), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_1473), .B(n_1449), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_1469), .B(n_1374), .Y(n_1518) );
OA22x2_ASAP7_75t_L g1519 ( .A1(n_1515), .A2(n_1495), .B1(n_1479), .B2(n_1428), .Y(n_1519) );
NAND2xp5_ASAP7_75t_L g1520 ( .A(n_1500), .B(n_1494), .Y(n_1520) );
AOI21xp5_ASAP7_75t_L g1521 ( .A1(n_1503), .A2(n_1478), .B(n_1495), .Y(n_1521) );
NAND3xp33_ASAP7_75t_L g1522 ( .A(n_1501), .B(n_1491), .C(n_1478), .Y(n_1522) );
OAI211xp5_ASAP7_75t_L g1523 ( .A1(n_1514), .A2(n_1491), .B(n_1257), .C(n_1369), .Y(n_1523) );
OAI21xp5_ASAP7_75t_SL g1524 ( .A1(n_1506), .A2(n_1460), .B(n_1428), .Y(n_1524) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1502), .Y(n_1525) );
A2O1A1Ixp33_ASAP7_75t_L g1526 ( .A1(n_1509), .A2(n_1344), .B(n_1439), .C(n_1497), .Y(n_1526) );
OAI21xp5_ASAP7_75t_SL g1527 ( .A1(n_1512), .A2(n_1439), .B(n_1315), .Y(n_1527) );
OAI21xp5_ASAP7_75t_L g1528 ( .A1(n_1509), .A2(n_1495), .B(n_1493), .Y(n_1528) );
BUFx3_ASAP7_75t_L g1529 ( .A(n_1513), .Y(n_1529) );
OAI21xp33_ASAP7_75t_L g1530 ( .A1(n_1504), .A2(n_1496), .B(n_1492), .Y(n_1530) );
AOI222xp33_ASAP7_75t_L g1531 ( .A1(n_1499), .A2(n_1490), .B1(n_1489), .B2(n_1486), .C1(n_1485), .C2(n_1463), .Y(n_1531) );
OAI22xp5_ASAP7_75t_L g1532 ( .A1(n_1505), .A2(n_1495), .B1(n_1486), .B2(n_1454), .Y(n_1532) );
OAI211xp5_ASAP7_75t_L g1533 ( .A1(n_1521), .A2(n_1257), .B(n_1326), .C(n_1282), .Y(n_1533) );
OAI222xp33_ASAP7_75t_L g1534 ( .A1(n_1519), .A2(n_1511), .B1(n_1508), .B2(n_1516), .C1(n_1517), .C2(n_1447), .Y(n_1534) );
AOI221xp5_ASAP7_75t_SL g1535 ( .A1(n_1528), .A2(n_1510), .B1(n_1518), .B2(n_1466), .C(n_1507), .Y(n_1535) );
AOI221xp5_ASAP7_75t_L g1536 ( .A1(n_1527), .A2(n_1375), .B1(n_1336), .B2(n_1402), .C(n_1401), .Y(n_1536) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1520), .Y(n_1537) );
NAND2xp5_ASAP7_75t_L g1538 ( .A(n_1531), .B(n_1331), .Y(n_1538) );
OAI22xp5_ASAP7_75t_L g1539 ( .A1(n_1522), .A2(n_1458), .B1(n_1457), .B2(n_1257), .Y(n_1539) );
NOR2xp33_ASAP7_75t_R g1540 ( .A(n_1529), .B(n_1293), .Y(n_1540) );
NAND4xp25_ASAP7_75t_SL g1541 ( .A(n_1526), .B(n_1375), .C(n_1401), .D(n_1402), .Y(n_1541) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1525), .Y(n_1542) );
OAI221xp5_ASAP7_75t_L g1543 ( .A1(n_1533), .A2(n_1524), .B1(n_1523), .B2(n_1532), .C(n_1530), .Y(n_1543) );
NOR2xp33_ASAP7_75t_L g1544 ( .A(n_1537), .B(n_1315), .Y(n_1544) );
NAND5xp2_ASAP7_75t_L g1545 ( .A(n_1533), .B(n_1132), .C(n_1231), .D(n_1332), .E(n_1334), .Y(n_1545) );
NOR3xp33_ASAP7_75t_SL g1546 ( .A(n_1534), .B(n_1284), .C(n_1385), .Y(n_1546) );
AOI221xp5_ASAP7_75t_SL g1547 ( .A1(n_1539), .A2(n_1412), .B1(n_1409), .B2(n_1408), .C(n_1334), .Y(n_1547) );
NAND4xp25_ASAP7_75t_L g1548 ( .A(n_1535), .B(n_1293), .C(n_1320), .D(n_1319), .Y(n_1548) );
NAND4xp25_ASAP7_75t_SL g1549 ( .A(n_1536), .B(n_1408), .C(n_1400), .D(n_1392), .Y(n_1549) );
AND2x4_ASAP7_75t_L g1550 ( .A(n_1544), .B(n_1542), .Y(n_1550) );
AND2x4_ASAP7_75t_L g1551 ( .A(n_1546), .B(n_1538), .Y(n_1551) );
NOR4xp25_ASAP7_75t_L g1552 ( .A(n_1543), .B(n_1541), .C(n_1540), .D(n_1284), .Y(n_1552) );
INVx4_ASAP7_75t_L g1553 ( .A(n_1548), .Y(n_1553) );
AOI211x1_ASAP7_75t_L g1554 ( .A1(n_1549), .A2(n_1409), .B(n_1412), .C(n_1398), .Y(n_1554) );
INVx2_ASAP7_75t_SL g1555 ( .A(n_1553), .Y(n_1555) );
AO22x2_ASAP7_75t_L g1556 ( .A1(n_1554), .A2(n_1547), .B1(n_1545), .B2(n_1318), .Y(n_1556) );
HB1xp67_ASAP7_75t_L g1557 ( .A(n_1550), .Y(n_1557) );
OAI211xp5_ASAP7_75t_L g1558 ( .A1(n_1552), .A2(n_1318), .B(n_1232), .C(n_1201), .Y(n_1558) );
AND2x2_ASAP7_75t_SL g1559 ( .A(n_1557), .B(n_1551), .Y(n_1559) );
INVx2_ASAP7_75t_SL g1560 ( .A(n_1555), .Y(n_1560) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1558), .Y(n_1561) );
INVx4_ASAP7_75t_L g1562 ( .A(n_1560), .Y(n_1562) );
OAI31xp33_ASAP7_75t_L g1563 ( .A1(n_1561), .A2(n_1556), .A3(n_1383), .B(n_1320), .Y(n_1563) );
XNOR2xp5_ASAP7_75t_L g1564 ( .A(n_1559), .B(n_1556), .Y(n_1564) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1562), .Y(n_1565) );
OAI21xp5_ASAP7_75t_SL g1566 ( .A1(n_1565), .A2(n_1564), .B(n_1563), .Y(n_1566) );
OR2x6_ASAP7_75t_L g1567 ( .A(n_1566), .B(n_1214), .Y(n_1567) );
AOI22xp33_ASAP7_75t_L g1568 ( .A1(n_1567), .A2(n_1430), .B1(n_1429), .B2(n_1427), .Y(n_1568) );
endmodule