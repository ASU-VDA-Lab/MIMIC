module fake_netlist_1_1788_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
NAND2xp5_ASAP7_75t_L g5 ( .A(n_1), .B(n_2), .Y(n_5) );
BUFx6f_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
HB1xp67_ASAP7_75t_L g7 ( .A(n_3), .Y(n_7) );
AO21x1_ASAP7_75t_L g8 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_9), .B(n_3), .Y(n_11) );
INVx2_ASAP7_75t_SL g12 ( .A(n_9), .Y(n_12) );
AOI222xp33_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_10), .B1(n_4), .B2(n_6), .C1(n_8), .C2(n_1), .Y(n_13) );
AOI21xp5_ASAP7_75t_SL g14 ( .A1(n_11), .A2(n_6), .B(n_0), .Y(n_14) );
NOR2xp33_ASAP7_75t_R g15 ( .A(n_13), .B(n_0), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_14), .B(n_0), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
AOI22xp33_ASAP7_75t_SL g18 ( .A1(n_17), .A2(n_15), .B1(n_6), .B2(n_2), .Y(n_18) );
endmodule