module fake_jpeg_15127_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_41),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_36),
.Y(n_60)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_22),
.B1(n_32),
.B2(n_30),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_55),
.B1(n_56),
.B2(n_67),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_32),
.B1(n_22),
.B2(n_21),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_63),
.B(n_28),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_22),
.B1(n_32),
.B2(n_30),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_22),
.B1(n_30),
.B2(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_65),
.Y(n_90)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_34),
.A2(n_32),
.B1(n_21),
.B2(n_20),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_21),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_20),
.B1(n_28),
.B2(n_19),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_79),
.Y(n_95)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_59),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_23),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_33),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_37),
.C(n_41),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_50),
.B1(n_66),
.B2(n_59),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_89),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_26),
.B1(n_19),
.B2(n_23),
.Y(n_107)
);

OAI32xp33_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_56),
.A3(n_48),
.B1(n_23),
.B2(n_28),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_120),
.B1(n_121),
.B2(n_74),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_102),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_46),
.B1(n_62),
.B2(n_58),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_103),
.A2(n_104),
.B1(n_76),
.B2(n_68),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_50),
.B1(n_39),
.B2(n_44),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_26),
.C(n_41),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_37),
.C(n_52),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_26),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_118),
.Y(n_139)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_69),
.A2(n_18),
.B1(n_24),
.B2(n_31),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_25),
.B(n_24),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_76),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_82),
.B1(n_73),
.B2(n_74),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_19),
.A3(n_18),
.B1(n_31),
.B2(n_25),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_123),
.B(n_25),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_64),
.C(n_52),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_129),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_101),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_37),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_126),
.C(n_132),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_100),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_31),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_133),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_71),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_72),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_140),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_137),
.B(n_142),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_64),
.B(n_37),
.Y(n_137)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_113),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_106),
.B(n_94),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_81),
.B(n_24),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_104),
.B(n_103),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_39),
.Y(n_167)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_108),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_98),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_81),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_147),
.B(n_102),
.Y(n_155)
);

AND2x4_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_37),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_101),
.A2(n_70),
.B1(n_85),
.B2(n_73),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_113),
.B1(n_114),
.B2(n_98),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_143),
.B1(n_146),
.B2(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_159),
.C(n_164),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_175),
.B(n_146),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_138),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_173),
.B1(n_148),
.B2(n_130),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_129),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_109),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_167),
.A2(n_140),
.B1(n_148),
.B2(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_169),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_115),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_116),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_132),
.C(n_139),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_134),
.B1(n_148),
.B2(n_99),
.Y(n_191)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_115),
.B1(n_99),
.B2(n_105),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_124),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_134),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_176),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_162),
.A2(n_137),
.B1(n_122),
.B2(n_149),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_178),
.A2(n_160),
.B1(n_163),
.B2(n_173),
.Y(n_206)
);

OR2x6_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_147),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_169),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_171),
.A2(n_146),
.B1(n_123),
.B2(n_147),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_191),
.B1(n_194),
.B2(n_199),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_147),
.B(n_125),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_183),
.Y(n_207)
);

NOR2x1_ASAP7_75t_R g183 ( 
.A(n_158),
.B(n_147),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_168),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_186),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_158),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_139),
.B1(n_148),
.B2(n_142),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_160),
.B1(n_183),
.B2(n_180),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_64),
.C(n_92),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_197),
.C(n_198),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_64),
.C(n_91),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_26),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_16),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_89),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_201),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_78),
.C(n_16),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_105),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_222),
.Y(n_241)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_211),
.A2(n_0),
.B(n_1),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_151),
.B1(n_194),
.B2(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_151),
.B1(n_161),
.B2(n_167),
.Y(n_213)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_179),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_215),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_174),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_197),
.C(n_196),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_203),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_217),
.B(n_221),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_180),
.A2(n_157),
.B1(n_172),
.B2(n_176),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_220),
.B1(n_223),
.B2(n_227),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_180),
.A2(n_157),
.B1(n_150),
.B2(n_138),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_177),
.B(n_150),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_180),
.A2(n_79),
.B1(n_27),
.B2(n_20),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_224),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_189),
.A2(n_17),
.B1(n_16),
.B2(n_2),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_201),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_177),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_232),
.C(n_233),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_184),
.Y(n_232)
);

AOI21x1_ASAP7_75t_SL g234 ( 
.A1(n_207),
.A2(n_199),
.B(n_182),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_250),
.B(n_211),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_236),
.B(n_239),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_198),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_219),
.C(n_225),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_244),
.C(n_246),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_178),
.C(n_17),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_17),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_205),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_224),
.B1(n_210),
.B2(n_209),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_17),
.C(n_16),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_220),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_15),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_249),
.B(n_227),
.Y(n_262)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_253),
.Y(n_282)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_235),
.B(n_226),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_258),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_257),
.B(n_269),
.Y(n_280)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_250),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_259),
.A2(n_260),
.B(n_264),
.Y(n_276)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_215),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_265),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_271),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_237),
.A2(n_204),
.B1(n_206),
.B2(n_218),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_258),
.B1(n_260),
.B2(n_259),
.Y(n_274)
);

AOI221xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_223),
.B1(n_210),
.B2(n_14),
.C(n_13),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_0),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_244),
.B(n_241),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_14),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_246),
.B(n_241),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_277),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_SL g283 ( 
.A1(n_254),
.A2(n_233),
.B(n_242),
.C(n_232),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_3),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_231),
.C(n_2),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_286),
.C(n_262),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_0),
.C(n_3),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_256),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_287),
.B(n_265),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_284),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_289),
.B(n_291),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_270),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_292),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_273),
.A2(n_252),
.B(n_268),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_296),
.B(n_301),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_270),
.C(n_261),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_297),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_263),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_275),
.Y(n_297)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_300),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_SL g306 ( 
.A1(n_299),
.A2(n_287),
.B(n_277),
.C(n_281),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_271),
.C(n_4),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_295),
.B(n_286),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_302),
.B(n_311),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_282),
.B1(n_274),
.B2(n_272),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_307),
.B1(n_290),
.B2(n_288),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_5),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_293),
.A2(n_283),
.B(n_301),
.Y(n_307)
);

OAI211xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_283),
.B(n_13),
.C(n_12),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_4),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_292),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_308),
.Y(n_314)
);

AOI21xp33_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_315),
.B(n_5),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_291),
.C(n_296),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_318),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_SL g323 ( 
.A1(n_317),
.A2(n_12),
.B(n_6),
.C(n_7),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_303),
.C(n_305),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_306),
.B(n_300),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_320),
.B(n_321),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_13),
.Y(n_320)
);

AO221x1_ASAP7_75t_L g330 ( 
.A1(n_323),
.A2(n_324),
.B1(n_325),
.B2(n_7),
.C(n_8),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_SL g324 ( 
.A1(n_321),
.A2(n_12),
.B(n_6),
.C(n_7),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_313),
.A2(n_5),
.B(n_7),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_326),
.Y(n_329)
);

AOI321xp33_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_314),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_329),
.B(n_330),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_9),
.B(n_10),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_10),
.Y(n_334)
);


endmodule