module fake_jpeg_18447_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_14),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_17),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx2_ASAP7_75t_SL g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_57),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_45),
.B1(n_24),
.B2(n_33),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_61),
.B1(n_73),
.B2(n_36),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_17),
.B1(n_27),
.B2(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_18),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_68),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_24),
.B(n_33),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_41),
.B(n_40),
.C(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_41),
.B1(n_40),
.B2(n_27),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_78),
.A2(n_84),
.B1(n_87),
.B2(n_91),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_81),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_24),
.B1(n_32),
.B2(n_29),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_29),
.B1(n_40),
.B2(n_41),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_106),
.B1(n_111),
.B2(n_44),
.Y(n_130)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_48),
.B1(n_47),
.B2(n_38),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_92),
.A2(n_25),
.B1(n_31),
.B2(n_16),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_68),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_101),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_46),
.B1(n_36),
.B2(n_22),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_21),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_59),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_103),
.A2(n_110),
.B1(n_31),
.B2(n_16),
.Y(n_142)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_68),
.Y(n_106)
);

AO22x1_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_48),
.B1(n_47),
.B2(n_38),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_44),
.B(n_16),
.C(n_31),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_21),
.Y(n_108)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

AOI22x1_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_39),
.B1(n_43),
.B2(n_48),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_47),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_113),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_30),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_55),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_19),
.B1(n_26),
.B2(n_20),
.Y(n_126)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

XNOR2x1_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_89),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_118),
.A2(n_126),
.B(n_151),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_36),
.B1(n_44),
.B2(n_34),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_139),
.B1(n_146),
.B2(n_99),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_30),
.B1(n_19),
.B2(n_26),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_120),
.A2(n_142),
.B1(n_148),
.B2(n_11),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_110),
.B(n_94),
.C(n_106),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_1),
.Y(n_183)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_20),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_95),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_78),
.A2(n_34),
.B1(n_25),
.B2(n_22),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_147),
.B1(n_152),
.B2(n_79),
.Y(n_168)
);

NOR2x1p5_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_23),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_140),
.B(n_1),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_107),
.B1(n_76),
.B2(n_77),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_91),
.A2(n_31),
.B1(n_16),
.B2(n_8),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_103),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_0),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_145),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_82),
.A2(n_107),
.B1(n_114),
.B2(n_83),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_114),
.C(n_96),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_158),
.C(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_155),
.B(n_167),
.Y(n_202)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_161),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_175),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_93),
.C(n_105),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_93),
.C(n_105),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_162),
.A2(n_140),
.B1(n_147),
.B2(n_124),
.Y(n_187)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_166),
.A2(n_168),
.B1(n_170),
.B2(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_173),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_135),
.A2(n_116),
.B1(n_104),
.B2(n_90),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_83),
.B(n_86),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_135),
.A2(n_86),
.B1(n_79),
.B2(n_3),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_12),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_184),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_12),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_176),
.A2(n_183),
.B1(n_141),
.B2(n_3),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_1),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_180),
.Y(n_191)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_182),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_133),
.A2(n_1),
.B(n_2),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_138),
.B(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_197),
.B1(n_201),
.B2(n_168),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_189),
.B(n_193),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_160),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_162),
.A2(n_130),
.B1(n_119),
.B2(n_117),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_134),
.Y(n_199)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_117),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_200),
.B(n_211),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_130),
.B1(n_126),
.B2(n_131),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_130),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_205),
.B(n_161),
.Y(n_228)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_141),
.B(n_127),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_216),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_127),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_212),
.A2(n_175),
.B1(n_182),
.B2(n_171),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_158),
.B(n_131),
.C(n_10),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_4),
.C(n_5),
.Y(n_234)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_165),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_157),
.B(n_2),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_190),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_225),
.B1(n_230),
.B2(n_212),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_227),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_155),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_228),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_224),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_209),
.A2(n_172),
.B1(n_183),
.B2(n_170),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_180),
.B1(n_181),
.B2(n_164),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_209),
.A2(n_178),
.B1(n_180),
.B2(n_169),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_232),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_186),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_187),
.A2(n_156),
.B1(n_10),
.B2(n_9),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_207),
.B(n_8),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_231),
.B(n_204),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_214),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_194),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_239),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_244),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_189),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_191),
.B1(n_216),
.B2(n_193),
.Y(n_252)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_5),
.C(n_6),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_240),
.C(n_241),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_6),
.C(n_7),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_208),
.C(n_213),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_206),
.C(n_190),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_217),
.C(n_196),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_206),
.B(n_191),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_257),
.B1(n_224),
.B2(n_226),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_201),
.Y(n_249)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_259),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_252),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_258),
.Y(n_266)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_218),
.A2(n_204),
.B1(n_194),
.B2(n_198),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_207),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_203),
.C(n_198),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_240),
.C(n_241),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_247),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_203),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_261),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_267),
.A2(n_279),
.B1(n_263),
.B2(n_257),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_253),
.C(n_265),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_262),
.A2(n_223),
.B(n_225),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_246),
.B(n_219),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_242),
.Y(n_270)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_255),
.B(n_244),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_277),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_273),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_210),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_276),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_248),
.B(n_238),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_255),
.B(n_221),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_245),
.A2(n_230),
.B1(n_232),
.B2(n_236),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_283),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_234),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_268),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_262),
.B1(n_249),
.B2(n_263),
.Y(n_287)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_269),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_278),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_298),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_246),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_297),
.B(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g299 ( 
.A(n_297),
.B(n_277),
.CI(n_283),
.CON(n_299),
.SN(n_299)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_303),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_304),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_298),
.A2(n_296),
.B1(n_292),
.B2(n_281),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_306),
.A2(n_293),
.B1(n_307),
.B2(n_291),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_266),
.C(n_253),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_289),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_312),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_305),
.A2(n_294),
.B(n_291),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_289),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_288),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

O2A1O1Ixp33_ASAP7_75t_SL g318 ( 
.A1(n_314),
.A2(n_301),
.B(n_290),
.C(n_267),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_315),
.B(n_285),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_279),
.B1(n_215),
.B2(n_266),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_322),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_302),
.C(n_299),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_288),
.C(n_311),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_323),
.B(n_321),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_325),
.Y(n_327)
);

AOI21x1_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_317),
.B(n_323),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_324),
.B(n_314),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_312),
.B(n_318),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_303),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_192),
.Y(n_333)
);


endmodule