module fake_jpeg_15016_n_42 (n_3, n_2, n_1, n_0, n_4, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

OR2x2_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

AOI21xp33_ASAP7_75t_L g12 ( 
.A1(n_0),
.A2(n_5),
.B(n_1),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_12),
.A2(n_1),
.B(n_2),
.Y(n_16)
);

OAI22x1_ASAP7_75t_L g29 ( 
.A1(n_16),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_3),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_6),
.A2(n_3),
.B(n_10),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_10),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_25),
.B1(n_13),
.B2(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_11),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_29),
.C(n_27),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_30),
.B1(n_29),
.B2(n_17),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_37),
.B1(n_23),
.B2(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_16),
.B(n_28),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_39),
.B(n_22),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_22),
.B(n_26),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_15),
.C(n_13),
.Y(n_42)
);


endmodule