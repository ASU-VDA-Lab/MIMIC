module fake_jpeg_2856_n_226 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_226);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_13),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_30),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_2),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_8),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_0),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_67),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_100),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_70),
.B1(n_58),
.B2(n_76),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_74),
.B1(n_69),
.B2(n_72),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_57),
.B1(n_56),
.B2(n_79),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_56),
.B1(n_57),
.B2(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_63),
.Y(n_114)
);

BUFx4f_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_76),
.B1(n_65),
.B2(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_74),
.B1(n_55),
.B2(n_77),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_103),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_57),
.B1(n_62),
.B2(n_79),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_116),
.Y(n_142)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_65),
.B1(n_73),
.B2(n_58),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_83),
.B1(n_55),
.B2(n_59),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_110),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_62),
.B1(n_64),
.B2(n_75),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_113),
.B1(n_118),
.B2(n_96),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_71),
.B1(n_66),
.B2(n_59),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_78),
.B1(n_68),
.B2(n_4),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_0),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_121),
.B(n_31),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_95),
.C(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_28),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_92),
.B(n_99),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_134),
.B(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_78),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_1),
.B(n_4),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_9),
.B(n_10),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_1),
.B(n_5),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_137),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_146),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g145 ( 
.A(n_138),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_16),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_26),
.B1(n_50),
.B2(n_49),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_149),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_12),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_154),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_15),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_159),
.Y(n_174)
);

HB1xp67_ASAP7_75t_SL g158 ( 
.A(n_122),
.Y(n_158)
);

AOI32xp33_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_142),
.A3(n_40),
.B1(n_36),
.B2(n_33),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_25),
.B1(n_48),
.B2(n_47),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_24),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_163),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_23),
.B1(n_45),
.B2(n_43),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_15),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_52),
.B1(n_42),
.B2(n_41),
.Y(n_165)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_179),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_157),
.A2(n_124),
.B1(n_142),
.B2(n_126),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_160),
.Y(n_190)
);

XNOR2x1_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_125),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_157),
.B(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_143),
.Y(n_179)
);

OA21x2_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_183),
.B(n_18),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_16),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_147),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_17),
.B(n_18),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_165),
.B(n_149),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_164),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_190),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_188),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_153),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_181),
.C(n_184),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_192),
.A2(n_194),
.B1(n_184),
.B2(n_185),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_166),
.B(n_150),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_206),
.B1(n_207),
.B2(n_191),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_201),
.B(n_167),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_193),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_205),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_166),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_191),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_187),
.C(n_175),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_209),
.C(n_213),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_198),
.A2(n_171),
.B1(n_169),
.B2(n_168),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_174),
.C(n_171),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_212),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_218),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_214),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_216),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_199),
.B(n_211),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

AOI21x1_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_204),
.B(n_199),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_204),
.A3(n_205),
.B1(n_169),
.B2(n_150),
.C1(n_22),
.C2(n_21),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_19),
.C(n_20),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_19),
.Y(n_226)
);


endmodule