module fake_ariane_2463_n_577 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_117, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_577);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_117;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_577;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_332;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_133;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_424;
wire n_528;
wire n_387;
wire n_406;
wire n_139;
wire n_524;
wire n_130;
wire n_349;
wire n_391;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_330;
wire n_400;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_136;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_565;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_448;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_475;
wire n_135;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_125;
wire n_407;
wire n_254;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_540;
wire n_216;
wire n_544;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_304;
wire n_509;
wire n_306;
wire n_313;
wire n_430;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_337;
wire n_437;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_494;
wire n_131;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_408;
wire n_322;
wire n_251;
wire n_506;
wire n_558;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_573;
wire n_127;
wire n_531;

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_87),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_45),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_12),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_46),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_17),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_40),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_39),
.Y(n_141)
);

BUFx2_ASAP7_75t_SL g142 ( 
.A(n_57),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_26),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_31),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_77),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_50),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_25),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_34),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_58),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_96),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_27),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_79),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_80),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_33),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_54),
.Y(n_157)
);

BUFx10_ASAP7_75t_L g158 ( 
.A(n_16),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_86),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_32),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_65),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_44),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_94),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_8),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_42),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_99),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_124),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_10),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

BUFx2_ASAP7_75t_SL g171 ( 
.A(n_121),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_0),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_10),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_108),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_101),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_73),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_24),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_82),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_76),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_1),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_29),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_129),
.B(n_0),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_127),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_132),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_182),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_136),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_138),
.B(n_1),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_154),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_166),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_134),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_2),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_142),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_150),
.Y(n_208)
);

NOR2xp67_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_2),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_3),
.Y(n_210)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_149),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_3),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_148),
.B(n_4),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

NOR2xp67_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_4),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_125),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_L g223 ( 
.A(n_149),
.B(n_5),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_128),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_135),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_137),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_139),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_149),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_207),
.B(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_140),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_141),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_216),
.B(n_183),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_178),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_224),
.B(n_143),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_218),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_187),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_195),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_186),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_144),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_195),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_199),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_212),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_194),
.Y(n_262)
);

AND2x4_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_178),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

AND2x4_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_203),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_226),
.B(n_146),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_223),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_189),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g270 ( 
.A1(n_226),
.A2(n_160),
.B(n_178),
.Y(n_270)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_227),
.B(n_151),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_200),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_256),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_201),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_273),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_242),
.Y(n_278)
);

AO22x2_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_152),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

BUFx4f_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_153),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_242),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_263),
.Y(n_286)
);

AND2x6_ASAP7_75t_L g287 ( 
.A(n_230),
.B(n_160),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_8),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_251),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_253),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_269),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_243),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_269),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_228),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_232),
.B(n_9),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

AND2x6_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_160),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_228),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_243),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_253),
.B(n_155),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_273),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_156),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_271),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_265),
.B(n_159),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_254),
.A2(n_180),
.B1(n_179),
.B2(n_177),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_257),
.B(n_163),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_272),
.B(n_164),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_229),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_262),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_258),
.B(n_167),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_262),
.B(n_168),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_266),
.A2(n_232),
.B1(n_240),
.B2(n_261),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_233),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_238),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_241),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_244),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_260),
.B(n_9),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_248),
.B(n_174),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_259),
.B(n_175),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_266),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_255),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_259),
.B(n_20),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_247),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_255),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_252),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_249),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

AO22x2_ASAP7_75t_L g333 ( 
.A1(n_296),
.A2(n_268),
.B1(n_236),
.B2(n_237),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_286),
.B(n_231),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_318),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_319),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_234),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_328),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_237),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_290),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_330),
.Y(n_344)
);

AO22x2_ASAP7_75t_L g345 ( 
.A1(n_296),
.A2(n_289),
.B1(n_276),
.B2(n_295),
.Y(n_345)
);

AO22x2_ASAP7_75t_L g346 ( 
.A1(n_289),
.A2(n_236),
.B1(n_235),
.B2(n_270),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_292),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_28),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_278),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_294),
.B(n_30),
.Y(n_351)
);

AO22x2_ASAP7_75t_L g352 ( 
.A1(n_276),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_278),
.Y(n_354)
);

NAND2x1p5_ASAP7_75t_L g355 ( 
.A(n_282),
.B(n_38),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_278),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_285),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_283),
.B(n_280),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_331),
.Y(n_359)
);

OR2x6_ASAP7_75t_L g360 ( 
.A(n_306),
.B(n_41),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_275),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_275),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_281),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_285),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_298),
.B(n_123),
.Y(n_368)
);

NAND2x1p5_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_43),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_298),
.B(n_122),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_291),
.B(n_47),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_298),
.B(n_117),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_297),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_309),
.B(n_115),
.Y(n_374)
);

NAND2x1p5_ASAP7_75t_L g375 ( 
.A(n_317),
.B(n_48),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_287),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_293),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_314),
.B(n_274),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_322),
.Y(n_379)
);

AO22x2_ASAP7_75t_L g380 ( 
.A1(n_279),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_324),
.B(n_114),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_284),
.B(n_59),
.Y(n_382)
);

OR2x6_ASAP7_75t_L g383 ( 
.A(n_279),
.B(n_60),
.Y(n_383)
);

AO22x2_ASAP7_75t_L g384 ( 
.A1(n_307),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_293),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_304),
.B(n_113),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_293),
.Y(n_387)
);

AO21x1_ASAP7_75t_L g388 ( 
.A1(n_326),
.A2(n_327),
.B(n_325),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_277),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_351),
.B(n_288),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_347),
.B(n_303),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_288),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_345),
.B(n_311),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_351),
.B(n_302),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_287),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_349),
.B(n_382),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_338),
.B(n_323),
.Y(n_397)
);

NAND2xp33_ASAP7_75t_SL g398 ( 
.A(n_386),
.B(n_315),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_371),
.B(n_308),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_371),
.B(n_301),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_287),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_359),
.B(n_301),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_361),
.B(n_329),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_341),
.B(n_335),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_336),
.B(n_287),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_337),
.B(n_64),
.Y(n_406)
);

NAND2xp33_ASAP7_75t_SL g407 ( 
.A(n_339),
.B(n_67),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_388),
.B(n_68),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_385),
.B(n_344),
.Y(n_409)
);

NAND2xp33_ASAP7_75t_SL g410 ( 
.A(n_374),
.B(n_69),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_SL g411 ( 
.A(n_342),
.B(n_363),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_334),
.B(n_362),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_333),
.B(n_71),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_333),
.B(n_72),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_364),
.B(n_350),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_354),
.B(n_74),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_356),
.B(n_75),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_357),
.B(n_78),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_366),
.B(n_83),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_367),
.B(n_84),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_377),
.B(n_387),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_381),
.B(n_85),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_408),
.A2(n_368),
.B(n_370),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_389),
.B(n_360),
.Y(n_424)
);

AO31x2_ASAP7_75t_L g425 ( 
.A1(n_413),
.A2(n_372),
.A3(n_373),
.B(n_365),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_401),
.B(n_355),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_401),
.B(n_353),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_395),
.A2(n_348),
.B(n_332),
.Y(n_429)
);

O2A1O1Ixp5_ASAP7_75t_L g430 ( 
.A1(n_398),
.A2(n_332),
.B(n_340),
.C(n_343),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g431 ( 
.A1(n_422),
.A2(n_369),
.B(n_375),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_397),
.B(n_345),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_396),
.A2(n_346),
.B(n_352),
.Y(n_433)
);

AOI221x1_ASAP7_75t_L g434 ( 
.A1(n_414),
.A2(n_352),
.B1(n_384),
.B2(n_380),
.C(n_346),
.Y(n_434)
);

AO31x2_ASAP7_75t_L g435 ( 
.A1(n_404),
.A2(n_384),
.A3(n_380),
.B(n_383),
.Y(n_435)
);

AOI21xp33_ASAP7_75t_L g436 ( 
.A1(n_399),
.A2(n_383),
.B(n_376),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_412),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_393),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_392),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g440 ( 
.A1(n_422),
.A2(n_88),
.B(n_89),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_403),
.A2(n_90),
.B(n_91),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_394),
.B(n_93),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_415),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_391),
.Y(n_444)
);

OAI21x1_ASAP7_75t_L g445 ( 
.A1(n_405),
.A2(n_95),
.B(n_97),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_400),
.A2(n_102),
.B(n_103),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_410),
.A2(n_107),
.B(n_407),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_402),
.A2(n_421),
.B(n_406),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_411),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_436),
.A2(n_433),
.B1(n_438),
.B2(n_434),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_438),
.A2(n_390),
.B1(n_416),
.B2(n_417),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_423),
.A2(n_418),
.B(n_419),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_427),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_420),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_437),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_439),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g458 ( 
.A1(n_431),
.A2(n_447),
.B(n_445),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_443),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_424),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_426),
.Y(n_461)
);

AOI21x1_ASAP7_75t_L g462 ( 
.A1(n_432),
.A2(n_441),
.B(n_442),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_435),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_430),
.Y(n_464)
);

BUFx2_ASAP7_75t_SL g465 ( 
.A(n_449),
.Y(n_465)
);

O2A1O1Ixp5_ASAP7_75t_SL g466 ( 
.A1(n_448),
.A2(n_435),
.B(n_425),
.C(n_440),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_435),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_446),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_425),
.B(n_389),
.Y(n_469)
);

OA21x2_ASAP7_75t_L g470 ( 
.A1(n_425),
.A2(n_429),
.B(n_433),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_436),
.A2(n_383),
.B1(n_380),
.B2(n_352),
.Y(n_471)
);

OA21x2_ASAP7_75t_L g472 ( 
.A1(n_429),
.A2(n_433),
.B(n_434),
.Y(n_472)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_423),
.A2(n_431),
.B(n_408),
.Y(n_473)
);

NAND2x1p5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_467),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_459),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_469),
.B(n_463),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_455),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_459),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_453),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_470),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_470),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_471),
.A2(n_450),
.B1(n_472),
.B2(n_461),
.Y(n_482)
);

AO21x2_ASAP7_75t_L g483 ( 
.A1(n_464),
.A2(n_473),
.B(n_462),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_461),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_460),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_468),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_457),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_465),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_468),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_452),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_452),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_458),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_468),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_461),
.B(n_456),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_450),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_461),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_456),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_451),
.A2(n_466),
.B(n_454),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_456),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_456),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_R g501 ( 
.A(n_494),
.B(n_488),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_451),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_468),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_484),
.B(n_478),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_498),
.B(n_487),
.Y(n_505)
);

OR2x6_ASAP7_75t_L g506 ( 
.A(n_484),
.B(n_496),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_497),
.B(n_475),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_475),
.B(n_496),
.Y(n_508)
);

OR2x4_ASAP7_75t_L g509 ( 
.A(n_476),
.B(n_481),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_479),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_478),
.B(n_476),
.Y(n_511)
);

BUFx8_ASAP7_75t_SL g512 ( 
.A(n_486),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_482),
.B(n_474),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_486),
.B(n_493),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_495),
.B(n_474),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_R g516 ( 
.A(n_486),
.B(n_489),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_495),
.B(n_481),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_R g518 ( 
.A(n_489),
.B(n_493),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_510),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_507),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_516),
.B(n_493),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_508),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_503),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_480),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_505),
.B(n_480),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_511),
.B(n_489),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_499),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_504),
.B(n_514),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_515),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_506),
.B(n_474),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_502),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_L g532 ( 
.A(n_525),
.B(n_518),
.C(n_501),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_483),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_526),
.B(n_513),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_525),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_519),
.Y(n_536)
);

NAND2x1p5_ASAP7_75t_L g537 ( 
.A(n_521),
.B(n_512),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_520),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_535),
.B(n_527),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_538),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_531),
.B(n_530),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_538),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_537),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_534),
.B(n_523),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_533),
.B(n_524),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_539),
.B(n_536),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_SL g547 ( 
.A(n_543),
.B(n_521),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_540),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_544),
.B(n_532),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_539),
.B(n_524),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_549),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_548),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_546),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_547),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_550),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_551),
.B(n_553),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_552),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_552),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_556),
.B(n_555),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_557),
.B(n_554),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_559),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_561),
.B(n_558),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_562),
.Y(n_563)
);

NAND4xp75_ASAP7_75t_L g564 ( 
.A(n_563),
.B(n_560),
.C(n_554),
.D(n_544),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_R g565 ( 
.A(n_564),
.B(n_542),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_565),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_566),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_567),
.Y(n_568)
);

AOI31xp33_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_545),
.A3(n_541),
.B(n_513),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_483),
.B1(n_522),
.B2(n_509),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_569),
.B(n_483),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_571),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_570),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_572),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_573),
.Y(n_575)
);

AOI221xp5_ASAP7_75t_L g576 ( 
.A1(n_574),
.A2(n_492),
.B1(n_491),
.B2(n_490),
.C(n_500),
.Y(n_576)
);

OA22x2_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_575),
.B1(n_492),
.B2(n_500),
.Y(n_577)
);


endmodule