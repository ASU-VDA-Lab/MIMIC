module fake_jpeg_16368_n_377 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_377);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_377;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_5),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_41),
.B(n_62),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_42),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_46),
.Y(n_67)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_48),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_51),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_57),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx5_ASAP7_75t_SL g102 ( 
.A(n_56),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_21),
.B1(n_23),
.B2(n_37),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_77),
.A2(n_88),
.B1(n_90),
.B2(n_93),
.Y(n_133)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_40),
.A2(n_18),
.B1(n_15),
.B2(n_35),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_85),
.B1(n_108),
.B2(n_33),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_44),
.A2(n_54),
.B1(n_59),
.B2(n_66),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_60),
.A2(n_37),
.B1(n_36),
.B2(n_18),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_41),
.A2(n_37),
.B1(n_29),
.B2(n_22),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_43),
.A2(n_35),
.B1(n_15),
.B2(n_19),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_41),
.B(n_22),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_101),
.Y(n_122)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

BUFx2_ASAP7_75t_SL g118 ( 
.A(n_99),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_46),
.B(n_62),
.Y(n_101)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_51),
.A2(n_29),
.B1(n_19),
.B2(n_16),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_110),
.B1(n_111),
.B2(n_26),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_53),
.A2(n_33),
.B1(n_31),
.B2(n_26),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_57),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_48),
.A2(n_16),
.B1(n_33),
.B2(n_31),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_55),
.A2(n_16),
.B1(n_33),
.B2(n_31),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_42),
.B(n_16),
.C(n_26),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_7),
.Y(n_124)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_117),
.B(n_137),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_119),
.A2(n_135),
.B1(n_152),
.B2(n_157),
.Y(n_168)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_125),
.Y(n_185)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_27),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_126),
.B(n_146),
.Y(n_191)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_71),
.B(n_70),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_134),
.A2(n_145),
.B(n_123),
.Y(n_206)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_136),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_104),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_7),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_83),
.Y(n_139)
);

INVx3_ASAP7_75t_SL g203 ( 
.A(n_139),
.Y(n_203)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_142),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_6),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_80),
.B(n_6),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_68),
.B(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_147),
.B(n_160),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_111),
.A2(n_50),
.B(n_27),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_0),
.C(n_162),
.Y(n_186)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_86),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_77),
.B(n_5),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_155),
.Y(n_183)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_112),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_157)
);

BUFx8_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_79),
.Y(n_159)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_68),
.B(n_25),
.Y(n_160)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_106),
.A2(n_5),
.B(n_2),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_161),
.A2(n_123),
.B(n_142),
.C(n_149),
.Y(n_209)
);

AND2x4_ASAP7_75t_L g162 ( 
.A(n_108),
.B(n_0),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_161),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_116),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_13),
.B1(n_6),
.B2(n_8),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_79),
.B(n_4),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_125),
.A2(n_116),
.B1(n_102),
.B2(n_69),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_167),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_153),
.A2(n_85),
.B1(n_78),
.B2(n_113),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_171),
.A2(n_177),
.B1(n_182),
.B2(n_187),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_162),
.A2(n_84),
.B1(n_98),
.B2(n_13),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_138),
.A2(n_81),
.B1(n_97),
.B2(n_84),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_119),
.A2(n_97),
.B1(n_98),
.B2(n_13),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_0),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_196),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_162),
.A2(n_0),
.B1(n_10),
.B2(n_133),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_127),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_124),
.A2(n_0),
.B1(n_134),
.B2(n_148),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_118),
.Y(n_188)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_150),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_124),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_190),
.A2(n_193),
.B(n_205),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_122),
.B(n_143),
.CI(n_164),
.CON(n_192),
.SN(n_192)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_192),
.B(n_178),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_117),
.A2(n_128),
.B1(n_130),
.B2(n_156),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_195),
.A2(n_205),
.B1(n_189),
.B2(n_188),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_136),
.B(n_144),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_131),
.B(n_140),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_202),
.C(n_206),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_141),
.Y(n_201)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_141),
.C(n_129),
.Y(n_202)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_158),
.A2(n_151),
.A3(n_145),
.B1(n_132),
.B2(n_139),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_204),
.B(n_206),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_128),
.B(n_130),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_204),
.B(n_178),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_159),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_127),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_212),
.A2(n_220),
.B(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_198),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_222),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_127),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_219),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_199),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_186),
.Y(n_220)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_175),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_224),
.A2(n_248),
.B(n_250),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_190),
.A2(n_188),
.B1(n_184),
.B2(n_168),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_225),
.A2(n_229),
.B1(n_233),
.B2(n_235),
.Y(n_254)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_205),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_183),
.B(n_176),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_230),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_209),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_175),
.B(n_192),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_238),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_198),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_207),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_185),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_245),
.C(n_249),
.Y(n_251)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_193),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_172),
.Y(n_239)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_185),
.B(n_193),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_246),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_243),
.B1(n_221),
.B2(n_229),
.Y(n_266)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_189),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_242),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_190),
.A2(n_182),
.B1(n_170),
.B2(n_177),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_244),
.A2(n_214),
.B1(n_222),
.B2(n_215),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_197),
.C(n_190),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_194),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_203),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_174),
.B(n_191),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_264),
.C(n_275),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_208),
.B1(n_169),
.B2(n_166),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_255),
.A2(n_269),
.B1(n_274),
.B2(n_254),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_232),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_257),
.B(n_251),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_212),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_270),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_203),
.C(n_208),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_258),
.B1(n_260),
.B2(n_252),
.Y(n_288)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_221),
.A2(n_180),
.B1(n_243),
.B2(n_248),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_224),
.B(n_180),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_238),
.A2(n_240),
.B1(n_216),
.B2(n_223),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_271),
.A2(n_278),
.B1(n_277),
.B2(n_262),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_219),
.B(n_218),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_220),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_220),
.A2(n_212),
.B(n_216),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_227),
.B(n_211),
.C(n_249),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_257),
.C(n_281),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_241),
.A2(n_211),
.B1(n_227),
.B2(n_213),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g280 ( 
.A(n_214),
.B(n_234),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_281),
.A2(n_283),
.B(n_267),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_247),
.A2(n_240),
.B(n_238),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_226),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_290),
.C(n_301),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_287),
.A2(n_288),
.B1(n_298),
.B2(n_285),
.Y(n_322)
);

NOR3xp33_ASAP7_75t_SL g289 ( 
.A(n_265),
.B(n_276),
.C(n_271),
.Y(n_289)
);

NAND3xp33_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_308),
.C(n_302),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_253),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_282),
.B(n_279),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_299),
.Y(n_316)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_252),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_296),
.A2(n_305),
.B(n_307),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_300),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_270),
.A2(n_260),
.B1(n_264),
.B2(n_262),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_263),
.Y(n_299)
);

AO21x2_ASAP7_75t_SL g302 ( 
.A1(n_283),
.A2(n_278),
.B(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_256),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_304),
.Y(n_324)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_282),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_273),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_306),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_280),
.A2(n_255),
.B(n_259),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_261),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_261),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_286),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_265),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_302),
.B(n_296),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_302),
.A2(n_288),
.B1(n_295),
.B2(n_298),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_312),
.A2(n_318),
.B1(n_329),
.B2(n_324),
.Y(n_340)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_314),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_290),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_317),
.B(n_323),
.C(n_327),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_310),
.A2(n_296),
.B1(n_304),
.B2(n_303),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_318),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_322),
.A2(n_320),
.B1(n_312),
.B2(n_313),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_291),
.B(n_297),
.Y(n_323)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_325),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_301),
.C(n_300),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_292),
.B(n_291),
.C(n_290),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_315),
.B(n_319),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_335),
.C(n_339),
.Y(n_351)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_333),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_330),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_316),
.Y(n_336)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_319),
.A2(n_320),
.B(n_321),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_338),
.B(n_340),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_323),
.B(n_327),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_311),
.A2(n_320),
.B1(n_318),
.B2(n_315),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_338),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_311),
.B(n_328),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_342),
.C(n_339),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_326),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_345),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_328),
.A2(n_254),
.B1(n_225),
.B2(n_316),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_346),
.B(n_332),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_340),
.B(n_337),
.Y(n_350)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_350),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_353),
.B(n_342),
.C(n_335),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_331),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_354),
.B(n_331),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_336),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_355),
.B(n_349),
.Y(n_359)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_356),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_351),
.B(n_343),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_358),
.C(n_362),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_334),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_359),
.B(n_361),
.C(n_347),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_360),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_349),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_366),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_367),
.B(n_354),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_363),
.A2(n_346),
.B(n_352),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_369),
.B(n_365),
.C(n_361),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_370),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_372),
.B(n_368),
.Y(n_373)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_373),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_371),
.C(n_353),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_375),
.B(n_351),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_357),
.Y(n_377)
);


endmodule