module fake_ariane_4_n_168 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_16, n_5, n_12, n_15, n_10, n_168);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_168;

wire n_83;
wire n_56;
wire n_60;
wire n_160;
wire n_64;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_34;
wire n_158;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_19;
wire n_40;
wire n_152;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_21;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_24;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_121;
wire n_93;
wire n_118;
wire n_23;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_28;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;
wire n_25;

INVxp33_ASAP7_75t_SL g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVxp33_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

AND2x4_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_19),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

AO22x2_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_30),
.B1(n_32),
.B2(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2x1p5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_27),
.B1(n_4),
.B2(n_5),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_17),
.Y(n_63)
);

AO22x2_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_64)
);

AO22x2_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_8),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_11),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2x1p5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_37),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_42),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_42),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_42),
.B1(n_48),
.B2(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2x1p5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_57),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_62),
.B(n_60),
.Y(n_86)
);

NOR2xp67_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_39),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_57),
.B(n_45),
.C(n_49),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_53),
.Y(n_94)
);

CKINVDCx6p67_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

OAI211xp5_ASAP7_75t_SL g97 ( 
.A1(n_91),
.A2(n_81),
.B(n_79),
.C(n_52),
.Y(n_97)
);

OAI21x1_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_82),
.B(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_76),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_81),
.B(n_74),
.Y(n_101)
);

OAI211xp5_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_79),
.B(n_51),
.C(n_80),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

NOR2x1_ASAP7_75t_SL g104 ( 
.A(n_85),
.B(n_82),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_77),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_77),
.B1(n_53),
.B2(n_64),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_71),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_53),
.Y(n_108)
);

AOI221xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_64),
.B1(n_65),
.B2(n_71),
.C(n_80),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_82),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_85),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_80),
.B(n_64),
.C(n_65),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_111),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_88),
.C(n_86),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_107),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_92),
.B(n_90),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_64),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_94),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

AOI31xp33_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_106),
.A3(n_109),
.B(n_108),
.Y(n_131)
);

NOR3xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_102),
.C(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_65),
.B1(n_107),
.B2(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_118),
.B(n_127),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_117),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_65),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_136),
.B(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_142),
.Y(n_150)
);

OAI222xp33_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_126),
.B1(n_135),
.B2(n_131),
.C1(n_133),
.C2(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

AOI221xp5_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_140),
.B1(n_141),
.B2(n_147),
.C(n_113),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_134),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_138),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_145),
.Y(n_156)
);

NAND3x2_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_152),
.C(n_149),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

NAND4xp75_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_152),
.C(n_151),
.D(n_110),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_155),
.B(n_98),
.Y(n_160)
);

OAI221xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_159),
.B1(n_157),
.B2(n_87),
.C(n_138),
.Y(n_161)
);

OAI211xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_11),
.B(n_125),
.C(n_87),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_128),
.B1(n_104),
.B2(n_110),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_162),
.A2(n_104),
.B1(n_122),
.B2(n_124),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_124),
.Y(n_166)
);

FAx1_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_164),
.CI(n_125),
.CON(n_167),
.SN(n_167)
);

AOI221xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_166),
.B1(n_90),
.B2(n_125),
.C(n_98),
.Y(n_168)
);


endmodule