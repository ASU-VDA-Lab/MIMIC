module fake_aes_7306_n_889 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_177, n_130, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_166, n_162, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_889);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_889;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_227;
wire n_476;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_818;
wire n_844;
wire n_725;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_828;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_357;
wire n_245;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_208;
wire n_200;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_875;
wire n_339;
wire n_657;
wire n_583;
wire n_728;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g182 ( .A(n_23), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_66), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_146), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_106), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_100), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_148), .B(n_82), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
INVx1_ASAP7_75t_SL g190 ( .A(n_44), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_94), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_167), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_5), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_83), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_181), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_46), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_162), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_140), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_33), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_5), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_157), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_110), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_103), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_166), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_61), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g206 ( .A(n_40), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g207 ( .A(n_89), .Y(n_207) );
BUFx10_ASAP7_75t_L g208 ( .A(n_98), .Y(n_208) );
INVxp67_ASAP7_75t_SL g209 ( .A(n_111), .Y(n_209) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_64), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_101), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_33), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_36), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_123), .B(n_172), .Y(n_214) );
INVxp67_ASAP7_75t_SL g215 ( .A(n_168), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_35), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_54), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_155), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_135), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_143), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_104), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_18), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_128), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_43), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_152), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_81), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_70), .Y(n_227) );
BUFx5_ASAP7_75t_L g228 ( .A(n_149), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_74), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_34), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_121), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_139), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_37), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_116), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_107), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_113), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_95), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_47), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_165), .Y(n_239) );
INVx1_ASAP7_75t_SL g240 ( .A(n_31), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_174), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_36), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_180), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_126), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_60), .Y(n_245) );
INVxp33_ASAP7_75t_SL g246 ( .A(n_118), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_96), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_22), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_56), .Y(n_249) );
BUFx10_ASAP7_75t_L g250 ( .A(n_93), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_127), .Y(n_251) );
CKINVDCx16_ASAP7_75t_R g252 ( .A(n_90), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_45), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_55), .Y(n_254) );
INVxp67_ASAP7_75t_SL g255 ( .A(n_147), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_67), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_31), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_71), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_109), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_3), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_108), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_145), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_112), .Y(n_263) );
INVxp67_ASAP7_75t_SL g264 ( .A(n_61), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g265 ( .A(n_57), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_42), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_129), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_178), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_30), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_75), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_153), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_80), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_8), .Y(n_273) );
BUFx10_ASAP7_75t_L g274 ( .A(n_32), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_62), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_97), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_120), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_154), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_82), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_138), .Y(n_280) );
CKINVDCx14_ASAP7_75t_R g281 ( .A(n_12), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_177), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_3), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_105), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_144), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_131), .Y(n_286) );
BUFx3_ASAP7_75t_L g287 ( .A(n_7), .Y(n_287) );
BUFx8_ASAP7_75t_SL g288 ( .A(n_117), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_173), .Y(n_289) );
NOR2x1_ASAP7_75t_L g290 ( .A(n_248), .B(n_0), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_210), .B(n_279), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_228), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_228), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_228), .Y(n_294) );
BUFx8_ASAP7_75t_L g295 ( .A(n_268), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_199), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_288), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_281), .Y(n_298) );
XNOR2xp5_ASAP7_75t_L g299 ( .A(n_254), .B(n_1), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_199), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_186), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_228), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_228), .Y(n_303) );
OA21x2_ASAP7_75t_L g304 ( .A1(n_189), .A2(n_85), .B(n_84), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_186), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_213), .Y(n_306) );
OA21x2_ASAP7_75t_L g307 ( .A1(n_189), .A2(n_87), .B(n_86), .Y(n_307) );
INVx5_ASAP7_75t_L g308 ( .A(n_186), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_248), .B(n_2), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_281), .B(n_2), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_213), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_206), .A2(n_7), .B1(n_4), .B2(n_6), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_287), .B(n_4), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_230), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_217), .Y(n_315) );
BUFx8_ASAP7_75t_SL g316 ( .A(n_254), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_265), .B(n_6), .Y(n_317) );
CKINVDCx8_ASAP7_75t_R g318 ( .A(n_207), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_288), .Y(n_319) );
NOR2x1_ASAP7_75t_L g320 ( .A(n_287), .B(n_8), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_217), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_186), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_274), .Y(n_323) );
AOI22xp5_ASAP7_75t_SL g324 ( .A1(n_260), .A2(n_11), .B1(n_9), .B2(n_10), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_252), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_274), .B(n_10), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_231), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_292), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_292), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_292), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_298), .B(n_246), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_293), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_309), .A2(n_183), .B1(n_193), .B2(n_182), .Y(n_333) );
AND3x2_ASAP7_75t_L g334 ( .A(n_325), .B(n_264), .C(n_215), .Y(n_334) );
INVx4_ASAP7_75t_L g335 ( .A(n_309), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_301), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_313), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_293), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_301), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_304), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_325), .B(n_208), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_301), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_291), .B(n_208), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_293), .B(n_192), .Y(n_344) );
OR2x6_ASAP7_75t_L g345 ( .A(n_312), .B(n_187), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_323), .B(n_246), .Y(n_346) );
OR2x6_ASAP7_75t_L g347 ( .A(n_312), .B(n_227), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_297), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_310), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_294), .B(n_192), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_295), .B(n_250), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_295), .Y(n_352) );
INVx4_ASAP7_75t_L g353 ( .A(n_313), .Y(n_353) );
BUFx2_ASAP7_75t_L g354 ( .A(n_295), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_313), .A2(n_222), .B1(n_233), .B2(n_226), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_296), .A2(n_245), .B1(n_253), .B2(n_238), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_310), .Y(n_357) );
INVx4_ASAP7_75t_L g358 ( .A(n_304), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_319), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_326), .B(n_250), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_305), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_305), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_302), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_361), .B(n_317), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_349), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_357), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_333), .A2(n_318), .B1(n_195), .B2(n_198), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_361), .B(n_295), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_335), .A2(n_303), .B1(n_296), .B2(n_300), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_343), .B(n_349), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_343), .A2(n_195), .B1(n_198), .B2(n_197), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_341), .A2(n_204), .B1(n_219), .B2(n_197), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_341), .B(n_318), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_346), .A2(n_219), .B1(n_235), .B2(n_204), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_340), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_352), .B(n_290), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_331), .B(n_300), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_335), .B(n_306), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_335), .B(n_290), .Y(n_380) );
NOR2xp33_ASAP7_75t_SL g381 ( .A(n_352), .B(n_354), .Y(n_381) );
INVx2_ASAP7_75t_SL g382 ( .A(n_354), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_353), .A2(n_303), .B1(n_315), .B2(n_311), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_337), .A2(n_307), .B(n_304), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_353), .B(n_320), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_345), .A2(n_247), .B1(n_284), .B2(n_235), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_337), .A2(n_303), .B1(n_321), .B2(n_266), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_364), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_328), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_333), .B(n_184), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_351), .B(n_321), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_328), .Y(n_392) );
INVx2_ASAP7_75t_SL g393 ( .A(n_334), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_355), .B(n_185), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_329), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_329), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_330), .B(n_188), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g398 ( .A1(n_345), .A2(n_324), .B1(n_260), .B2(n_283), .Y(n_398) );
INVxp67_ASAP7_75t_L g399 ( .A(n_345), .Y(n_399) );
AND2x4_ASAP7_75t_SL g400 ( .A(n_345), .B(n_314), .Y(n_400) );
NOR3xp33_ASAP7_75t_L g401 ( .A(n_348), .B(n_240), .C(n_190), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_359), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_347), .A2(n_269), .B1(n_270), .B2(n_256), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_340), .A2(n_307), .B(n_304), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g405 ( .A1(n_358), .A2(n_307), .B(n_191), .Y(n_405) );
OAI22xp33_ASAP7_75t_SL g406 ( .A1(n_345), .A2(n_196), .B1(n_205), .B2(n_200), .Y(n_406) );
NAND2x2_ASAP7_75t_L g407 ( .A(n_334), .B(n_316), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_344), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_332), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_338), .Y(n_410) );
NOR2xp67_ASAP7_75t_L g411 ( .A(n_344), .B(n_299), .Y(n_411) );
AND2x2_ASAP7_75t_SL g412 ( .A(n_356), .B(n_307), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_350), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_350), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_345), .Y(n_415) );
INVx1_ASAP7_75t_SL g416 ( .A(n_364), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_347), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_347), .A2(n_284), .B1(n_247), .B2(n_212), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_360), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_340), .B(n_324), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_358), .B(n_194), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_336), .A2(n_275), .B1(n_272), .B2(n_227), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_336), .B(n_299), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_339), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_339), .A2(n_216), .B1(n_229), .B2(n_224), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_342), .Y(n_426) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_376), .Y(n_427) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_376), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_388), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_369), .B(n_283), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_374), .B(n_273), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_404), .A2(n_255), .B(n_209), .Y(n_432) );
NOR2x1_ASAP7_75t_R g433 ( .A(n_420), .B(n_221), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_381), .B(n_236), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_408), .Y(n_435) );
O2A1O1Ixp33_ASAP7_75t_L g436 ( .A1(n_371), .A2(n_249), .B(n_257), .C(n_242), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_414), .Y(n_437) );
INVx4_ASAP7_75t_L g438 ( .A(n_388), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_405), .A2(n_202), .B(n_201), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_366), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_419), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_416), .B(n_251), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_419), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_379), .Y(n_444) );
BUFx8_ASAP7_75t_L g445 ( .A(n_420), .Y(n_445) );
OA22x2_ASAP7_75t_L g446 ( .A1(n_373), .A2(n_220), .B1(n_223), .B2(n_218), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_403), .A2(n_417), .B1(n_415), .B2(n_412), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_380), .A2(n_234), .B(n_232), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_377), .B(n_237), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_400), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_385), .A2(n_243), .B(n_241), .Y(n_451) );
INVx4_ASAP7_75t_L g452 ( .A(n_409), .Y(n_452) );
BUFx3_ASAP7_75t_L g453 ( .A(n_400), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_372), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_411), .B(n_258), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_410), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_410), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_379), .Y(n_458) );
AO22x1_ASAP7_75t_L g459 ( .A1(n_368), .A2(n_214), .B1(n_263), .B2(n_261), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_389), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_391), .B(n_258), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_393), .B(n_276), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_392), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_423), .B(n_277), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_395), .Y(n_465) );
AND2x2_ASAP7_75t_SL g466 ( .A(n_386), .B(n_214), .Y(n_466) );
AOI21xp5_ASAP7_75t_SL g467 ( .A1(n_396), .A2(n_239), .B(n_203), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_418), .A2(n_285), .B1(n_286), .B2(n_282), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_391), .B(n_289), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_387), .A2(n_211), .B1(n_244), .B2(n_225), .Y(n_470) );
OR2x6_ASAP7_75t_SL g471 ( .A(n_398), .B(n_262), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_394), .A2(n_383), .B1(n_370), .B2(n_387), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_425), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_383), .A2(n_278), .B1(n_280), .B2(n_271), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_422), .A2(n_280), .B1(n_278), .B2(n_259), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_397), .A2(n_267), .B1(n_231), .B2(n_305), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_424), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_401), .B(n_13), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_407), .Y(n_479) );
AO21x1_ASAP7_75t_L g480 ( .A1(n_424), .A2(n_363), .B(n_362), .Y(n_480) );
AOI33xp33_ASAP7_75t_L g481 ( .A1(n_407), .A2(n_363), .A3(n_362), .B1(n_15), .B2(n_16), .B3(n_17), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_426), .Y(n_482) );
AO21x1_ASAP7_75t_L g483 ( .A1(n_404), .A2(n_363), .B(n_362), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_413), .B(n_14), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_403), .A2(n_267), .B1(n_308), .B2(n_322), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_413), .B(n_15), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_404), .A2(n_308), .B(n_267), .Y(n_487) );
NAND3xp33_ASAP7_75t_L g488 ( .A(n_378), .B(n_308), .C(n_322), .Y(n_488) );
AO32x1_ASAP7_75t_L g489 ( .A1(n_413), .A2(n_327), .A3(n_322), .B1(n_308), .B2(n_19), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_413), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_420), .A2(n_327), .B1(n_322), .B2(n_18), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_366), .B(n_16), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_404), .A2(n_327), .B(n_88), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_399), .A2(n_327), .B1(n_20), .B2(n_17), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_413), .Y(n_495) );
OR2x6_ASAP7_75t_SL g496 ( .A(n_402), .B(n_20), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_366), .B(n_21), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_399), .A2(n_25), .B1(n_22), .B2(n_24), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_413), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_404), .A2(n_92), .B(n_91), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_413), .B(n_24), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_382), .B(n_26), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_388), .Y(n_503) );
BUFx3_ASAP7_75t_L g504 ( .A(n_402), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_366), .B(n_26), .Y(n_505) );
CKINVDCx6p67_ASAP7_75t_R g506 ( .A(n_366), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_420), .A2(n_29), .B1(n_27), .B2(n_28), .Y(n_507) );
AOI21x1_ASAP7_75t_L g508 ( .A1(n_404), .A2(n_102), .B(n_99), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_413), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_440), .Y(n_510) );
BUFx2_ASAP7_75t_R g511 ( .A(n_471), .Y(n_511) );
AO31x2_ASAP7_75t_L g512 ( .A1(n_483), .A2(n_480), .A3(n_439), .B(n_493), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_435), .Y(n_513) );
AO31x2_ASAP7_75t_L g514 ( .A1(n_500), .A2(n_38), .A3(n_39), .B(n_40), .Y(n_514) );
AO32x2_ASAP7_75t_L g515 ( .A1(n_474), .A2(n_38), .A3(n_39), .B1(n_41), .B2(n_42), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_490), .Y(n_516) );
OR2x6_ASAP7_75t_L g517 ( .A(n_453), .B(n_41), .Y(n_517) );
INVxp67_ASAP7_75t_SL g518 ( .A(n_445), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_495), .Y(n_519) );
AO31x2_ASAP7_75t_L g520 ( .A1(n_470), .A2(n_48), .A3(n_49), .B(n_50), .Y(n_520) );
AOI211x1_ASAP7_75t_L g521 ( .A1(n_459), .A2(n_48), .B(n_49), .C(n_50), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_444), .B(n_51), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_458), .B(n_51), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_454), .A2(n_52), .B1(n_53), .B2(n_54), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_436), .A2(n_56), .B(n_57), .C(n_58), .Y(n_525) );
AO32x2_ASAP7_75t_L g526 ( .A1(n_470), .A2(n_58), .A3(n_59), .B1(n_60), .B2(n_63), .Y(n_526) );
INVx8_ASAP7_75t_L g527 ( .A(n_502), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_427), .Y(n_528) );
OAI21x1_ASAP7_75t_L g529 ( .A1(n_508), .A2(n_115), .B(n_114), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_477), .A2(n_461), .B(n_457), .Y(n_530) );
INVx6_ASAP7_75t_SL g531 ( .A(n_449), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_456), .A2(n_141), .B(n_179), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_460), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_499), .B(n_65), .Y(n_534) );
AO32x2_ASAP7_75t_L g535 ( .A1(n_475), .A2(n_68), .A3(n_69), .B1(n_71), .B2(n_72), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_441), .A2(n_443), .B(n_469), .Y(n_536) );
CKINVDCx11_ASAP7_75t_R g537 ( .A(n_496), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_504), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_509), .B(n_73), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_484), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_472), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_464), .B(n_77), .Y(n_542) );
AND2x4_ASAP7_75t_L g543 ( .A(n_450), .B(n_78), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_438), .B(n_449), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_473), .B(n_79), .Y(n_545) );
OAI21x1_ASAP7_75t_L g546 ( .A1(n_488), .A2(n_142), .B(n_176), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_486), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_431), .B(n_80), .Y(n_548) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_428), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_501), .Y(n_550) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_428), .Y(n_551) );
INVx3_ASAP7_75t_SL g552 ( .A(n_479), .Y(n_552) );
INVxp67_ASAP7_75t_SL g553 ( .A(n_438), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_463), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_466), .B(n_119), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_465), .Y(n_556) );
AO31x2_ASAP7_75t_L g557 ( .A1(n_485), .A2(n_122), .A3(n_124), .B(n_125), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_507), .Y(n_558) );
INVx5_ASAP7_75t_L g559 ( .A(n_428), .Y(n_559) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_448), .A2(n_130), .B(n_132), .C(n_133), .Y(n_560) );
OR2x6_ASAP7_75t_L g561 ( .A(n_446), .B(n_134), .Y(n_561) );
NAND3xp33_ASAP7_75t_L g562 ( .A(n_491), .B(n_136), .C(n_137), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_482), .B(n_156), .Y(n_563) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_451), .A2(n_158), .B(n_159), .C(n_160), .Y(n_564) );
INVx3_ASAP7_75t_SL g565 ( .A(n_455), .Y(n_565) );
BUFx2_ASAP7_75t_L g566 ( .A(n_433), .Y(n_566) );
AO22x2_ASAP7_75t_L g567 ( .A1(n_498), .A2(n_161), .B1(n_163), .B2(n_164), .Y(n_567) );
INVx6_ASAP7_75t_SL g568 ( .A(n_467), .Y(n_568) );
AOI221x1_ASAP7_75t_L g569 ( .A1(n_494), .A2(n_169), .B1(n_170), .B2(n_171), .C(n_175), .Y(n_569) );
CKINVDCx16_ASAP7_75t_R g570 ( .A(n_492), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_497), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_505), .B(n_462), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_442), .A2(n_429), .B(n_503), .Y(n_573) );
NOR2x1_ASAP7_75t_R g574 ( .A(n_434), .B(n_478), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_481), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_476), .Y(n_576) );
AOI21x1_ASAP7_75t_L g577 ( .A1(n_489), .A2(n_404), .B(n_487), .Y(n_577) );
OAI21x1_ASAP7_75t_L g578 ( .A1(n_489), .A2(n_487), .B(n_404), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_489), .Y(n_579) );
BUFx2_ASAP7_75t_L g580 ( .A(n_506), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_440), .B(n_365), .Y(n_581) );
AO31x2_ASAP7_75t_L g582 ( .A1(n_483), .A2(n_480), .A3(n_439), .B(n_487), .Y(n_582) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_440), .Y(n_583) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_506), .Y(n_584) );
NAND2x1_ASAP7_75t_L g585 ( .A(n_452), .B(n_438), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_487), .A2(n_404), .B(n_384), .Y(n_586) );
BUFx3_ASAP7_75t_L g587 ( .A(n_506), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_435), .B(n_437), .Y(n_588) );
AO31x2_ASAP7_75t_L g589 ( .A1(n_483), .A2(n_480), .A3(n_439), .B(n_487), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_487), .A2(n_404), .B(n_384), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_452), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_487), .A2(n_404), .B(n_384), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_487), .A2(n_404), .B(n_384), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_435), .B(n_437), .Y(n_594) );
AOI21x1_ASAP7_75t_L g595 ( .A1(n_487), .A2(n_404), .B(n_483), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g596 ( .A1(n_432), .A2(n_439), .B(n_421), .Y(n_596) );
OAI22xp33_ASAP7_75t_L g597 ( .A1(n_506), .A2(n_386), .B1(n_375), .B2(n_418), .Y(n_597) );
OAI21x1_ASAP7_75t_L g598 ( .A1(n_487), .A2(n_404), .B(n_493), .Y(n_598) );
AOI211x1_ASAP7_75t_L g599 ( .A1(n_459), .A2(n_498), .B(n_390), .C(n_394), .Y(n_599) );
INVx2_ASAP7_75t_SL g600 ( .A(n_506), .Y(n_600) );
BUFx10_ASAP7_75t_L g601 ( .A(n_440), .Y(n_601) );
AOI221xp5_ASAP7_75t_L g602 ( .A1(n_464), .A2(n_406), .B1(n_468), .B2(n_430), .C(n_367), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_558), .B(n_513), .Y(n_603) );
INVx3_ASAP7_75t_L g604 ( .A(n_585), .Y(n_604) );
AO31x2_ASAP7_75t_L g605 ( .A1(n_586), .A2(n_590), .A3(n_593), .B(n_592), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_588), .A2(n_561), .B1(n_511), .B2(n_599), .Y(n_606) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_510), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_594), .B(n_602), .Y(n_608) );
OA21x2_ASAP7_75t_L g609 ( .A1(n_529), .A2(n_569), .B(n_546), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_594), .B(n_540), .Y(n_610) );
NAND2x1p5_ASAP7_75t_L g611 ( .A(n_559), .B(n_584), .Y(n_611) );
CKINVDCx6p67_ASAP7_75t_R g612 ( .A(n_587), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_516), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_583), .B(n_545), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_519), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_531), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_576), .A2(n_536), .B(n_530), .Y(n_617) );
BUFx12f_ASAP7_75t_L g618 ( .A(n_537), .Y(n_618) );
INVx3_ASAP7_75t_L g619 ( .A(n_559), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_543), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_547), .B(n_550), .Y(n_621) );
BUFx10_ASAP7_75t_L g622 ( .A(n_517), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_554), .Y(n_623) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_528), .Y(n_624) );
NAND2x1p5_ASAP7_75t_L g625 ( .A(n_559), .B(n_544), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_556), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_570), .B(n_527), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_597), .B(n_522), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_523), .B(n_571), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_534), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_572), .B(n_548), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_553), .B(n_591), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_539), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_525), .A2(n_562), .B(n_573), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_533), .Y(n_635) );
INVx4_ASAP7_75t_SL g636 ( .A(n_552), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_580), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_601), .B(n_600), .Y(n_638) );
BUFx3_ASAP7_75t_L g639 ( .A(n_538), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_518), .B(n_566), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_574), .B(n_542), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_567), .A2(n_563), .B1(n_521), .B2(n_541), .Y(n_642) );
AND2x6_ASAP7_75t_L g643 ( .A(n_528), .B(n_551), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_567), .A2(n_524), .B1(n_565), .B2(n_568), .Y(n_644) );
OA21x2_ASAP7_75t_L g645 ( .A1(n_560), .A2(n_564), .B(n_532), .Y(n_645) );
CKINVDCx6p67_ASAP7_75t_R g646 ( .A(n_531), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_582), .B(n_589), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_582), .B(n_589), .Y(n_648) );
BUFx8_ASAP7_75t_L g649 ( .A(n_526), .Y(n_649) );
OR2x6_ASAP7_75t_L g650 ( .A(n_549), .B(n_535), .Y(n_650) );
AO21x2_ASAP7_75t_L g651 ( .A1(n_512), .A2(n_582), .B(n_557), .Y(n_651) );
NAND2x1p5_ASAP7_75t_L g652 ( .A(n_535), .B(n_515), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_535), .B(n_515), .Y(n_653) );
OA21x2_ASAP7_75t_L g654 ( .A1(n_514), .A2(n_520), .B(n_515), .Y(n_654) );
OA21x2_ASAP7_75t_L g655 ( .A1(n_520), .A2(n_579), .B(n_578), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_526), .B(n_558), .Y(n_656) );
OA21x2_ASAP7_75t_L g657 ( .A1(n_526), .A2(n_579), .B(n_578), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_513), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_596), .A2(n_412), .B(n_439), .Y(n_659) );
OA21x2_ASAP7_75t_L g660 ( .A1(n_579), .A2(n_578), .B(n_598), .Y(n_660) );
NAND2x1p5_ASAP7_75t_L g661 ( .A(n_559), .B(n_438), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_513), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_558), .B(n_435), .Y(n_663) );
BUFx3_ASAP7_75t_L g664 ( .A(n_584), .Y(n_664) );
AOI21xp33_ASAP7_75t_SL g665 ( .A1(n_552), .A2(n_402), .B(n_299), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_594), .B(n_435), .Y(n_666) );
INVx2_ASAP7_75t_SL g667 ( .A(n_584), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_583), .B(n_440), .Y(n_668) );
AOI21xp33_ASAP7_75t_L g669 ( .A1(n_558), .A2(n_575), .B(n_555), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_558), .A2(n_447), .B1(n_386), .B2(n_420), .Y(n_670) );
INVx3_ASAP7_75t_L g671 ( .A(n_585), .Y(n_671) );
AND2x4_ASAP7_75t_L g672 ( .A(n_594), .B(n_435), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_510), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_581), .B(n_440), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_594), .B(n_435), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_558), .B(n_435), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_581), .B(n_440), .Y(n_677) );
INVxp67_ASAP7_75t_SL g678 ( .A(n_583), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_594), .B(n_435), .Y(n_679) );
INVx3_ASAP7_75t_L g680 ( .A(n_585), .Y(n_680) );
INVx3_ASAP7_75t_L g681 ( .A(n_585), .Y(n_681) );
INVx8_ASAP7_75t_L g682 ( .A(n_527), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_513), .Y(n_683) );
AOI21x1_ASAP7_75t_L g684 ( .A1(n_577), .A2(n_595), .B(n_579), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_623), .B(n_626), .Y(n_685) );
OR2x6_ASAP7_75t_L g686 ( .A(n_644), .B(n_682), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_617), .B(n_624), .Y(n_687) );
INVx4_ASAP7_75t_L g688 ( .A(n_682), .Y(n_688) );
BUFx3_ASAP7_75t_L g689 ( .A(n_682), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_608), .B(n_656), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_605), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_608), .B(n_656), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_605), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_660), .Y(n_694) );
OR2x6_ASAP7_75t_L g695 ( .A(n_644), .B(n_606), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_670), .B(n_658), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_674), .B(n_677), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_670), .B(n_662), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_603), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_683), .B(n_663), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_652), .Y(n_701) );
OR2x6_ASAP7_75t_L g702 ( .A(n_606), .B(n_650), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_668), .Y(n_703) );
BUFx2_ASAP7_75t_L g704 ( .A(n_649), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_663), .B(n_676), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_652), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_610), .B(n_666), .Y(n_707) );
OR2x6_ASAP7_75t_L g708 ( .A(n_650), .B(n_625), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_610), .B(n_666), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_678), .B(n_631), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_631), .B(n_628), .Y(n_711) );
AO21x2_ASAP7_75t_L g712 ( .A1(n_617), .A2(n_647), .B(n_648), .Y(n_712) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_672), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_621), .B(n_672), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_653), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_654), .Y(n_716) );
BUFx2_ASAP7_75t_L g717 ( .A(n_649), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_654), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_675), .B(n_679), .Y(n_719) );
INVx2_ASAP7_75t_SL g720 ( .A(n_611), .Y(n_720) );
AO21x2_ASAP7_75t_L g721 ( .A1(n_648), .A2(n_684), .B(n_659), .Y(n_721) );
AO21x2_ASAP7_75t_L g722 ( .A1(n_669), .A2(n_651), .B(n_634), .Y(n_722) );
AO21x2_ASAP7_75t_L g723 ( .A1(n_669), .A2(n_651), .B(n_634), .Y(n_723) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_607), .Y(n_724) );
BUFx4f_ASAP7_75t_SL g725 ( .A(n_618), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_613), .B(n_615), .Y(n_726) );
OR2x6_ASAP7_75t_L g727 ( .A(n_642), .B(n_661), .Y(n_727) );
INVx3_ASAP7_75t_L g728 ( .A(n_643), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_657), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_614), .B(n_629), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_657), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_655), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_630), .B(n_633), .Y(n_733) );
BUFx3_ASAP7_75t_L g734 ( .A(n_661), .Y(n_734) );
BUFx3_ASAP7_75t_L g735 ( .A(n_643), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_632), .B(n_635), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_673), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_620), .B(n_641), .Y(n_738) );
INVx3_ASAP7_75t_L g739 ( .A(n_619), .Y(n_739) );
OR2x6_ASAP7_75t_L g740 ( .A(n_604), .B(n_681), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_710), .B(n_641), .Y(n_741) );
BUFx2_ASAP7_75t_L g742 ( .A(n_708), .Y(n_742) );
OR2x2_ASAP7_75t_L g743 ( .A(n_710), .B(n_627), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_686), .B(n_680), .Y(n_744) );
BUFx3_ASAP7_75t_L g745 ( .A(n_689), .Y(n_745) );
BUFx3_ASAP7_75t_L g746 ( .A(n_689), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_715), .B(n_609), .Y(n_747) );
BUFx2_ASAP7_75t_L g748 ( .A(n_686), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_696), .B(n_680), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_694), .Y(n_750) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_724), .Y(n_751) );
AND2x4_ASAP7_75t_L g752 ( .A(n_686), .B(n_671), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_729), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_700), .B(n_637), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_730), .B(n_622), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_731), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_731), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_698), .B(n_622), .Y(n_758) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_737), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_695), .B(n_645), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_695), .B(n_645), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_733), .B(n_667), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_716), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_695), .B(n_664), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_716), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_718), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_726), .B(n_616), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_726), .B(n_640), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_736), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_701), .B(n_639), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_718), .Y(n_771) );
OR2x2_ASAP7_75t_L g772 ( .A(n_690), .B(n_638), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_706), .B(n_646), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_711), .B(n_665), .Y(n_774) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_736), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_732), .Y(n_776) );
AND2x4_ASAP7_75t_L g777 ( .A(n_704), .B(n_636), .Y(n_777) );
INVxp67_ASAP7_75t_L g778 ( .A(n_703), .Y(n_778) );
NAND2x1p5_ASAP7_75t_L g779 ( .A(n_734), .B(n_636), .Y(n_779) );
OR2x2_ASAP7_75t_L g780 ( .A(n_692), .B(n_612), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_732), .Y(n_781) );
CKINVDCx16_ASAP7_75t_R g782 ( .A(n_688), .Y(n_782) );
AND2x4_ASAP7_75t_L g783 ( .A(n_717), .B(n_687), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_699), .B(n_707), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_709), .B(n_685), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_709), .B(n_685), .Y(n_786) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_714), .Y(n_787) );
OR2x2_ASAP7_75t_L g788 ( .A(n_692), .B(n_705), .Y(n_788) );
NOR2x1_ASAP7_75t_SL g789 ( .A(n_727), .B(n_740), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_760), .B(n_712), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_760), .B(n_712), .Y(n_791) );
OR2x2_ASAP7_75t_L g792 ( .A(n_788), .B(n_717), .Y(n_792) );
OR2x2_ASAP7_75t_L g793 ( .A(n_788), .B(n_702), .Y(n_793) );
AND2x2_ASAP7_75t_L g794 ( .A(n_761), .B(n_712), .Y(n_794) );
OR2x2_ASAP7_75t_L g795 ( .A(n_741), .B(n_702), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_741), .B(n_702), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_761), .B(n_722), .Y(n_797) );
HB1xp67_ASAP7_75t_L g798 ( .A(n_751), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_785), .B(n_722), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_785), .B(n_722), .Y(n_800) );
OR2x2_ASAP7_75t_L g801 ( .A(n_769), .B(n_702), .Y(n_801) );
OR2x2_ASAP7_75t_L g802 ( .A(n_775), .B(n_723), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_786), .B(n_723), .Y(n_803) );
AND2x4_ASAP7_75t_L g804 ( .A(n_789), .B(n_687), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_749), .B(n_691), .Y(n_805) );
INVxp67_ASAP7_75t_L g806 ( .A(n_759), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_750), .Y(n_807) );
AND2x4_ASAP7_75t_L g808 ( .A(n_789), .B(n_687), .Y(n_808) );
OR2x2_ASAP7_75t_L g809 ( .A(n_787), .B(n_693), .Y(n_809) );
OR2x2_ASAP7_75t_L g810 ( .A(n_754), .B(n_721), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_782), .B(n_697), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_784), .B(n_721), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_753), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_753), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_756), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_799), .B(n_747), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_800), .B(n_757), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_807), .Y(n_818) );
INVx1_ASAP7_75t_SL g819 ( .A(n_792), .Y(n_819) );
INVxp67_ASAP7_75t_L g820 ( .A(n_811), .Y(n_820) );
AND2x4_ASAP7_75t_L g821 ( .A(n_804), .B(n_748), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_803), .B(n_763), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_798), .B(n_778), .Y(n_823) );
OR2x2_ASAP7_75t_L g824 ( .A(n_810), .B(n_765), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_790), .B(n_766), .Y(n_825) );
AND2x4_ASAP7_75t_L g826 ( .A(n_804), .B(n_783), .Y(n_826) );
INVx1_ASAP7_75t_SL g827 ( .A(n_792), .Y(n_827) );
INVx1_ASAP7_75t_SL g828 ( .A(n_809), .Y(n_828) );
OR2x2_ASAP7_75t_L g829 ( .A(n_812), .B(n_766), .Y(n_829) );
OR2x2_ASAP7_75t_L g830 ( .A(n_802), .B(n_771), .Y(n_830) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_806), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_790), .B(n_771), .Y(n_832) );
INVx3_ASAP7_75t_L g833 ( .A(n_804), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_791), .B(n_776), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_791), .B(n_776), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_794), .B(n_781), .Y(n_836) );
INVxp67_ASAP7_75t_SL g837 ( .A(n_809), .Y(n_837) );
AND2x2_ASAP7_75t_L g838 ( .A(n_797), .B(n_783), .Y(n_838) );
NOR2x1_ASAP7_75t_L g839 ( .A(n_833), .B(n_777), .Y(n_839) );
INVx4_ASAP7_75t_L g840 ( .A(n_833), .Y(n_840) );
INVxp67_ASAP7_75t_L g841 ( .A(n_831), .Y(n_841) );
OAI32xp33_ASAP7_75t_L g842 ( .A1(n_819), .A2(n_779), .A3(n_801), .B1(n_745), .B2(n_746), .Y(n_842) );
NAND2x1p5_ASAP7_75t_L g843 ( .A(n_826), .B(n_745), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_822), .B(n_813), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_825), .B(n_814), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_818), .Y(n_846) );
NAND3xp33_ASAP7_75t_SL g847 ( .A(n_827), .B(n_779), .C(n_780), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_832), .B(n_814), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_816), .B(n_805), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_832), .B(n_815), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_834), .B(n_815), .Y(n_851) );
AOI21xp33_ASAP7_75t_L g852 ( .A1(n_841), .A2(n_823), .B(n_780), .Y(n_852) );
OAI32xp33_ASAP7_75t_L g853 ( .A1(n_840), .A2(n_820), .A3(n_828), .B1(n_829), .B2(n_779), .Y(n_853) );
INVxp67_ASAP7_75t_L g854 ( .A(n_841), .Y(n_854) );
NAND3xp33_ASAP7_75t_L g855 ( .A(n_840), .B(n_830), .C(n_824), .Y(n_855) );
O2A1O1Ixp33_ASAP7_75t_L g856 ( .A1(n_847), .A2(n_774), .B(n_755), .C(n_767), .Y(n_856) );
INVx2_ASAP7_75t_SL g857 ( .A(n_843), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_844), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_846), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_843), .A2(n_826), .B1(n_821), .B2(n_837), .Y(n_860) );
AOI21xp5_ASAP7_75t_L g861 ( .A1(n_842), .A2(n_821), .B(n_808), .Y(n_861) );
AND2x4_ASAP7_75t_L g862 ( .A(n_839), .B(n_821), .Y(n_862) );
NOR2xp33_ASAP7_75t_L g863 ( .A(n_854), .B(n_852), .Y(n_863) );
NOR3xp33_ASAP7_75t_L g864 ( .A(n_856), .B(n_773), .C(n_762), .Y(n_864) );
AOI221xp5_ASAP7_75t_L g865 ( .A1(n_855), .A2(n_848), .B1(n_851), .B2(n_850), .C(n_845), .Y(n_865) );
OAI21xp33_ASAP7_75t_L g866 ( .A1(n_860), .A2(n_817), .B(n_849), .Y(n_866) );
OAI211xp5_ASAP7_75t_SL g867 ( .A1(n_861), .A2(n_772), .B(n_768), .C(n_725), .Y(n_867) );
OAI22xp33_ASAP7_75t_SL g868 ( .A1(n_857), .A2(n_793), .B1(n_796), .B2(n_795), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_858), .A2(n_835), .B1(n_836), .B2(n_838), .Y(n_869) );
NAND4xp25_ASAP7_75t_L g870 ( .A(n_853), .B(n_764), .C(n_758), .D(n_772), .Y(n_870) );
OAI22xp5_ASAP7_75t_SL g871 ( .A1(n_862), .A2(n_688), .B1(n_743), .B2(n_742), .Y(n_871) );
AOI211xp5_ASAP7_75t_L g872 ( .A1(n_862), .A2(n_744), .B(n_752), .C(n_793), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_863), .B(n_865), .Y(n_873) );
NAND3xp33_ASAP7_75t_SL g874 ( .A(n_866), .B(n_864), .C(n_872), .Y(n_874) );
NOR2x1_ASAP7_75t_L g875 ( .A(n_867), .B(n_870), .Y(n_875) );
NOR3xp33_ASAP7_75t_L g876 ( .A(n_874), .B(n_871), .C(n_868), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_875), .B(n_869), .Y(n_877) );
NOR3xp33_ASAP7_75t_L g878 ( .A(n_873), .B(n_739), .C(n_728), .Y(n_878) );
AND2x4_ASAP7_75t_L g879 ( .A(n_878), .B(n_876), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_877), .Y(n_880) );
AOI31xp33_ASAP7_75t_L g881 ( .A1(n_880), .A2(n_770), .A3(n_713), .B(n_720), .Y(n_881) );
NOR2x1_ASAP7_75t_L g882 ( .A(n_879), .B(n_735), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_881), .Y(n_883) );
INVx3_ASAP7_75t_L g884 ( .A(n_882), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_883), .B(n_859), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_885), .B(n_884), .Y(n_886) );
XNOR2xp5_ASAP7_75t_L g887 ( .A(n_886), .B(n_719), .Y(n_887) );
NAND2xp5_ASAP7_75t_SL g888 ( .A(n_887), .B(n_735), .Y(n_888) );
AOI21xp33_ASAP7_75t_SL g889 ( .A1(n_888), .A2(n_738), .B(n_728), .Y(n_889) );
endmodule