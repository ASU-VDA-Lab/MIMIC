module fake_jpeg_2141_n_71 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_71);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_71;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

BUFx24_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_31),
.Y(n_35)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_23),
.B1(n_22),
.B2(n_26),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_37),
.B1(n_31),
.B2(n_25),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_22),
.B(n_21),
.C(n_25),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_35),
.C(n_33),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_31),
.B1(n_28),
.B2(n_21),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_33),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

BUFx2_ASAP7_75t_SL g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_19),
.C(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_48),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_17),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_1),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_57),
.B(n_55),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

AO22x1_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_56)
);

AO22x1_ASAP7_75t_SL g60 ( 
.A1(n_56),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_60)
);

OAI211xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_47),
.B(n_48),
.C(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_60),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

A2O1A1O1Ixp25_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_56),
.B(n_55),
.C(n_57),
.D(n_10),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_60),
.C(n_62),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_65),
.C(n_63),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_SL g68 ( 
.A1(n_67),
.A2(n_61),
.B(n_12),
.C(n_11),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_9),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_69),
.A2(n_9),
.B(n_10),
.Y(n_70)
);

BUFx24_ASAP7_75t_SL g71 ( 
.A(n_70),
.Y(n_71)
);


endmodule