module fake_jpeg_1687_n_92 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_92);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_92;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_11),
.B(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_5),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_22),
.A2(n_18),
.B1(n_15),
.B2(n_20),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_40),
.B1(n_4),
.B2(n_8),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_21),
.B1(n_13),
.B2(n_3),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_21),
.B1(n_4),
.B2(n_1),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_1),
.B(n_4),
.Y(n_50)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_29),
.B1(n_25),
.B2(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_34),
.B(n_40),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_34),
.B1(n_42),
.B2(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_8),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_44),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_44),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_50),
.B(n_48),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_48),
.B1(n_57),
.B2(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_65),
.B(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_70),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_62),
.B1(n_61),
.B2(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_72),
.Y(n_76)
);

INVxp33_ASAP7_75t_SL g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_66),
.C(n_61),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_65),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_73),
.B1(n_47),
.B2(n_59),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_77),
.A2(n_69),
.B1(n_74),
.B2(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_76),
.C(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_83),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_81),
.C(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_88),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_76),
.A3(n_83),
.B1(n_59),
.B2(n_60),
.C1(n_56),
.C2(n_42),
.Y(n_88)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_85),
.A3(n_60),
.B1(n_56),
.B2(n_42),
.C1(n_64),
.C2(n_33),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_90),
.A2(n_60),
.B(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_46),
.Y(n_92)
);


endmodule