module fake_jpeg_20801_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_43),
.Y(n_46)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_22),
.B1(n_33),
.B2(n_20),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_37),
.B1(n_40),
.B2(n_36),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_63),
.B(n_71),
.Y(n_105)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_57),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_75),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_80),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_78),
.A2(n_93),
.B1(n_51),
.B2(n_55),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_40),
.B1(n_22),
.B2(n_44),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_82),
.B1(n_31),
.B2(n_21),
.Y(n_109)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_44),
.B1(n_22),
.B2(n_33),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_87),
.B1(n_51),
.B2(n_16),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_22),
.B1(n_33),
.B2(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_88),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_17),
.B1(n_26),
.B2(n_29),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_17),
.B1(n_26),
.B2(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_16),
.B1(n_21),
.B2(n_25),
.Y(n_89)
);

AOI32xp33_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_30),
.A3(n_32),
.B1(n_16),
.B2(n_25),
.Y(n_100)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_43),
.C(n_45),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_43),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_30),
.B1(n_17),
.B2(n_32),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_102),
.B(n_89),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_43),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_73),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_109),
.B1(n_114),
.B2(n_115),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_106),
.A2(n_71),
.B1(n_68),
.B2(n_91),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_74),
.A2(n_47),
.B1(n_30),
.B2(n_32),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_112),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_64),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_69),
.A2(n_38),
.B1(n_21),
.B2(n_31),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_31),
.B1(n_25),
.B2(n_18),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_64),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_118),
.Y(n_149)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_28),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_28),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_125),
.B1(n_124),
.B2(n_119),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_128),
.A2(n_151),
.B1(n_121),
.B2(n_28),
.Y(n_176)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_115),
.B(n_109),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_95),
.C(n_83),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_74),
.C(n_70),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_143),
.C(n_99),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_139),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_67),
.B1(n_65),
.B2(n_80),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_121),
.B1(n_97),
.B2(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_84),
.C(n_91),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_90),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_110),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_97),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_43),
.B(n_34),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_153),
.A2(n_34),
.B(n_104),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_84),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_66),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_149),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_155),
.B(n_173),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_112),
.B1(n_117),
.B2(n_100),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_161),
.B1(n_163),
.B2(n_178),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_157),
.A2(n_159),
.B(n_164),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_182),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_145),
.B(n_153),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_162),
.A2(n_172),
.B(n_3),
.Y(n_218)
);

OAI22x1_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_96),
.B1(n_88),
.B2(n_101),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_152),
.A2(n_101),
.B(n_118),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_171),
.C(n_166),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_96),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_170),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_0),
.B(n_1),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_126),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_140),
.B1(n_146),
.B2(n_137),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_135),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_131),
.A2(n_27),
.B1(n_24),
.B2(n_2),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_179),
.A2(n_180),
.B1(n_3),
.B2(n_4),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_131),
.A2(n_27),
.B1(n_24),
.B2(n_2),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_0),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_0),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_186),
.Y(n_209)
);

AO22x1_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_1),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_187),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_196),
.B1(n_180),
.B2(n_179),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_165),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_191),
.B(n_198),
.Y(n_227)
);

A2O1A1O1Ixp25_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_136),
.B(n_143),
.C(n_126),
.D(n_133),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_192),
.B(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_185),
.A2(n_130),
.B1(n_129),
.B2(n_139),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_148),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_206),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_174),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_147),
.A3(n_141),
.B1(n_15),
.B2(n_14),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_169),
.C(n_183),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_15),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_167),
.B(n_14),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_210),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

INVxp67_ASAP7_75t_SL g238 ( 
.A(n_211),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_176),
.A2(n_13),
.B(n_4),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_233)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

OAI22x1_ASAP7_75t_SL g216 ( 
.A1(n_159),
.A2(n_164),
.B1(n_186),
.B2(n_167),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_5),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_166),
.B(n_182),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_222),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_224),
.C(n_244),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_184),
.B1(n_181),
.B2(n_161),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_223),
.A2(n_231),
.B1(n_235),
.B2(n_237),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_187),
.C(n_184),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_187),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_230),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_172),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_202),
.A2(n_181),
.B1(n_186),
.B2(n_6),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_195),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_237)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_192),
.B(n_199),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_236),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_190),
.B(n_13),
.C(n_8),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_216),
.B1(n_197),
.B2(n_196),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_247),
.B1(n_248),
.B2(n_222),
.Y(n_268)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_189),
.C(n_194),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_246),
.A2(n_250),
.B(n_8),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_227),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_197),
.B1(n_188),
.B2(n_209),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_200),
.B(n_201),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_253),
.B(n_226),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_226),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_263),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_242),
.B(n_193),
.CI(n_209),
.CON(n_257),
.SN(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_213),
.C(n_203),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_262),
.C(n_265),
.Y(n_267)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_259),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_218),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_264),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_215),
.C(n_193),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_228),
.B(n_220),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_219),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_7),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_244),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_279),
.Y(n_298)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_275),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_281),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_243),
.C(n_234),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_283),
.C(n_262),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_231),
.B1(n_225),
.B2(n_240),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_280),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_251),
.B(n_253),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_240),
.B1(n_243),
.B2(n_237),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_252),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_282),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_9),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_270),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_284),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_272),
.A2(n_248),
.B(n_245),
.Y(n_287)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_294),
.C(n_285),
.Y(n_306)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_274),
.A2(n_257),
.B(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_266),
.A2(n_257),
.B(n_251),
.Y(n_292)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_256),
.C(n_11),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_267),
.C(n_283),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g295 ( 
.A(n_275),
.B(n_10),
.CI(n_12),
.CON(n_295),
.SN(n_295)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_271),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_273),
.A2(n_10),
.B(n_12),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_12),
.B(n_290),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_299),
.B(n_306),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_305),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_277),
.C(n_279),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_277),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_310),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_278),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_308),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_12),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_295),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_311),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_305),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_293),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_317),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_290),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_302),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_304),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_323),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_298),
.C(n_309),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_325),
.C(n_319),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_286),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_328),
.B(n_320),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_315),
.B(n_291),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_327),
.B(n_322),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_325),
.C(n_289),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_289),
.Y(n_334)
);


endmodule