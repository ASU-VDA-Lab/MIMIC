module fake_jpeg_3503_n_44 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_4),
.B(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_6),
.B(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_19),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_31)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_25),
.C(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx2_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_9),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_31),
.C(n_21),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_25),
.Y(n_32)
);

XOR2x2_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_21),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_30),
.B1(n_23),
.B2(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_20),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_27),
.B1(n_18),
.B2(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_26),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

NAND2xp67_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_24),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_40),
.A2(n_37),
.B1(n_12),
.B2(n_29),
.Y(n_42)
);

AOI322xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_13),
.A3(n_14),
.B1(n_17),
.B2(n_35),
.C1(n_36),
.C2(n_42),
.Y(n_43)
);

NAND4xp25_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_17),
.C(n_30),
.D(n_35),
.Y(n_44)
);


endmodule