module fake_jpeg_21836_n_109 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_26),
.B(n_34),
.Y(n_47)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_35),
.Y(n_45)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_30),
.A2(n_12),
.B1(n_16),
.B2(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

NAND2x1p5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_49),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_57),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_55),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_43),
.B1(n_27),
.B2(n_32),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_64),
.B1(n_18),
.B2(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_12),
.B1(n_29),
.B2(n_22),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_14),
.Y(n_63)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_21),
.B1(n_20),
.B2(n_18),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_47),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_50),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_47),
.C(n_61),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_74),
.C(n_75),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_49),
.B1(n_47),
.B2(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_75),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_45),
.B(n_20),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_45),
.B1(n_15),
.B2(n_31),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_13),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_78),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_50),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_81),
.B(n_84),
.Y(n_87)
);

MAJx2_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_52),
.C(n_31),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_65),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_58),
.B1(n_70),
.B2(n_53),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_92),
.C(n_86),
.Y(n_94)
);

XNOR2x2_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_80),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_25),
.Y(n_97)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_89),
.B(n_68),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_66),
.B1(n_86),
.B2(n_57),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_74),
.B(n_70),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_97),
.B(n_15),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_95),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_67),
.C(n_85),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_14),
.B(n_25),
.Y(n_99)
);

AO21x1_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_7),
.B(n_9),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_101),
.Y(n_104)
);

AOI32xp33_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_25),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_100),
.B(n_1),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_9),
.B(n_104),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_106),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);


endmodule