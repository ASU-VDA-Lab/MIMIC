module fake_jpeg_861_n_214 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_214);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_31),
.Y(n_63)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

INVx11_ASAP7_75t_SL g67 ( 
.A(n_21),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_18),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_19),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_12),
.Y(n_77)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_1),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_1),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_65),
.B(n_75),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_86),
.B1(n_80),
.B2(n_79),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_96),
.B1(n_101),
.B2(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_69),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_62),
.B1(n_79),
.B2(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_75),
.B1(n_77),
.B2(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_105),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_72),
.B(n_55),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_104),
.B(n_107),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_64),
.B(n_72),
.C(n_56),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_76),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_60),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_78),
.B1(n_64),
.B2(n_73),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_60),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_57),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_115),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_54),
.C(n_69),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_114),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_58),
.C(n_63),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_29),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_56),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_120),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_114),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_138),
.B1(n_142),
.B2(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_132),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_78),
.B(n_73),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_7),
.B(n_8),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_120),
.Y(n_132)
);

OR2x6_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_60),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_134),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_62),
.B1(n_3),
.B2(n_4),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_6),
.Y(n_148)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_105),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_13),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_148),
.B(n_156),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_28),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_150),
.C(n_159),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_160),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_30),
.B1(n_52),
.B2(n_51),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_159),
.B1(n_164),
.B2(n_168),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_133),
.B1(n_141),
.B2(n_130),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_154),
.A2(n_36),
.B(n_35),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_7),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_27),
.B1(n_48),
.B2(n_47),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_13),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_162),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_26),
.B1(n_45),
.B2(n_42),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_165),
.B(n_53),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_123),
.B(n_136),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_32),
.B(n_23),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_25),
.B1(n_41),
.B2(n_40),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_39),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_174),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_162),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_173),
.A2(n_179),
.B(n_168),
.Y(n_190)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_33),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_176),
.B(n_182),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_178),
.A2(n_180),
.B1(n_167),
.B2(n_157),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_155),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_175),
.B(n_149),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_188),
.B(n_194),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_151),
.B(n_164),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_190),
.B(n_178),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_179),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_193),
.B1(n_183),
.B2(n_153),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_173),
.B1(n_176),
.B2(n_184),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_177),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_186),
.B(n_182),
.CI(n_147),
.CON(n_195),
.SN(n_195)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_199),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_171),
.C(n_145),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_198),
.C(n_189),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_173),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_201),
.Y(n_204)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_203),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_204),
.A2(n_201),
.B1(n_195),
.B2(n_191),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_206),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_185),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_209),
.A2(n_207),
.B(n_205),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_211),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_206),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_18),
.Y(n_214)
);


endmodule