module fake_jpeg_20073_n_238 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_31),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_21),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_33),
.Y(n_82)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_23),
.B1(n_32),
.B2(n_30),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_53),
.A2(n_64),
.B1(n_68),
.B2(n_29),
.Y(n_90)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_65),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_23),
.B1(n_30),
.B2(n_17),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_59),
.A2(n_61),
.B1(n_9),
.B2(n_10),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_23),
.B1(n_17),
.B2(n_28),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_18),
.B(n_28),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_3),
.B(n_4),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_71),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_18),
.B1(n_27),
.B2(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_22),
.Y(n_65)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_69),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_27),
.B1(n_20),
.B2(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_22),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_39),
.B(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_20),
.Y(n_72)
);

NAND2x2_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_33),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_29),
.B(n_24),
.C(n_19),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_15),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_13),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_29),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_98),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_73),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_92),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_56),
.B(n_62),
.C(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_77),
.B(n_79),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_1),
.B(n_2),
.Y(n_78)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_78),
.A2(n_86),
.B(n_91),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_15),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_33),
.B1(n_24),
.B2(n_19),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_87),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_29),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_96),
.B1(n_101),
.B2(n_49),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_24),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_19),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_2),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_98),
.C(n_49),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_3),
.C(n_5),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_14),
.Y(n_112)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_58),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_109),
.B(n_111),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_58),
.B(n_51),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_48),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_99),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_67),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_91),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_126),
.B1(n_129),
.B2(n_131),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_125),
.B1(n_108),
.B2(n_127),
.Y(n_153)
);

OR2x4_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_12),
.Y(n_123)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_84),
.B(n_86),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_82),
.A2(n_96),
.B1(n_91),
.B2(n_87),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_132),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_94),
.B1(n_105),
.B2(n_88),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_81),
.A2(n_89),
.B1(n_85),
.B2(n_103),
.Y(n_131)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_130),
.B(n_106),
.Y(n_165)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_104),
.C(n_85),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_118),
.C(n_106),
.Y(n_160)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_99),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_143),
.B(n_146),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_92),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_144),
.B(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_147),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_83),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_83),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_121),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_130),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_150),
.B1(n_111),
.B2(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_155),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_132),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_154),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_177),
.C(n_133),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_171),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_164),
.A2(n_165),
.B(n_168),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_149),
.A2(n_111),
.B1(n_148),
.B2(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_167),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_125),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_120),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_170),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_122),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_131),
.B(n_137),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_174),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_141),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_172),
.C(n_168),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_162),
.B(n_134),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_181),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_148),
.B1(n_157),
.B2(n_152),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_157),
.B1(n_156),
.B2(n_137),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_185),
.B1(n_166),
.B2(n_169),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_151),
.B1(n_136),
.B2(n_139),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_135),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_193),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_135),
.Y(n_193)
);

INVxp33_ASAP7_75t_SL g196 ( 
.A(n_184),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_183),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_160),
.C(n_177),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_197),
.B(n_206),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_184),
.A2(n_167),
.B(n_162),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_201),
.B(n_187),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_163),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_204),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_190),
.A2(n_186),
.B(n_175),
.Y(n_201)
);

OAI321xp33_ASAP7_75t_L g205 ( 
.A1(n_180),
.A2(n_175),
.A3(n_168),
.B1(n_161),
.B2(n_138),
.C(n_158),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_182),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_209),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_195),
.B(n_185),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_212),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_194),
.B(n_192),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_204),
.B(n_190),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_215),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_179),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_187),
.C(n_202),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_194),
.B1(n_179),
.B2(n_203),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_222),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_213),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_216),
.A2(n_201),
.B1(n_200),
.B2(n_188),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_221),
.A2(n_189),
.B(n_169),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_227),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_217),
.B(n_213),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_226),
.B(n_220),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_142),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_214),
.C(n_223),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_225),
.B(n_223),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_232),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_218),
.B(n_138),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_235),
.A2(n_228),
.B1(n_218),
.B2(n_145),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_237),
.C(n_233),
.Y(n_238)
);


endmodule