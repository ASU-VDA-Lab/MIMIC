module fake_netlist_6_3246_n_1488 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_376, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_364, n_295, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1488);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_364;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1488;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_1371;
wire n_1285;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_1485;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_1408;
wire n_1196;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1109;
wire n_712;
wire n_1276;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_L g384 ( 
.A(n_103),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_221),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_252),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_276),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_172),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_288),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_353),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_284),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_312),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_36),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_240),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_31),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_109),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_366),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_177),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_346),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_304),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_359),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_6),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_188),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_63),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_344),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_333),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_295),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_331),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_97),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_134),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_41),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_143),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_235),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_230),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_47),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_150),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_377),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_124),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_52),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_0),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_264),
.B(n_335),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_110),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_75),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_285),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_94),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_327),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_350),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_20),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_78),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_374),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_247),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_130),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_380),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_123),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_347),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_302),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_33),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_99),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_261),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_94),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_37),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_148),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_233),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_112),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_220),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_292),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_314),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_370),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_281),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_187),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_41),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_375),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_64),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_12),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_51),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_325),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_82),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_311),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_117),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_297),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_202),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_339),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_125),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_330),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_92),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_107),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_149),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_255),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_319),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_206),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_140),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_256),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_334),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_267),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_263),
.B(n_128),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_300),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_3),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_28),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_303),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_315),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_141),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_243),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_345),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_47),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_298),
.B(n_153),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_207),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_251),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_10),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_277),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_273),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_234),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_260),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_289),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_114),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_205),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_100),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_169),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_164),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_106),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_167),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_357),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_232),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_5),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_163),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_342),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_L g509 ( 
.A(n_217),
.B(n_12),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_361),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_343),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_323),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_111),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_253),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_33),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_84),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_20),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_248),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_309),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_61),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_103),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_245),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_105),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_127),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_10),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_11),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_126),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_57),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_161),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_24),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_192),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_50),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_166),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_80),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_272),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_364),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_106),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_59),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_84),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_85),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_95),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_354),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_82),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_100),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_27),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_196),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_78),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_139),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_378),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_291),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_270),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_332),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_171),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_258),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_74),
.B(n_215),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_326),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_257),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_294),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_72),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_278),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_254),
.B(n_286),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_73),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_244),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_52),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_165),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_56),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_54),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_168),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_63),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_28),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_174),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_265),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_89),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_310),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_552),
.B(n_0),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_491),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_569),
.Y(n_577)
);

OAI22x1_ASAP7_75t_R g578 ( 
.A1(n_395),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_552),
.B(n_2),
.Y(n_579)
);

OA21x2_ASAP7_75t_L g580 ( 
.A1(n_388),
.A2(n_4),
.B(n_5),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_569),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_502),
.Y(n_582)
);

BUFx12f_ASAP7_75t_L g583 ( 
.A(n_386),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_502),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_394),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_502),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_502),
.Y(n_587)
);

BUFx8_ASAP7_75t_L g588 ( 
.A(n_447),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_414),
.B(n_4),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_425),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_590)
);

BUFx8_ASAP7_75t_L g591 ( 
.A(n_411),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_384),
.Y(n_592)
);

INVx6_ASAP7_75t_L g593 ( 
.A(n_386),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_393),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_411),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_432),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_462),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_414),
.B(n_7),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_415),
.B(n_8),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_462),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_394),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_415),
.B(n_442),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_497),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_396),
.Y(n_604)
);

OA21x2_ASAP7_75t_L g605 ( 
.A1(n_388),
.A2(n_9),
.B(n_11),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_497),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_442),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_394),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_394),
.Y(n_609)
);

BUFx8_ASAP7_75t_L g610 ( 
.A(n_534),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_448),
.Y(n_611)
);

AND2x2_ASAP7_75t_SL g612 ( 
.A(n_407),
.B(n_470),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_404),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_408),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_409),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_416),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_408),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_408),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_408),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_568),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_L g621 ( 
.A(n_570),
.B(n_13),
.Y(n_621)
);

OA21x2_ASAP7_75t_L g622 ( 
.A1(n_397),
.A2(n_13),
.B(n_14),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_402),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_422),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_426),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_472),
.B(n_15),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_538),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_547),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_547),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_423),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_428),
.B(n_16),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_562),
.Y(n_632)
);

AND2x6_ASAP7_75t_L g633 ( 
.A(n_568),
.B(n_119),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_397),
.B(n_17),
.Y(n_634)
);

OA21x2_ASAP7_75t_L g635 ( 
.A1(n_418),
.A2(n_18),
.B(n_19),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_448),
.B(n_18),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_431),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_562),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_441),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_567),
.Y(n_640)
);

AND2x6_ASAP7_75t_L g641 ( 
.A(n_568),
.B(n_120),
.Y(n_641)
);

BUFx8_ASAP7_75t_L g642 ( 
.A(n_567),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_563),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_443),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_548),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_563),
.B(n_21),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_440),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_418),
.B(n_22),
.Y(n_648)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_419),
.A2(n_122),
.B(n_121),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_456),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_481),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_499),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_419),
.B(n_23),
.Y(n_653)
);

BUFx12f_ASAP7_75t_L g654 ( 
.A(n_444),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_593),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_586),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_609),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_602),
.B(n_506),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_598),
.B(n_599),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_596),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_609),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_612),
.A2(n_406),
.B1(n_410),
.B2(n_390),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_607),
.B(n_515),
.Y(n_663)
);

INVx5_ASAP7_75t_L g664 ( 
.A(n_633),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_609),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_582),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_609),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_589),
.B(n_446),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_614),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_588),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_607),
.B(n_611),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_643),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_611),
.B(n_421),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_612),
.B(n_555),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_643),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_593),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_643),
.B(n_619),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_584),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_577),
.B(n_520),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_643),
.B(n_421),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_587),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_614),
.Y(n_682)
);

CKINVDCx6p67_ASAP7_75t_R g683 ( 
.A(n_583),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_588),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_601),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_601),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_633),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_575),
.B(n_387),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_619),
.B(n_438),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_601),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_591),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_589),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_625),
.B(n_539),
.C(n_469),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_608),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_608),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_608),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_617),
.Y(n_697)
);

NOR2x1p5_ASAP7_75t_L g698 ( 
.A(n_575),
.B(n_541),
.Y(n_698)
);

NOR2x1p5_ASAP7_75t_L g699 ( 
.A(n_579),
.B(n_424),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_617),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_626),
.B(n_509),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_617),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_581),
.Y(n_703)
);

CKINVDCx6p67_ASAP7_75t_R g704 ( 
.A(n_654),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_579),
.B(n_454),
.Y(n_705)
);

NAND3xp33_ASAP7_75t_L g706 ( 
.A(n_626),
.B(n_458),
.C(n_457),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_697),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_697),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_671),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_688),
.B(n_675),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_701),
.B(n_623),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_677),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_671),
.B(n_647),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_658),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_699),
.B(n_585),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_697),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_685),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_706),
.B(n_692),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_685),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_668),
.B(n_585),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_690),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_686),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_674),
.B(n_576),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_698),
.A2(n_645),
.B1(n_590),
.B2(n_634),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_668),
.B(n_585),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_668),
.B(n_585),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_658),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_692),
.B(n_636),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_700),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_692),
.B(n_636),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_659),
.B(n_698),
.Y(n_731)
);

OAI221xp5_ASAP7_75t_L g732 ( 
.A1(n_705),
.A2(n_653),
.B1(n_648),
.B2(n_621),
.C(n_594),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_693),
.A2(n_705),
.B1(n_660),
.B2(n_451),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_679),
.A2(n_605),
.B1(n_622),
.B2(n_580),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_672),
.B(n_618),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_694),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_667),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_673),
.B(n_646),
.Y(n_738)
);

O2A1O1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_680),
.A2(n_648),
.B(n_653),
.C(n_621),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_703),
.B(n_591),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_655),
.B(n_435),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_702),
.B(n_618),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_662),
.A2(n_514),
.B1(n_549),
.B2(n_473),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_694),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_679),
.A2(n_649),
.B(n_561),
.C(n_604),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_695),
.Y(n_746)
);

OR2x6_ASAP7_75t_L g747 ( 
.A(n_655),
.B(n_625),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_695),
.B(n_618),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_696),
.B(n_620),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_676),
.B(n_550),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_676),
.B(n_385),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_663),
.Y(n_752)
);

BUFx8_ASAP7_75t_L g753 ( 
.A(n_691),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_696),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_687),
.A2(n_605),
.B1(n_622),
.B2(n_580),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_663),
.B(n_595),
.Y(n_756)
);

NAND3xp33_ASAP7_75t_L g757 ( 
.A(n_703),
.B(n_642),
.C(n_610),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_689),
.B(n_610),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_691),
.B(n_595),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_704),
.B(n_650),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_657),
.B(n_665),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_704),
.A2(n_523),
.B1(n_650),
.B2(n_540),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_666),
.B(n_597),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_665),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_669),
.B(n_392),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_666),
.Y(n_766)
);

NAND2xp33_ASAP7_75t_SL g767 ( 
.A(n_687),
.B(n_460),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_664),
.B(n_633),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_678),
.B(n_681),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_661),
.B(n_437),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_731),
.B(n_687),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_739),
.A2(n_561),
.B(n_488),
.C(n_445),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_713),
.B(n_683),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_723),
.B(n_631),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_756),
.B(n_683),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_766),
.Y(n_776)
);

O2A1O1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_732),
.A2(n_564),
.B(n_566),
.C(n_530),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_738),
.B(n_682),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_745),
.A2(n_664),
.B(n_635),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_732),
.A2(n_641),
.B1(n_633),
.B2(n_445),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_759),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_709),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_712),
.B(n_682),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_714),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_752),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_711),
.B(n_664),
.Y(n_786)
);

OAI21xp33_ASAP7_75t_L g787 ( 
.A1(n_723),
.A2(n_613),
.B(n_592),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_720),
.A2(n_667),
.B(n_478),
.Y(n_788)
);

AOI21x1_ASAP7_75t_L g789 ( 
.A1(n_761),
.A2(n_764),
.B(n_748),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_739),
.A2(n_449),
.B(n_453),
.C(n_438),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_727),
.B(n_615),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_755),
.A2(n_734),
.B(n_752),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_711),
.A2(n_479),
.B1(n_459),
.B2(n_391),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_728),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_728),
.B(n_715),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_730),
.B(n_468),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_724),
.A2(n_573),
.B(n_624),
.C(n_616),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_758),
.B(n_389),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_733),
.A2(n_718),
.B1(n_743),
.B2(n_726),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_725),
.A2(n_667),
.B(n_656),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_749),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_741),
.B(n_480),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_770),
.B(n_656),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_735),
.A2(n_667),
.B(n_681),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_747),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_717),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_765),
.A2(n_400),
.B(n_398),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_758),
.B(n_630),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_750),
.B(n_487),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_747),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_769),
.B(n_449),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_721),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_740),
.B(n_637),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_747),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_762),
.B(n_399),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_736),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_751),
.B(n_513),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_744),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_768),
.A2(n_413),
.B(n_412),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_762),
.B(n_651),
.C(n_639),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_719),
.B(n_516),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_746),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_722),
.B(n_482),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_754),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_760),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_729),
.B(n_517),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_767),
.A2(n_420),
.B(n_417),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_742),
.A2(n_430),
.B(n_427),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_757),
.B(n_521),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_707),
.B(n_525),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_737),
.B(n_484),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_708),
.A2(n_716),
.B(n_737),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_760),
.B(n_644),
.Y(n_833)
);

AOI21xp33_ASAP7_75t_L g834 ( 
.A1(n_760),
.A2(n_528),
.B(n_526),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_753),
.A2(n_434),
.B(n_433),
.Y(n_835)
);

INVx4_ASAP7_75t_L g836 ( 
.A(n_753),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_709),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_710),
.A2(n_452),
.B(n_436),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_731),
.B(n_532),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_710),
.A2(n_466),
.B(n_461),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_763),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_738),
.B(n_484),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_710),
.A2(n_475),
.B(n_467),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_713),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_709),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_709),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_766),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_738),
.B(n_496),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_763),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_731),
.B(n_537),
.Y(n_850)
);

O2A1O1Ixp5_ASAP7_75t_L g851 ( 
.A1(n_731),
.A2(n_496),
.B(n_490),
.C(n_492),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_710),
.A2(n_495),
.B(n_489),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_731),
.B(n_543),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_709),
.Y(n_854)
);

NOR2xp67_ASAP7_75t_L g855 ( 
.A(n_743),
.B(n_401),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_709),
.B(n_644),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_710),
.A2(n_503),
.B(n_501),
.Y(n_857)
);

OAI321xp33_ASAP7_75t_L g858 ( 
.A1(n_732),
.A2(n_524),
.A3(n_511),
.B1(n_527),
.B2(n_519),
.C(n_508),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_731),
.B(n_544),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_713),
.B(n_652),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_731),
.B(n_545),
.Y(n_861)
);

BUFx4f_ASAP7_75t_L g862 ( 
.A(n_760),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_763),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_710),
.A2(n_531),
.B(n_529),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_732),
.A2(n_641),
.B1(n_533),
.B2(n_536),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_738),
.B(n_551),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_710),
.A2(n_560),
.B(n_558),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_710),
.A2(n_574),
.B(n_565),
.Y(n_868)
);

AND2x2_ASAP7_75t_SL g869 ( 
.A(n_743),
.B(n_578),
.Y(n_869)
);

NOR2xp67_ASAP7_75t_L g870 ( 
.A(n_743),
.B(n_403),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_710),
.A2(n_429),
.B(n_405),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_723),
.B(n_642),
.C(n_559),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_789),
.A2(n_606),
.B(n_600),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_792),
.A2(n_641),
.B(n_450),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_781),
.B(n_670),
.Y(n_875)
);

AO21x1_ASAP7_75t_L g876 ( 
.A1(n_777),
.A2(n_848),
.B(n_842),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_839),
.B(n_439),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_850),
.B(n_455),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_784),
.B(n_782),
.Y(n_879)
);

BUFx12f_ASAP7_75t_L g880 ( 
.A(n_836),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_860),
.B(n_670),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_844),
.B(n_684),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_853),
.B(n_463),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_805),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_784),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_795),
.A2(n_465),
.B1(n_471),
.B2(n_464),
.Y(n_886)
);

AOI21xp33_ASAP7_75t_L g887 ( 
.A1(n_802),
.A2(n_476),
.B(n_474),
.Y(n_887)
);

OAI21x1_ASAP7_75t_L g888 ( 
.A1(n_832),
.A2(n_628),
.B(n_627),
.Y(n_888)
);

O2A1O1Ixp5_ASAP7_75t_L g889 ( 
.A1(n_772),
.A2(n_629),
.B(n_632),
.C(n_628),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_771),
.A2(n_483),
.B(n_477),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_865),
.A2(n_486),
.B1(n_493),
.B2(n_485),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_785),
.B(n_684),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_779),
.A2(n_498),
.B(n_494),
.Y(n_893)
);

AO31x2_ASAP7_75t_L g894 ( 
.A1(n_866),
.A2(n_632),
.A3(n_638),
.B(n_629),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_813),
.B(n_603),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_784),
.Y(n_896)
);

OAI21xp33_ASAP7_75t_L g897 ( 
.A1(n_809),
.A2(n_640),
.B(n_638),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_776),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_859),
.A2(n_504),
.B(n_505),
.C(n_500),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_861),
.B(n_507),
.Y(n_900)
);

NOR2xp67_ASAP7_75t_SL g901 ( 
.A(n_858),
.B(n_510),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_800),
.A2(n_788),
.B(n_804),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_808),
.B(n_512),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_778),
.A2(n_803),
.B(n_783),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_841),
.B(n_518),
.Y(n_905)
);

AO31x2_ASAP7_75t_L g906 ( 
.A1(n_811),
.A2(n_25),
.A3(n_23),
.B(n_24),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_849),
.B(n_522),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_863),
.B(n_535),
.Y(n_908)
);

OAI21x1_ASAP7_75t_SL g909 ( 
.A1(n_827),
.A2(n_131),
.B(n_129),
.Y(n_909)
);

OA22x2_ASAP7_75t_L g910 ( 
.A1(n_810),
.A2(n_546),
.B1(n_553),
.B2(n_542),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_801),
.B(n_554),
.Y(n_911)
);

OAI21x1_ASAP7_75t_L g912 ( 
.A1(n_831),
.A2(n_133),
.B(n_132),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_847),
.B(n_556),
.Y(n_913)
);

AO21x2_ASAP7_75t_L g914 ( 
.A1(n_786),
.A2(n_136),
.B(n_135),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_780),
.A2(n_571),
.B(n_557),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_791),
.B(n_572),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_782),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_851),
.A2(n_138),
.B(n_137),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_812),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_782),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_796),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_799),
.A2(n_144),
.B(n_142),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_837),
.Y(n_923)
);

AO31x2_ASAP7_75t_L g924 ( 
.A1(n_838),
.A2(n_30),
.A3(n_26),
.B(n_29),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_794),
.A2(n_146),
.B1(n_147),
.B2(n_145),
.Y(n_925)
);

AOI21x1_ASAP7_75t_SL g926 ( 
.A1(n_823),
.A2(n_29),
.B(n_30),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_822),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_856),
.B(n_791),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_793),
.A2(n_152),
.B1(n_154),
.B2(n_151),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_775),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_837),
.A2(n_156),
.B1(n_157),
.B2(n_155),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_840),
.A2(n_159),
.B(n_158),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_843),
.A2(n_162),
.B(n_160),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_852),
.A2(n_173),
.B(n_170),
.Y(n_934)
);

OAI21xp33_ASAP7_75t_L g935 ( 
.A1(n_787),
.A2(n_31),
.B(n_32),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_856),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_819),
.A2(n_176),
.B(n_175),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_833),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_836),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_837),
.A2(n_179),
.B1(n_180),
.B2(n_178),
.Y(n_940)
);

OAI21xp33_ASAP7_75t_L g941 ( 
.A1(n_774),
.A2(n_32),
.B(n_34),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_846),
.A2(n_182),
.B1(n_183),
.B2(n_181),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_857),
.B(n_34),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_816),
.A2(n_185),
.B(n_184),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_864),
.B(n_35),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_824),
.A2(n_189),
.B(n_186),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_867),
.B(n_35),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_868),
.B(n_36),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_806),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_871),
.A2(n_191),
.B(n_190),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_846),
.Y(n_951)
);

AO21x2_ASAP7_75t_L g952 ( 
.A1(n_798),
.A2(n_194),
.B(n_193),
.Y(n_952)
);

AO31x2_ASAP7_75t_L g953 ( 
.A1(n_807),
.A2(n_39),
.A3(n_37),
.B(n_38),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_854),
.B(n_845),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_854),
.B(n_38),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_814),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_812),
.A2(n_197),
.B(n_195),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_854),
.B(n_39),
.Y(n_958)
);

AOI221xp5_ASAP7_75t_L g959 ( 
.A1(n_797),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.C(n_44),
.Y(n_959)
);

NAND2x1_ASAP7_75t_L g960 ( 
.A(n_812),
.B(n_198),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_818),
.A2(n_200),
.B(n_199),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_773),
.B(n_40),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_855),
.B(n_201),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_817),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_964)
);

AO21x2_ASAP7_75t_L g965 ( 
.A1(n_870),
.A2(n_204),
.B(n_203),
.Y(n_965)
);

OAI21xp33_ASAP7_75t_L g966 ( 
.A1(n_815),
.A2(n_45),
.B(n_46),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_862),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_821),
.B(n_45),
.Y(n_968)
);

AO31x2_ASAP7_75t_L g969 ( 
.A1(n_826),
.A2(n_49),
.A3(n_46),
.B(n_48),
.Y(n_969)
);

AO31x2_ASAP7_75t_L g970 ( 
.A1(n_830),
.A2(n_50),
.A3(n_48),
.B(n_49),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_820),
.B(n_51),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_818),
.B(n_53),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_872),
.A2(n_209),
.B(n_208),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_828),
.A2(n_835),
.B(n_829),
.Y(n_974)
);

NAND2x1p5_ASAP7_75t_L g975 ( 
.A(n_825),
.B(n_210),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_834),
.A2(n_383),
.B(n_212),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_869),
.B(n_53),
.Y(n_977)
);

AO31x2_ASAP7_75t_L g978 ( 
.A1(n_790),
.A2(n_56),
.A3(n_54),
.B(n_55),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_792),
.A2(n_213),
.B(n_211),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_784),
.B(n_214),
.Y(n_980)
);

AO32x2_ASAP7_75t_L g981 ( 
.A1(n_799),
.A2(n_55),
.A3(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_981)
);

NOR2xp67_ASAP7_75t_L g982 ( 
.A(n_872),
.B(n_216),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_799),
.A2(n_219),
.B1(n_222),
.B2(n_218),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_771),
.A2(n_224),
.B(n_223),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_792),
.A2(n_226),
.B(n_225),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_839),
.B(n_58),
.Y(n_986)
);

AO31x2_ASAP7_75t_L g987 ( 
.A1(n_790),
.A2(n_60),
.A3(n_61),
.B(n_62),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_784),
.B(n_227),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_839),
.B(n_60),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_844),
.Y(n_990)
);

OAI21x1_ASAP7_75t_SL g991 ( 
.A1(n_792),
.A2(n_229),
.B(n_228),
.Y(n_991)
);

AOI221xp5_ASAP7_75t_SL g992 ( 
.A1(n_777),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.C(n_66),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_792),
.A2(n_271),
.B1(n_381),
.B2(n_379),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_812),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_784),
.B(n_231),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_839),
.B(n_65),
.Y(n_996)
);

AO31x2_ASAP7_75t_L g997 ( 
.A1(n_790),
.A2(n_66),
.A3(n_67),
.B(n_68),
.Y(n_997)
);

BUFx12f_ASAP7_75t_L g998 ( 
.A(n_836),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_839),
.B(n_67),
.Y(n_999)
);

AO22x2_ASAP7_75t_L g1000 ( 
.A1(n_799),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_839),
.B(n_69),
.Y(n_1001)
);

OAI31xp33_ASAP7_75t_SL g1002 ( 
.A1(n_799),
.A2(n_70),
.A3(n_71),
.B(n_72),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_792),
.A2(n_279),
.B1(n_373),
.B2(n_372),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_771),
.A2(n_237),
.B(n_236),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_839),
.B(n_73),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_839),
.B(n_74),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_792),
.A2(n_239),
.B(n_238),
.Y(n_1007)
);

AND3x4_ASAP7_75t_L g1008 ( 
.A(n_820),
.B(n_75),
.C(n_76),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_860),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_839),
.B(n_76),
.Y(n_1010)
);

NOR2x1_ASAP7_75t_SL g1011 ( 
.A(n_771),
.B(n_241),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_SL g1012 ( 
.A1(n_792),
.A2(n_246),
.B(n_242),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_771),
.A2(n_250),
.B(n_249),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_839),
.B(n_77),
.Y(n_1014)
);

BUFx10_ASAP7_75t_L g1015 ( 
.A(n_829),
.Y(n_1015)
);

INVxp67_ASAP7_75t_SL g1016 ( 
.A(n_896),
.Y(n_1016)
);

AO21x1_ASAP7_75t_L g1017 ( 
.A1(n_986),
.A2(n_79),
.B(n_80),
.Y(n_1017)
);

NAND2x1p5_ASAP7_75t_L g1018 ( 
.A(n_896),
.B(n_259),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_895),
.B(n_79),
.Y(n_1019)
);

INVx3_ASAP7_75t_SL g1020 ( 
.A(n_967),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_888),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_919),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_904),
.A2(n_299),
.B(n_369),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_956),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_898),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_930),
.B(n_81),
.Y(n_1026)
);

NAND3xp33_ASAP7_75t_L g1027 ( 
.A(n_968),
.B(n_81),
.C(n_83),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_927),
.Y(n_1028)
);

OR2x6_ASAP7_75t_L g1029 ( 
.A(n_880),
.B(n_83),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_903),
.A2(n_296),
.B1(n_368),
.B2(n_365),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_884),
.Y(n_1031)
);

BUFx12f_ASAP7_75t_L g1032 ( 
.A(n_998),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_874),
.A2(n_290),
.B(n_363),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_989),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_1034)
);

AO21x2_ASAP7_75t_L g1035 ( 
.A1(n_876),
.A2(n_293),
.B(n_362),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_939),
.Y(n_1036)
);

AOI221xp5_ASAP7_75t_L g1037 ( 
.A1(n_941),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.C(n_89),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_938),
.B(n_262),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1009),
.B(n_88),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_928),
.B(n_877),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_893),
.A2(n_301),
.B(n_360),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_889),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_990),
.Y(n_1043)
);

CKINVDCx16_ASAP7_75t_R g1044 ( 
.A(n_875),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_916),
.B(n_90),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_954),
.B(n_90),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_936),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_999),
.A2(n_287),
.B1(n_358),
.B2(n_356),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1001),
.A2(n_283),
.B(n_355),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_1005),
.A2(n_91),
.B(n_92),
.C(n_93),
.Y(n_1050)
);

CKINVDCx11_ASAP7_75t_R g1051 ( 
.A(n_1015),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_1015),
.B(n_91),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1006),
.A2(n_282),
.B1(n_352),
.B2(n_351),
.Y(n_1053)
);

BUFx2_ASAP7_75t_SL g1054 ( 
.A(n_917),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_894),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_878),
.B(n_93),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_994),
.Y(n_1057)
);

AO21x1_ASAP7_75t_L g1058 ( 
.A1(n_1010),
.A2(n_1014),
.B(n_922),
.Y(n_1058)
);

BUFx4_ASAP7_75t_SL g1059 ( 
.A(n_951),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_881),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_917),
.B(n_266),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_917),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_949),
.B(n_882),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_894),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_892),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_883),
.A2(n_305),
.B1(n_349),
.B2(n_348),
.Y(n_1066)
);

CKINVDCx16_ASAP7_75t_R g1067 ( 
.A(n_920),
.Y(n_1067)
);

OR2x6_ASAP7_75t_L g1068 ( 
.A(n_920),
.B(n_95),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_900),
.A2(n_280),
.B1(n_341),
.B2(n_340),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_920),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_911),
.B(n_96),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_SL g1072 ( 
.A1(n_979),
.A2(n_275),
.B(n_338),
.C(n_337),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_885),
.B(n_96),
.Y(n_1073)
);

OA21x2_ASAP7_75t_L g1074 ( 
.A1(n_918),
.A2(n_274),
.B(n_336),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_SL g1075 ( 
.A1(n_901),
.A2(n_269),
.B(n_329),
.C(n_328),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_SL g1076 ( 
.A1(n_962),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_894),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_923),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_985),
.A2(n_1007),
.B(n_915),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_912),
.A2(n_268),
.B(n_324),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_971),
.B(n_98),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_978),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_955),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_978),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_978),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_879),
.B(n_101),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_972),
.Y(n_1087)
);

INVx4_ASAP7_75t_L g1088 ( 
.A(n_975),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_958),
.B(n_306),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_913),
.B(n_905),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_910),
.Y(n_1091)
);

BUFx10_ASAP7_75t_L g1092 ( 
.A(n_926),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_987),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_977),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_987),
.Y(n_1095)
);

BUFx12f_ASAP7_75t_L g1096 ( 
.A(n_1008),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_987),
.Y(n_1097)
);

NOR2xp67_ASAP7_75t_L g1098 ( 
.A(n_907),
.B(n_371),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_997),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_960),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_SL g1101 ( 
.A1(n_991),
.A2(n_322),
.B(n_321),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_908),
.B(n_101),
.Y(n_1102)
);

NAND2x1p5_ASAP7_75t_L g1103 ( 
.A(n_963),
.B(n_320),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_997),
.Y(n_1104)
);

BUFx12f_ASAP7_75t_L g1105 ( 
.A(n_982),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_983),
.A2(n_318),
.B1(n_317),
.B2(n_316),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_935),
.B(n_102),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_966),
.B(n_102),
.Y(n_1108)
);

OAI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_943),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_887),
.B(n_104),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_974),
.B(n_1011),
.Y(n_1111)
);

AOI21xp33_ASAP7_75t_L g1112 ( 
.A1(n_886),
.A2(n_108),
.B(n_109),
.Y(n_1112)
);

CKINVDCx11_ASAP7_75t_R g1113 ( 
.A(n_929),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_897),
.B(n_108),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_980),
.B(n_988),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_914),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_995),
.B(n_313),
.Y(n_1117)
);

INVx6_ASAP7_75t_L g1118 ( 
.A(n_1000),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_899),
.A2(n_308),
.B(n_307),
.Y(n_1119)
);

OA21x2_ASAP7_75t_L g1120 ( 
.A1(n_950),
.A2(n_110),
.B(n_111),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_976),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_SL g1122 ( 
.A1(n_909),
.A2(n_112),
.B(n_113),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_1000),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_945),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_1124)
);

AOI221xp5_ASAP7_75t_L g1125 ( 
.A1(n_959),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.C(n_118),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_952),
.B(n_116),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_947),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_948),
.Y(n_1128)
);

OAI222xp33_ASAP7_75t_L g1129 ( 
.A1(n_993),
.A2(n_1003),
.B1(n_1002),
.B2(n_925),
.C1(n_940),
.C2(n_942),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_891),
.B(n_921),
.Y(n_1130)
);

OA21x2_ASAP7_75t_L g1131 ( 
.A1(n_932),
.A2(n_933),
.B(n_934),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_981),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_964),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_984),
.A2(n_1013),
.B(n_1004),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_973),
.B(n_890),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_944),
.A2(n_946),
.B(n_937),
.C(n_961),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_992),
.B(n_970),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1012),
.A2(n_931),
.B(n_957),
.Y(n_1138)
);

OR2x6_ASAP7_75t_L g1139 ( 
.A(n_981),
.B(n_965),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_981),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_924),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_953),
.A2(n_906),
.B(n_970),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_969),
.A2(n_873),
.B(n_902),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_969),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_930),
.B(n_774),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_990),
.Y(n_1146)
);

BUFx5_ASAP7_75t_L g1147 ( 
.A(n_951),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_895),
.B(n_839),
.Y(n_1148)
);

AO21x1_ASAP7_75t_L g1149 ( 
.A1(n_986),
.A2(n_996),
.B(n_989),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_1146),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1022),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1094),
.B(n_1145),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1025),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_1031),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1044),
.B(n_1060),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1025),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1090),
.B(n_1040),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1125),
.A2(n_1037),
.B1(n_1112),
.B2(n_1133),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1081),
.B(n_1044),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_1079),
.A2(n_1058),
.B(n_1143),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1045),
.B(n_1102),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1148),
.B(n_1087),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1063),
.B(n_1043),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_1024),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1067),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1083),
.B(n_1026),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_1020),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1028),
.B(n_1108),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1067),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1057),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1047),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1065),
.B(n_1046),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1135),
.A2(n_1021),
.B(n_1042),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1091),
.B(n_1019),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1114),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1052),
.B(n_1068),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1062),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1100),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1107),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1100),
.Y(n_1180)
);

AO21x2_ASAP7_75t_L g1181 ( 
.A1(n_1149),
.A2(n_1137),
.B(n_1141),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1088),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_1071),
.B(n_1056),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1127),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1128),
.B(n_1140),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1039),
.Y(n_1186)
);

AO21x2_ASAP7_75t_L g1187 ( 
.A1(n_1141),
.A2(n_1055),
.B(n_1077),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1033),
.A2(n_1129),
.B(n_1041),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1073),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1068),
.B(n_1123),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1036),
.B(n_1070),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1082),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1147),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1082),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1147),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1084),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1105),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1084),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1085),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1147),
.Y(n_1200)
);

AOI211xp5_ASAP7_75t_L g1201 ( 
.A1(n_1109),
.A2(n_1110),
.B(n_1027),
.C(n_1017),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1097),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1059),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1113),
.A2(n_1034),
.B1(n_1124),
.B2(n_1076),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1078),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1089),
.B(n_1147),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1097),
.Y(n_1207)
);

BUFx8_ASAP7_75t_L g1208 ( 
.A(n_1032),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1054),
.B(n_1016),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1086),
.B(n_1096),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1051),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1089),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1131),
.A2(n_1134),
.B(n_1136),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1093),
.Y(n_1214)
);

AO21x2_ASAP7_75t_L g1215 ( 
.A1(n_1055),
.A2(n_1064),
.B(n_1077),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1118),
.A2(n_1139),
.B1(n_1132),
.B2(n_1130),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1118),
.B(n_1050),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1104),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1104),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1144),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1144),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1049),
.A2(n_1119),
.B(n_1072),
.C(n_1023),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1095),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1099),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1029),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1115),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1139),
.A2(n_1132),
.B1(n_1131),
.B2(n_1120),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1018),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1142),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1115),
.B(n_1117),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1080),
.A2(n_1138),
.B(n_1116),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1092),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1092),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1117),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1029),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1061),
.B(n_1098),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1126),
.B(n_1103),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1126),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1122),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1111),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1101),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1106),
.A2(n_1048),
.B1(n_1069),
.B2(n_1030),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1053),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1035),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1066),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1074),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1121),
.B(n_1075),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1038),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1024),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1145),
.B(n_774),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_1146),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1025),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1157),
.B(n_1179),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1157),
.B(n_1175),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1167),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1214),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1159),
.B(n_1161),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1163),
.B(n_1162),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1162),
.B(n_1152),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1164),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1168),
.B(n_1172),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1167),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1183),
.B(n_1191),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1185),
.B(n_1252),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1214),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1166),
.B(n_1250),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1250),
.B(n_1174),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1153),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1156),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1155),
.B(n_1217),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1155),
.B(n_1230),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1248),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1154),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1185),
.B(n_1150),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1230),
.B(n_1226),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1249),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1158),
.B(n_1226),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1169),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1165),
.B(n_1176),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1165),
.B(n_1210),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1223),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1251),
.B(n_1234),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1186),
.B(n_1189),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1248),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1212),
.B(n_1228),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1150),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1184),
.Y(n_1287)
);

INVxp67_ASAP7_75t_SL g1288 ( 
.A(n_1224),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1251),
.B(n_1204),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1238),
.B(n_1204),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1190),
.B(n_1171),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1158),
.B(n_1243),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1192),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1194),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1187),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1205),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1196),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1198),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1199),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1177),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1187),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1245),
.B(n_1188),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1209),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1188),
.B(n_1206),
.Y(n_1304)
);

INVx5_ASAP7_75t_SL g1305 ( 
.A(n_1197),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1202),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1197),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1215),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1215),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1206),
.B(n_1232),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1201),
.B(n_1233),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1228),
.B(n_1182),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1201),
.B(n_1237),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1235),
.B(n_1151),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1207),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1173),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1218),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1170),
.B(n_1216),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1216),
.B(n_1181),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1219),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1220),
.B(n_1221),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1236),
.B(n_1178),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1180),
.B(n_1197),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1180),
.B(n_1239),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1229),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1296),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1258),
.B(n_1259),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1293),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1304),
.B(n_1181),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1294),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1304),
.B(n_1227),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1297),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1315),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1298),
.B(n_1227),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1319),
.B(n_1160),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1299),
.B(n_1160),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1325),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1267),
.B(n_1225),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1266),
.B(n_1225),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1306),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1261),
.Y(n_1341)
);

NOR2x1p5_ASAP7_75t_L g1342 ( 
.A(n_1292),
.B(n_1211),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1317),
.B(n_1320),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1319),
.B(n_1213),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1275),
.B(n_1240),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1253),
.B(n_1213),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1253),
.B(n_1240),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1321),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1315),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1254),
.B(n_1241),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1313),
.B(n_1246),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1300),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1254),
.B(n_1193),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1281),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1289),
.B(n_1195),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1289),
.B(n_1200),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1286),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_1303),
.B(n_1211),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1283),
.B(n_1263),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1274),
.B(n_1244),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1271),
.B(n_1290),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1281),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1301),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1301),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1256),
.B(n_1265),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1268),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1270),
.B(n_1242),
.Y(n_1367)
);

BUFx2_ASAP7_75t_SL g1368 ( 
.A(n_1255),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1311),
.B(n_1247),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1288),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1324),
.B(n_1231),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1292),
.B(n_1242),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1286),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1269),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1264),
.B(n_1222),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1327),
.B(n_1303),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1345),
.B(n_1279),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1331),
.B(n_1308),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1337),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1345),
.B(n_1257),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1359),
.B(n_1302),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1337),
.Y(n_1382)
);

NOR2x1_ASAP7_75t_L g1383 ( 
.A(n_1368),
.B(n_1310),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1360),
.B(n_1277),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1370),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1333),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1331),
.B(n_1309),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1371),
.B(n_1309),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1357),
.B(n_1264),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1333),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1360),
.B(n_1277),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1343),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1354),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1373),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1329),
.B(n_1295),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1362),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1349),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1328),
.Y(n_1398)
);

NAND3xp33_ASAP7_75t_L g1399 ( 
.A(n_1372),
.B(n_1222),
.C(n_1282),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1369),
.B(n_1280),
.Y(n_1400)
);

AND2x2_ASAP7_75t_SL g1401 ( 
.A(n_1370),
.B(n_1318),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1369),
.B(n_1367),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1347),
.B(n_1287),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1330),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1344),
.B(n_1295),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1332),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1371),
.B(n_1288),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1329),
.B(n_1316),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1340),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1351),
.B(n_1291),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1351),
.B(n_1278),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1334),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1392),
.B(n_1334),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1395),
.B(n_1336),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1379),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1382),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1398),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1381),
.B(n_1346),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1402),
.B(n_1326),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1404),
.Y(n_1420)
);

INVxp33_ASAP7_75t_L g1421 ( 
.A(n_1402),
.Y(n_1421)
);

AOI211xp5_ASAP7_75t_SL g1422 ( 
.A1(n_1405),
.A2(n_1344),
.B(n_1335),
.C(n_1358),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1412),
.B(n_1335),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1395),
.B(n_1336),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1412),
.B(n_1363),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1408),
.B(n_1363),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1408),
.B(n_1364),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1378),
.B(n_1364),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1376),
.B(n_1341),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1385),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1380),
.B(n_1338),
.Y(n_1431)
);

AOI22x1_ASAP7_75t_SL g1432 ( 
.A1(n_1386),
.A2(n_1348),
.B1(n_1374),
.B2(n_1366),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1390),
.B(n_1365),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1389),
.B(n_1375),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1406),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1432),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1434),
.B(n_1394),
.Y(n_1437)
);

AOI21xp33_ASAP7_75t_L g1438 ( 
.A1(n_1421),
.A2(n_1399),
.B(n_1383),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1421),
.A2(n_1342),
.B1(n_1401),
.B2(n_1407),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1422),
.A2(n_1350),
.B(n_1356),
.C(n_1355),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1430),
.Y(n_1441)
);

NOR2x1p5_ASAP7_75t_SL g1442 ( 
.A(n_1423),
.B(n_1384),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1415),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1414),
.B(n_1401),
.Y(n_1444)
);

OAI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1418),
.A2(n_1361),
.B1(n_1391),
.B2(n_1394),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1419),
.B(n_1392),
.Y(n_1446)
);

NOR3xp33_ASAP7_75t_L g1447 ( 
.A(n_1429),
.B(n_1339),
.C(n_1262),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1431),
.A2(n_1407),
.B1(n_1400),
.B2(n_1388),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1414),
.B(n_1407),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1416),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1417),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1420),
.Y(n_1452)
);

AOI32xp33_ASAP7_75t_L g1453 ( 
.A1(n_1445),
.A2(n_1413),
.A3(n_1411),
.B1(n_1424),
.B2(n_1410),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1446),
.B(n_1423),
.Y(n_1454)
);

OAI21xp33_ASAP7_75t_L g1455 ( 
.A1(n_1442),
.A2(n_1403),
.B(n_1435),
.Y(n_1455)
);

AOI322xp5_ASAP7_75t_L g1456 ( 
.A1(n_1436),
.A2(n_1424),
.A3(n_1413),
.B1(n_1377),
.B2(n_1428),
.C1(n_1427),
.C2(n_1426),
.Y(n_1456)
);

OAI311xp33_ASAP7_75t_L g1457 ( 
.A1(n_1436),
.A2(n_1314),
.A3(n_1425),
.B1(n_1433),
.C1(n_1353),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1437),
.B(n_1438),
.Y(n_1458)
);

OAI21xp33_ASAP7_75t_L g1459 ( 
.A1(n_1440),
.A2(n_1397),
.B(n_1396),
.Y(n_1459)
);

AOI322xp5_ASAP7_75t_L g1460 ( 
.A1(n_1447),
.A2(n_1413),
.A3(n_1428),
.B1(n_1427),
.B2(n_1426),
.C1(n_1378),
.C2(n_1387),
.Y(n_1460)
);

NAND4xp25_ASAP7_75t_L g1461 ( 
.A(n_1459),
.B(n_1440),
.C(n_1439),
.D(n_1282),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1458),
.B(n_1441),
.Y(n_1462)
);

NAND4xp25_ASAP7_75t_L g1463 ( 
.A(n_1456),
.B(n_1453),
.C(n_1460),
.D(n_1455),
.Y(n_1463)
);

AOI211xp5_ASAP7_75t_L g1464 ( 
.A1(n_1457),
.A2(n_1452),
.B(n_1451),
.C(n_1448),
.Y(n_1464)
);

AOI221xp5_ASAP7_75t_L g1465 ( 
.A1(n_1454),
.A2(n_1450),
.B1(n_1443),
.B2(n_1444),
.C(n_1276),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1464),
.B(n_1449),
.Y(n_1466)
);

AOI211xp5_ASAP7_75t_L g1467 ( 
.A1(n_1463),
.A2(n_1307),
.B(n_1409),
.C(n_1393),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1462),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1465),
.B(n_1433),
.Y(n_1469)
);

NOR3xp33_ASAP7_75t_L g1470 ( 
.A(n_1461),
.B(n_1273),
.C(n_1322),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1462),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1468),
.B(n_1260),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1467),
.B(n_1260),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1470),
.B(n_1208),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1473),
.B(n_1471),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1472),
.Y(n_1476)
);

XOR2x1_ASAP7_75t_L g1477 ( 
.A(n_1475),
.B(n_1203),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1477),
.A2(n_1476),
.B1(n_1466),
.B2(n_1474),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1478),
.Y(n_1479)
);

NOR2xp67_ASAP7_75t_SL g1480 ( 
.A(n_1478),
.B(n_1208),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1479),
.A2(n_1469),
.B(n_1323),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1480),
.Y(n_1482)
);

AO21x2_ASAP7_75t_L g1483 ( 
.A1(n_1482),
.A2(n_1305),
.B(n_1323),
.Y(n_1483)
);

XOR2x1_ASAP7_75t_L g1484 ( 
.A(n_1481),
.B(n_1305),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1483),
.A2(n_1481),
.B1(n_1484),
.B2(n_1305),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1485),
.A2(n_1285),
.B(n_1312),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1486),
.B(n_1300),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1487),
.A2(n_1352),
.B1(n_1272),
.B2(n_1284),
.Y(n_1488)
);


endmodule