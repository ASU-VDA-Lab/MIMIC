module real_aes_8985_n_12 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10, n_11, n_12);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
input n_10;
input n_11;
output n_12;
wire n_28;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_19;
wire n_25;
wire n_14;
wire n_16;
wire n_15;
wire n_27;
wire n_23;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
NOR2xp33_ASAP7_75t_R g27 ( .A(n_0), .B(n_28), .Y(n_27) );
NAND2xp33_ASAP7_75t_SL g16 ( .A(n_1), .B(n_17), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_2), .Y(n_22) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_3), .B(n_7), .C(n_21), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_4), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_5), .Y(n_21) );
AOI22xp5_ASAP7_75t_SL g12 ( .A1(n_6), .A2(n_8), .B1(n_13), .B2(n_29), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g25 ( .A(n_9), .Y(n_25) );
CKINVDCx20_ASAP7_75t_R g28 ( .A(n_10), .Y(n_28) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_11), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_14), .Y(n_13) );
CKINVDCx16_ASAP7_75t_R g14 ( .A(n_15), .Y(n_14) );
INVx1_ASAP7_75t_SL g29 ( .A(n_15), .Y(n_29) );
NOR2xp33_ASAP7_75t_R g15 ( .A(n_16), .B(n_18), .Y(n_15) );
NAND2xp33_ASAP7_75t_SL g18 ( .A(n_19), .B(n_23), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_20), .B(n_22), .Y(n_19) );
NOR3xp33_ASAP7_75t_SL g23 ( .A(n_24), .B(n_25), .C(n_26), .Y(n_23) );
CKINVDCx16_ASAP7_75t_R g26 ( .A(n_27), .Y(n_26) );
endmodule