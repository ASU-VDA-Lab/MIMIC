module fake_jpeg_26344_n_227 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_25),
.Y(n_47)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_53),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_30),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_63),
.B(n_33),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_58),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_34),
.B1(n_27),
.B2(n_30),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_34),
.B1(n_27),
.B2(n_32),
.Y(n_67)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_28),
.Y(n_68)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_30),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_50),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_44),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_72),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_34),
.B1(n_26),
.B2(n_25),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_26),
.B1(n_42),
.B2(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_74),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_25),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_65),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_87),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_21),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_25),
.C(n_21),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_88),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_21),
.B1(n_28),
.B2(n_18),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_24),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_24),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_56),
.B(n_22),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_19),
.B(n_33),
.C(n_17),
.Y(n_88)
);

AOI22x1_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_28),
.B1(n_19),
.B2(n_33),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_89),
.A2(n_90),
.B1(n_87),
.B2(n_19),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_23),
.B1(n_18),
.B2(n_29),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_50),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_103),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_74),
.A2(n_61),
.B1(n_48),
.B2(n_58),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_75),
.B1(n_78),
.B2(n_61),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_108),
.Y(n_133)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_71),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_59),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_111),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_108),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_122),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_73),
.B1(n_78),
.B2(n_89),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_121),
.B1(n_104),
.B2(n_97),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_79),
.C(n_81),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_120),
.C(n_103),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_83),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_88),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_23),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_88),
.B(n_77),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_93),
.B(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_84),
.Y(n_141)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_52),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_75),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_137),
.B(n_29),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_79),
.B1(n_62),
.B2(n_52),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_136),
.A2(n_112),
.B1(n_106),
.B2(n_96),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_67),
.B(n_84),
.Y(n_137)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_113),
.B(n_98),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_143),
.B(n_149),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_99),
.B1(n_92),
.B2(n_95),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_144),
.B1(n_148),
.B2(n_158),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_135),
.B(n_125),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_146),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_97),
.B(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_147),
.B(n_134),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_102),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_102),
.C(n_96),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_120),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_153),
.B(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_156),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_86),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_0),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_159),
.Y(n_162)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_158),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_163),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_132),
.Y(n_163)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_170),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_126),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_149),
.B(n_117),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_148),
.A3(n_151),
.B1(n_155),
.B2(n_153),
.C1(n_149),
.C2(n_143),
.Y(n_174)
);

OAI21x1_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_15),
.B(n_13),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_177),
.C(n_5),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_124),
.B(n_117),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_176),
.A2(n_124),
.B1(n_145),
.B2(n_147),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_128),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_144),
.B1(n_157),
.B2(n_134),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_178),
.Y(n_193)
);

OAI321xp33_ASAP7_75t_L g180 ( 
.A1(n_176),
.A2(n_138),
.A3(n_145),
.B1(n_152),
.B2(n_157),
.C(n_150),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_171),
.A2(n_131),
.B1(n_136),
.B2(n_127),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_171),
.A2(n_127),
.B1(n_29),
.B2(n_17),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_187),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_185),
.A2(n_189),
.B(n_190),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_0),
.A3(n_1),
.B1(n_3),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_3),
.B(n_5),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_173),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_186),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_198),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_177),
.C(n_175),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_196),
.C(n_199),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_168),
.C(n_170),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_168),
.C(n_162),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_190),
.C(n_179),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_183),
.B1(n_184),
.B2(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_208),
.B1(n_200),
.B2(n_160),
.Y(n_213)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_204),
.Y(n_214)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_207),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_179),
.C(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_199),
.Y(n_208)
);

OAI221xp5_ASAP7_75t_L g212 ( 
.A1(n_209),
.A2(n_161),
.B1(n_181),
.B2(n_178),
.C(n_196),
.Y(n_212)
);

AOI31xp67_ASAP7_75t_SL g211 ( 
.A1(n_206),
.A2(n_194),
.A3(n_161),
.B(n_181),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_211),
.B(n_213),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

NOR2xp67_ASAP7_75t_SL g215 ( 
.A(n_206),
.B(n_6),
.Y(n_215)
);

AOI21x1_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_9),
.B(n_10),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_6),
.C(n_8),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_217),
.B(n_219),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_218),
.A2(n_216),
.B1(n_214),
.B2(n_11),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_9),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_10),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_221),
.C(n_220),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_223),
.B(n_10),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_12),
.Y(n_227)
);


endmodule