module fake_jpeg_8166_n_225 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_42),
.Y(n_55)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_23),
.B1(n_27),
.B2(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_45),
.B1(n_63),
.B2(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_20),
.B1(n_16),
.B2(n_19),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_41),
.B1(n_42),
.B2(n_40),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_26),
.B1(n_31),
.B2(n_21),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_58),
.B1(n_25),
.B2(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_56),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_21),
.B1(n_29),
.B2(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_26),
.B1(n_31),
.B2(n_29),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_16),
.B1(n_19),
.B2(n_24),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_42),
.C(n_33),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_80),
.Y(n_104)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_70),
.B1(n_76),
.B2(n_79),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_40),
.B1(n_38),
.B2(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_82),
.Y(n_89)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_83),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_43),
.B1(n_49),
.B2(n_59),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_33),
.B(n_22),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_22),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_53),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_1),
.B(n_2),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

OA21x2_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_50),
.B(n_32),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_67),
.B(n_80),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_66),
.B1(n_15),
.B2(n_28),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_96),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_61),
.B1(n_52),
.B2(n_46),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_105),
.B1(n_61),
.B2(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_61),
.B1(n_50),
.B2(n_62),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_107),
.B1(n_115),
.B2(n_99),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_95),
.B1(n_98),
.B2(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_114),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_30),
.B(n_4),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_73),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_71),
.B1(n_68),
.B2(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_118),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_124),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_28),
.C(n_15),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_126),
.C(n_25),
.Y(n_141)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_28),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_97),
.B1(n_103),
.B2(n_90),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_135),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_SL g130 ( 
.A(n_126),
.B(n_109),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_120),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_143),
.B1(n_125),
.B2(n_113),
.Y(n_151)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_146),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_89),
.B(n_90),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_138),
.B(n_139),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_144),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_93),
.B1(n_101),
.B2(n_15),
.Y(n_137)
);

AOI221xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_111),
.B1(n_30),
.B2(n_5),
.C(n_6),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_15),
.B1(n_25),
.B2(n_18),
.Y(n_138)
);

NOR2xp67_ASAP7_75t_R g139 ( 
.A(n_113),
.B(n_93),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_30),
.C(n_6),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_25),
.B1(n_30),
.B2(n_13),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_145),
.A2(n_3),
.B(n_4),
.Y(n_160)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_128),
.B1(n_131),
.B2(n_142),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_154),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_134),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_151),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_124),
.B1(n_115),
.B2(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_108),
.B1(n_117),
.B2(n_122),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_158),
.B(n_160),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_30),
.B1(n_12),
.B2(n_5),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_163),
.C(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_162),
.B(n_164),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_3),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

OA21x2_ASAP7_75t_SL g165 ( 
.A1(n_163),
.A2(n_139),
.B(n_129),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_167),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_173),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_174),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_145),
.C(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_143),
.C(n_138),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_3),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_7),
.Y(n_176)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_9),
.C(n_10),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_177),
.Y(n_181)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_186),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_155),
.B(n_159),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_183),
.A2(n_9),
.B(n_10),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_157),
.B(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_170),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_166),
.A2(n_154),
.B1(n_151),
.B2(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_161),
.B1(n_10),
.B2(n_11),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_191),
.B(n_175),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_169),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_195),
.C(n_198),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_168),
.C(n_181),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_185),
.A2(n_175),
.B(n_177),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_200),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_176),
.C(n_174),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

OAI221xp5_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_183),
.B1(n_190),
.B2(n_189),
.C(n_184),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_204),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_197),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_208),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_192),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_200),
.C(n_193),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_198),
.B(n_182),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_212),
.A2(n_190),
.B(n_207),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_216),
.A2(n_214),
.B(n_213),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_190),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_217),
.B(n_213),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_218),
.C(n_9),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_11),
.C(n_223),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_224),
.Y(n_225)
);


endmodule