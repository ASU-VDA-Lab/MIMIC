module fake_jpeg_11239_n_105 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_105);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_52),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_36),
.B1(n_38),
.B2(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_1),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_54),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_3),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_54),
.A2(n_45),
.B1(n_36),
.B2(n_46),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_41),
.B1(n_8),
.B2(n_7),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_64),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_66),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_4),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_5),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_7),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_14),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_41),
.B1(n_8),
.B2(n_12),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_10),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_79),
.C(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_13),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_15),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_85),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_26),
.C(n_27),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_28),
.B(n_29),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_88),
.B(n_89),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_34),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_84),
.Y(n_92)
);

NAND2xp67_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

OAI21x1_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_81),
.B(n_90),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_74),
.Y(n_98)
);

NAND2xp67_ASAP7_75t_SL g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

OAI21x1_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_93),
.B(n_98),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_94),
.B(n_88),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_94),
.B(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_35),
.Y(n_105)
);


endmodule