module fake_jpeg_31369_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

AOI21xp33_ASAP7_75t_L g8 ( 
.A1(n_6),
.A2(n_4),
.B(n_1),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx8_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_1),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx4_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_21),
.Y(n_26)
);

CKINVDCx12_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_15),
.B(n_2),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

AO22x1_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_13),
.B1(n_9),
.B2(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_27),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_17),
.B1(n_16),
.B2(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_11),
.Y(n_27)
);

AND2x6_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_16),
.Y(n_28)
);

NOR2xp67_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_13),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_19),
.B1(n_22),
.B2(n_3),
.Y(n_35)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_24),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_35),
.B(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_26),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_47),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_35),
.B(n_40),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_31),
.C(n_3),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_51),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_5),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_46),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

AO21x1_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_50),
.B(n_45),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_54),
.C(n_55),
.Y(n_57)
);

INVxp67_ASAP7_75t_SL g58 ( 
.A(n_57),
.Y(n_58)
);


endmodule