module fake_ariane_1041_n_1718 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_345, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_361, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_1718);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_345;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_1718;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_1716;
wire n_380;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_436;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1674;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_1687;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_1686;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_933;
wire n_954;
wire n_596;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_1569;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_234),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_39),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_356),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_317),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_43),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_260),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_81),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_115),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_39),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_60),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_92),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_138),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_142),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_190),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_319),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_122),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_318),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_341),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_264),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_74),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_199),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_210),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_312),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_240),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_307),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_29),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_172),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_177),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_337),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_211),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_116),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_88),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_129),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_182),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_227),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_56),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_78),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_220),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_82),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_214),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_108),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_32),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_225),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_57),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_203),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_137),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_344),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_163),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_198),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_313),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_186),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_269),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_311),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_102),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_327),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_156),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_322),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_324),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_332),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_237),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_286),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_36),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_348),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_126),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_152),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_338),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_94),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_347),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_105),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_183),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_72),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_263),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_49),
.Y(n_438)
);

BUFx10_ASAP7_75t_L g439 ( 
.A(n_25),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_147),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_253),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_79),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_330),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_59),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_325),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_169),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_70),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_8),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_185),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_131),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_320),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_65),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_294),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_53),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_146),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_34),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_204),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_34),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_148),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_21),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_331),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_48),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_140),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_46),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_101),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_329),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_154),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_241),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_47),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_46),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_14),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_106),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_21),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_215),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_16),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_113),
.Y(n_476)
);

BUFx10_ASAP7_75t_L g477 ( 
.A(n_361),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_135),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_328),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_144),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_358),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_68),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_45),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_13),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_251),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_255),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_64),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_302),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_168),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_28),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_268),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_143),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_239),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_292),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_90),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_301),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_179),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_273),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_83),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_54),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_128),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_162),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_123),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_224),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_316),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_343),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_35),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_150),
.Y(n_508)
);

BUFx5_ASAP7_75t_L g509 ( 
.A(n_118),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_17),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_221),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_226),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_261),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_175),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_25),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_18),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_336),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_259),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_271),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_306),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_194),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_287),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_288),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_355),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_29),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_132),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_62),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_173),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_293),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_171),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_334),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_195),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_280),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_352),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_26),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_242),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_201),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_161),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_321),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_340),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_184),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_3),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_73),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_174),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_1),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_206),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_134),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_89),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_258),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_97),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_323),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_266),
.Y(n_552)
);

BUFx10_ASAP7_75t_L g553 ( 
.A(n_23),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_354),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_244),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_3),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_55),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_256),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_110),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_217),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_357),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_229),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_10),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_136),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_9),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_291),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_196),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_188),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_180),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_187),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_333),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_170),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_84),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_149),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_11),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_32),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_309),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_277),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_339),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_335),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_103),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_202),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_326),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_30),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_117),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_125),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_235),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_120),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_26),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_213),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_95),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_218),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_290),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_315),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_314),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_236),
.Y(n_596)
);

BUFx10_ASAP7_75t_L g597 ( 
.A(n_299),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_274),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_228),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_363),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_310),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_104),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_484),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_495),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_495),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_386),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_391),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_448),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_427),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_460),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_367),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_462),
.Y(n_612)
);

INVxp33_ASAP7_75t_SL g613 ( 
.A(n_370),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_374),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_412),
.Y(n_615)
);

CKINVDCx16_ASAP7_75t_R g616 ( 
.A(n_434),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_452),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_464),
.B(n_0),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_543),
.B(n_0),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_472),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_489),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_508),
.Y(n_622)
);

INVxp33_ASAP7_75t_L g623 ( 
.A(n_475),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_519),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_526),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_537),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_507),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_544),
.Y(n_628)
);

CKINVDCx16_ASAP7_75t_R g629 ( 
.A(n_444),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_510),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g631 ( 
.A(n_407),
.B(n_1),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_542),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_558),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_556),
.Y(n_634)
);

INVxp33_ASAP7_75t_SL g635 ( 
.A(n_456),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_585),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_576),
.B(n_2),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_484),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_586),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_484),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_591),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_484),
.Y(n_642)
);

INVxp33_ASAP7_75t_L g643 ( 
.A(n_563),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_563),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_563),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_563),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_413),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_413),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_477),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_387),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_377),
.B(n_378),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_595),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_600),
.Y(n_653)
);

INVxp67_ASAP7_75t_SL g654 ( 
.A(n_394),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_469),
.Y(n_655)
);

NOR2xp67_ASAP7_75t_L g656 ( 
.A(n_458),
.B(n_470),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_471),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_473),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_477),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_483),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_597),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_490),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_597),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_439),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_439),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_375),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_553),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_515),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_553),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_383),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_516),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_525),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_535),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_389),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_390),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_396),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_545),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_397),
.Y(n_678)
);

CKINVDCx16_ASAP7_75t_R g679 ( 
.A(n_375),
.Y(n_679)
);

INVxp67_ASAP7_75t_SL g680 ( 
.A(n_488),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_565),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_400),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_575),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_584),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_405),
.B(n_2),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_589),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_366),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_369),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_409),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_421),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_554),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_555),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_376),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_423),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_435),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_379),
.Y(n_696)
);

NOR2xp67_ASAP7_75t_L g697 ( 
.A(n_446),
.B(n_4),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_450),
.B(n_4),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_380),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_560),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_463),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_467),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_474),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_381),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_382),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_385),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_592),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_392),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_R g709 ( 
.A(n_393),
.B(n_50),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_395),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_480),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_398),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_399),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_481),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_485),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_401),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_402),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_486),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_494),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_403),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_404),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_406),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_499),
.B(n_5),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_410),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_414),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_509),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_416),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_509),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_509),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_501),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_417),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_418),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_502),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_518),
.B(n_5),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_521),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_531),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_532),
.B(n_6),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_372),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_419),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_420),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_533),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_509),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_534),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_373),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_538),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_422),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_424),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_388),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_509),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_546),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_425),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_426),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_547),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_509),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_577),
.B(n_6),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_582),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_428),
.Y(n_757)
);

CKINVDCx16_ASAP7_75t_R g758 ( 
.A(n_505),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_587),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_368),
.B(n_7),
.Y(n_760)
);

INVxp33_ASAP7_75t_SL g761 ( 
.A(n_430),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_431),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_594),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_603),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_603),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_645),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_644),
.B(n_602),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_607),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_645),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_683),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_609),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_610),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_638),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_650),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_640),
.Y(n_775)
);

OA21x2_ASAP7_75t_L g776 ( 
.A1(n_726),
.A2(n_415),
.B(n_411),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_651),
.B(n_487),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_758),
.B(n_371),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_627),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_738),
.B(n_408),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_642),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_651),
.B(n_536),
.Y(n_782)
);

AND2x6_ASAP7_75t_L g783 ( 
.A(n_760),
.B(n_505),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_630),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_SL g785 ( 
.A(n_619),
.B(n_561),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_744),
.B(n_443),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_726),
.A2(n_729),
.B(n_728),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_646),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_632),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_634),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_748),
.B(n_493),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_670),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_674),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_655),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_675),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_728),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_650),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_679),
.B(n_548),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_676),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_729),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_742),
.Y(n_801)
);

OA21x2_ASAP7_75t_L g802 ( 
.A1(n_742),
.A2(n_442),
.B(n_429),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_749),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_647),
.B(n_482),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_678),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_749),
.Y(n_806)
);

BUFx8_ASAP7_75t_L g807 ( 
.A(n_611),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_754),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_682),
.B(n_568),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_689),
.B(n_384),
.Y(n_810)
);

BUFx8_ASAP7_75t_L g811 ( 
.A(n_658),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_700),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_690),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_648),
.B(n_514),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_754),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_616),
.A2(n_527),
.B1(n_599),
.B2(n_557),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_694),
.B(n_432),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_629),
.B(n_433),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_657),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_695),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_623),
.B(n_436),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_743),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_743),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_701),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_702),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_703),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_763),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_671),
.B(n_437),
.Y(n_828)
);

CKINVDCx16_ASAP7_75t_R g829 ( 
.A(n_666),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_613),
.A2(n_635),
.B1(n_710),
.B2(n_708),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_711),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_677),
.B(n_438),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_714),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_763),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_715),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_718),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_719),
.B(n_440),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_660),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_730),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_735),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_614),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_736),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_745),
.Y(n_843)
);

OA21x2_ASAP7_75t_L g844 ( 
.A1(n_685),
.A2(n_566),
.B(n_517),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_750),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_756),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_618),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_637),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_759),
.B(n_441),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_654),
.B(n_445),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_643),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_SL g852 ( 
.A(n_604),
.B(n_505),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_668),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_649),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_680),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_659),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_733),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_661),
.B(n_447),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_741),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_692),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_698),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_753),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_608),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_698),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_723),
.Y(n_865)
);

BUFx8_ASAP7_75t_L g866 ( 
.A(n_664),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_723),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_612),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_605),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_663),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_687),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_778),
.B(n_761),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_822),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_861),
.B(n_688),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_861),
.B(n_693),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_797),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_871),
.B(n_696),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_796),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_774),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_796),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_787),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_766),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_864),
.A2(n_861),
.B1(n_867),
.B2(n_865),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_768),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_766),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_780),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_786),
.Y(n_887)
);

AND2x2_ASAP7_75t_SL g888 ( 
.A(n_791),
.B(n_737),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_766),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_772),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_779),
.Y(n_891)
);

INVx1_ASAP7_75t_SL g892 ( 
.A(n_770),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_766),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_774),
.B(n_665),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_784),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_773),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_775),
.Y(n_897)
);

INVx5_ASAP7_75t_L g898 ( 
.A(n_783),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_789),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_797),
.B(n_667),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_790),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_822),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_843),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_822),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_822),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_794),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_812),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_871),
.B(n_699),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_843),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_778),
.B(n_704),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_823),
.B(n_669),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_843),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_781),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_855),
.B(n_705),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_843),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_823),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_808),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_861),
.B(n_706),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_794),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_850),
.B(n_717),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_831),
.Y(n_921)
);

INVx5_ASAP7_75t_L g922 ( 
.A(n_783),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_798),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_827),
.B(n_720),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_827),
.B(n_834),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_821),
.B(n_724),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_831),
.Y(n_927)
);

BUFx6f_ASAP7_75t_SL g928 ( 
.A(n_857),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_792),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_788),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_793),
.Y(n_931)
);

BUFx10_ASAP7_75t_L g932 ( 
.A(n_858),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_795),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_839),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_808),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_818),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_850),
.B(n_725),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_800),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_834),
.B(n_727),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_801),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_803),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_806),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_815),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_828),
.B(n_731),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_799),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_764),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_805),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_769),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_851),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_864),
.A2(n_755),
.B1(n_737),
.B2(n_734),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_765),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_840),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_860),
.B(n_691),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_813),
.Y(n_954)
);

BUFx10_ASAP7_75t_L g955 ( 
.A(n_858),
.Y(n_955)
);

AND2x2_ASAP7_75t_SL g956 ( 
.A(n_829),
.B(n_755),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_765),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_820),
.Y(n_958)
);

NAND2xp33_ASAP7_75t_L g959 ( 
.A(n_783),
.B(n_732),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_812),
.B(n_841),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_776),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_839),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_776),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_824),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_802),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_825),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_802),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_844),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_826),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_783),
.Y(n_970)
);

AO21x2_ASAP7_75t_L g971 ( 
.A1(n_817),
.A2(n_709),
.B(n_697),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_833),
.Y(n_972)
);

AO22x2_ASAP7_75t_L g973 ( 
.A1(n_923),
.A2(n_841),
.B1(n_869),
.B2(n_615),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_969),
.Y(n_974)
);

AO22x2_ASAP7_75t_L g975 ( 
.A1(n_886),
.A2(n_617),
.B1(n_621),
.B2(n_606),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_960),
.B(n_907),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_969),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_879),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_941),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_920),
.B(n_847),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_892),
.B(n_953),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_874),
.B(n_819),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_941),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_937),
.B(n_847),
.Y(n_984)
);

AO22x2_ASAP7_75t_L g985 ( 
.A1(n_887),
.A2(n_625),
.B1(n_628),
.B2(n_624),
.Y(n_985)
);

NAND2x1p5_ASAP7_75t_L g986 ( 
.A(n_953),
.B(n_936),
.Y(n_986)
);

NAND2x1p5_ASAP7_75t_L g987 ( 
.A(n_949),
.B(n_830),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_884),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_890),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_891),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_888),
.A2(n_782),
.B1(n_777),
.B2(n_819),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_883),
.B(n_847),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_895),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_872),
.B(n_910),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_899),
.Y(n_995)
);

AND2x6_ASAP7_75t_L g996 ( 
.A(n_963),
.B(n_847),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_917),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_901),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_929),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_906),
.Y(n_1000)
);

OAI221xp5_ASAP7_75t_L g1001 ( 
.A1(n_950),
.A2(n_777),
.B1(n_782),
.B2(n_816),
.C(n_810),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_875),
.B(n_838),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_918),
.B(n_848),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_931),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_911),
.B(n_639),
.Y(n_1005)
);

AO22x2_ASAP7_75t_L g1006 ( 
.A1(n_956),
.A2(n_652),
.B1(n_862),
.B2(n_859),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_917),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_917),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_933),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_945),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_914),
.A2(n_853),
.B1(n_838),
.B2(n_713),
.Y(n_1011)
);

AO22x2_ASAP7_75t_L g1012 ( 
.A1(n_964),
.A2(n_804),
.B1(n_814),
.B2(n_870),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_916),
.B(n_854),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_919),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_878),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_934),
.B(n_848),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_934),
.B(n_848),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_902),
.Y(n_1018)
);

AO22x2_ASAP7_75t_L g1019 ( 
.A1(n_966),
.A2(n_804),
.B1(n_814),
.B2(n_662),
.Y(n_1019)
);

NOR2xp67_ASAP7_75t_L g1020 ( 
.A(n_877),
.B(n_853),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_908),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_947),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_954),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_970),
.B(n_894),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_878),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_958),
.Y(n_1026)
);

NOR2xp67_ASAP7_75t_L g1027 ( 
.A(n_924),
.B(n_771),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_911),
.B(n_854),
.Y(n_1028)
);

OA22x2_ASAP7_75t_L g1029 ( 
.A1(n_894),
.A2(n_622),
.B1(n_626),
.B2(n_620),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_972),
.B(n_848),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_972),
.B(n_832),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_921),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_932),
.B(n_849),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_900),
.B(n_856),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_927),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_900),
.B(n_633),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_932),
.B(n_771),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_955),
.B(n_849),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_926),
.B(n_636),
.Y(n_1039)
);

NAND2x1p5_ASAP7_75t_L g1040 ( 
.A(n_970),
.B(n_856),
.Y(n_1040)
);

AO22x2_ASAP7_75t_L g1041 ( 
.A1(n_963),
.A2(n_809),
.B1(n_641),
.B2(n_653),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_928),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_938),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_955),
.B(n_863),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_940),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_898),
.B(n_868),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_952),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_876),
.B(n_809),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_944),
.B(n_672),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_880),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_880),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_942),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_962),
.B(n_707),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_943),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_SL g1055 ( 
.A(n_928),
.Y(n_1055)
);

AO22x2_ASAP7_75t_L g1056 ( 
.A1(n_896),
.A2(n_810),
.B1(n_836),
.B2(n_835),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_952),
.Y(n_1057)
);

AO22x2_ASAP7_75t_L g1058 ( 
.A1(n_897),
.A2(n_930),
.B1(n_913),
.B2(n_845),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_952),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_925),
.B(n_817),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_939),
.Y(n_1061)
);

BUFx8_ASAP7_75t_L g1062 ( 
.A(n_902),
.Y(n_1062)
);

NAND2x1p5_ASAP7_75t_L g1063 ( 
.A(n_898),
.B(n_922),
.Y(n_1063)
);

AO22x2_ASAP7_75t_L g1064 ( 
.A1(n_948),
.A2(n_846),
.B1(n_842),
.B2(n_811),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_935),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_873),
.B(n_712),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_951),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_971),
.B(n_673),
.Y(n_1068)
);

INVxp67_ASAP7_75t_L g1069 ( 
.A(n_873),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_912),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_957),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_959),
.A2(n_716),
.B1(n_722),
.B2(n_721),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_903),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_909),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_915),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_912),
.Y(n_1076)
);

BUFx8_ASAP7_75t_L g1077 ( 
.A(n_902),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_946),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_946),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_946),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_994),
.B(n_837),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_980),
.B(n_837),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_984),
.B(n_904),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_SL g1084 ( 
.A(n_1031),
.B(n_740),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_1011),
.B(n_904),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_991),
.B(n_904),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_976),
.B(n_905),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_1072),
.B(n_905),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_1061),
.B(n_905),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1048),
.B(n_767),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_1024),
.B(n_747),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1003),
.B(n_752),
.Y(n_1092)
);

NAND2xp33_ASAP7_75t_SL g1093 ( 
.A(n_1037),
.B(n_762),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1030),
.B(n_767),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_1027),
.B(n_739),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_1044),
.B(n_746),
.Y(n_1096)
);

NAND2xp33_ASAP7_75t_SL g1097 ( 
.A(n_1033),
.B(n_881),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1060),
.B(n_974),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_1028),
.B(n_751),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_1028),
.B(n_757),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1034),
.B(n_898),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_1014),
.B(n_684),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_1034),
.B(n_922),
.Y(n_1103)
);

NAND2xp33_ASAP7_75t_SL g1104 ( 
.A(n_1038),
.B(n_881),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_1068),
.B(n_922),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1036),
.B(n_686),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1020),
.B(n_881),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1013),
.B(n_992),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1013),
.B(n_807),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1016),
.B(n_807),
.Y(n_1110)
);

NAND2xp33_ASAP7_75t_SL g1111 ( 
.A(n_1017),
.B(n_709),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_1049),
.B(n_811),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_982),
.B(n_785),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_1002),
.B(n_785),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_978),
.B(n_882),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_987),
.B(n_1005),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_977),
.B(n_882),
.Y(n_1117)
);

NAND2xp33_ASAP7_75t_SL g1118 ( 
.A(n_1021),
.B(n_882),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_1066),
.B(n_885),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_1039),
.B(n_885),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_981),
.B(n_885),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_1047),
.B(n_893),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_1040),
.B(n_893),
.Y(n_1123)
);

NAND2xp33_ASAP7_75t_SL g1124 ( 
.A(n_988),
.B(n_893),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1056),
.B(n_783),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_989),
.B(n_866),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_990),
.B(n_866),
.Y(n_1127)
);

NAND2xp33_ASAP7_75t_SL g1128 ( 
.A(n_993),
.B(n_968),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_995),
.B(n_968),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_998),
.B(n_999),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1004),
.B(n_968),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_986),
.B(n_681),
.Y(n_1132)
);

NAND2xp33_ASAP7_75t_L g1133 ( 
.A(n_996),
.B(n_967),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_1022),
.B(n_1023),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1026),
.B(n_631),
.Y(n_1136)
);

NAND2xp33_ASAP7_75t_SL g1137 ( 
.A(n_1070),
.B(n_889),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1056),
.B(n_961),
.Y(n_1138)
);

NAND2xp33_ASAP7_75t_SL g1139 ( 
.A(n_1042),
.B(n_1059),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1057),
.B(n_961),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1018),
.B(n_961),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_1018),
.B(n_965),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1001),
.B(n_965),
.Y(n_1143)
);

NAND2xp33_ASAP7_75t_SL g1144 ( 
.A(n_1055),
.B(n_965),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1053),
.B(n_967),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1062),
.B(n_967),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1077),
.B(n_852),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1069),
.B(n_852),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_979),
.B(n_656),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_983),
.B(n_1032),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_1035),
.B(n_449),
.Y(n_1151)
);

NAND2xp33_ASAP7_75t_SL g1152 ( 
.A(n_1076),
.B(n_451),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1078),
.B(n_453),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1079),
.B(n_454),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1080),
.B(n_455),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1015),
.B(n_457),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1025),
.B(n_459),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1050),
.B(n_461),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1051),
.B(n_465),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_997),
.B(n_466),
.Y(n_1160)
);

NAND2xp33_ASAP7_75t_SL g1161 ( 
.A(n_1000),
.B(n_468),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1007),
.B(n_505),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1008),
.B(n_476),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_973),
.B(n_844),
.Y(n_1164)
);

NAND2xp33_ASAP7_75t_SL g1165 ( 
.A(n_1073),
.B(n_478),
.Y(n_1165)
);

NAND2xp33_ASAP7_75t_SL g1166 ( 
.A(n_1074),
.B(n_601),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1075),
.B(n_479),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1065),
.B(n_511),
.Y(n_1168)
);

NAND2xp33_ASAP7_75t_SL g1169 ( 
.A(n_1043),
.B(n_598),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_1138),
.A2(n_1071),
.A3(n_1067),
.B(n_1045),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1150),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1102),
.B(n_1052),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1098),
.A2(n_1054),
.B(n_1058),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_1132),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1130),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1081),
.A2(n_1046),
.B(n_1041),
.C(n_1006),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1146),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1082),
.A2(n_1058),
.B(n_1063),
.Y(n_1178)
);

AOI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1083),
.A2(n_1041),
.B(n_1012),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_1116),
.B(n_1006),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1134),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1090),
.B(n_1012),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1143),
.A2(n_1094),
.B1(n_1135),
.B2(n_1086),
.Y(n_1183)
);

AND3x4_ASAP7_75t_L g1184 ( 
.A(n_1093),
.B(n_1084),
.C(n_1106),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1149),
.A2(n_973),
.B1(n_1019),
.B2(n_1029),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1108),
.B(n_996),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1145),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_1118),
.Y(n_1188)
);

O2A1O1Ixp5_ASAP7_75t_L g1189 ( 
.A1(n_1097),
.A2(n_996),
.B(n_1064),
.C(n_1019),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1133),
.A2(n_492),
.B(n_491),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_1129),
.A2(n_497),
.B(n_496),
.Y(n_1191)
);

OAI21xp33_ASAP7_75t_L g1192 ( 
.A1(n_1151),
.A2(n_1064),
.B(n_985),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1085),
.B(n_975),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1104),
.A2(n_500),
.B(n_498),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1164),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1131),
.A2(n_52),
.B(n_51),
.Y(n_1196)
);

NOR2xp67_ASAP7_75t_L g1197 ( 
.A(n_1112),
.B(n_975),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1125),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1121),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1144),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1128),
.A2(n_985),
.A3(n_520),
.B(n_564),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1117),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1107),
.A2(n_504),
.B(n_503),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1092),
.B(n_7),
.Y(n_1204)
);

BUFx2_ASAP7_75t_SL g1205 ( 
.A(n_1109),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1088),
.B(n_8),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1139),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1119),
.Y(n_1208)
);

AO22x2_ASAP7_75t_L g1209 ( 
.A1(n_1126),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1141),
.A2(n_512),
.B(n_506),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1120),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1096),
.B(n_12),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1168),
.A2(n_520),
.A3(n_564),
.B(n_511),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1091),
.B(n_12),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1161),
.B(n_513),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1165),
.B(n_1166),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1142),
.A2(n_61),
.B(n_58),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1168),
.A2(n_66),
.B(n_63),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1127),
.B(n_13),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1140),
.A2(n_69),
.B(n_67),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1110),
.B(n_14),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1099),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1111),
.A2(n_523),
.B(n_522),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_SL g1224 ( 
.A1(n_1124),
.A2(n_15),
.B(n_16),
.Y(n_1224)
);

OA21x2_ASAP7_75t_L g1225 ( 
.A1(n_1162),
.A2(n_528),
.B(n_524),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1087),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1162),
.A2(n_75),
.B(n_71),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1105),
.A2(n_77),
.B(n_76),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1123),
.A2(n_530),
.B(n_529),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1136),
.A2(n_511),
.A3(n_564),
.B(n_520),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1113),
.B(n_15),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1122),
.A2(n_85),
.B(n_80),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1089),
.A2(n_540),
.B(n_539),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1167),
.A2(n_1115),
.B(n_1137),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1114),
.B(n_17),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1156),
.A2(n_549),
.B(n_541),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1100),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1148),
.Y(n_1238)
);

NAND3xp33_ASAP7_75t_L g1239 ( 
.A(n_1169),
.B(n_551),
.C(n_550),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1147),
.B(n_18),
.Y(n_1240)
);

OAI21xp33_ASAP7_75t_L g1241 ( 
.A1(n_1095),
.A2(n_559),
.B(n_552),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1157),
.A2(n_596),
.B1(n_593),
.B2(n_590),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1101),
.Y(n_1243)
);

AOI21xp33_ASAP7_75t_L g1244 ( 
.A1(n_1158),
.A2(n_567),
.B(n_562),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1183),
.A2(n_1154),
.B(n_1153),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1200),
.B(n_1103),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1172),
.B(n_1159),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1222),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1196),
.A2(n_1163),
.B(n_1160),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1217),
.A2(n_1155),
.B(n_1152),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1177),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1174),
.B(n_1188),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1220),
.A2(n_87),
.B(n_86),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1175),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1211),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1207),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1170),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1228),
.A2(n_93),
.B(n_91),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1238),
.A2(n_570),
.B(n_569),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1182),
.B(n_19),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1219),
.B(n_19),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1231),
.A2(n_572),
.B(n_571),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1176),
.A2(n_588),
.B(n_583),
.C(n_581),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1177),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_1177),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1243),
.B(n_96),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1199),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1181),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_SL g1269 ( 
.A1(n_1216),
.A2(n_1215),
.B(n_1235),
.C(n_1212),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1243),
.B(n_98),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1171),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1232),
.A2(n_100),
.B(n_99),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1218),
.A2(n_109),
.B(n_107),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1243),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1178),
.A2(n_574),
.B(n_573),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1192),
.A2(n_564),
.B1(n_520),
.B2(n_511),
.Y(n_1276)
);

AOI22x1_ASAP7_75t_L g1277 ( 
.A1(n_1234),
.A2(n_580),
.B1(n_579),
.B2(n_578),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1206),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1173),
.A2(n_112),
.B(n_111),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1170),
.Y(n_1280)
);

INVx6_ASAP7_75t_L g1281 ( 
.A(n_1184),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1223),
.A2(n_20),
.B(n_22),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1210),
.A2(n_233),
.B(n_364),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1237),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1170),
.Y(n_1285)
);

AO32x2_ASAP7_75t_L g1286 ( 
.A1(n_1185),
.A2(n_20),
.A3(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_1286)
);

AO21x2_ASAP7_75t_L g1287 ( 
.A1(n_1179),
.A2(n_238),
.B(n_362),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1189),
.A2(n_24),
.B(n_27),
.C(n_28),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1187),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1180),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1239),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1198),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1214),
.A2(n_1204),
.B(n_1244),
.C(n_1241),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1193),
.A2(n_246),
.A3(n_360),
.B(n_359),
.Y(n_1294)
);

NAND3xp33_ASAP7_75t_L g1295 ( 
.A(n_1203),
.B(n_33),
.C(n_36),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1208),
.B(n_114),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1195),
.B(n_365),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1205),
.Y(n_1298)
);

BUFx2_ASAP7_75t_SL g1299 ( 
.A(n_1240),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1226),
.B(n_119),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1221),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1242),
.B(n_37),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1186),
.A2(n_38),
.B(n_40),
.C(n_41),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1202),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1209),
.B(n_1197),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1230),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1209),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1191),
.A2(n_250),
.B(n_351),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1201),
.B(n_42),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_SL g1310 ( 
.A(n_1224),
.B(n_121),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1230),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1190),
.B(n_44),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1201),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1233),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1229),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1227),
.A2(n_252),
.B(n_350),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1236),
.B(n_44),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1233),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1230),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1191),
.A2(n_249),
.B(n_349),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1311),
.A2(n_1194),
.B(n_1213),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1254),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1292),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1280),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1255),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1285),
.Y(n_1326)
);

A2O1A1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1302),
.A2(n_1201),
.B(n_1225),
.C(n_48),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1257),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1300),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1304),
.B(n_1225),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1257),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1273),
.A2(n_1213),
.B(n_254),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1306),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1311),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1248),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1267),
.Y(n_1336)
);

AO21x2_ASAP7_75t_L g1337 ( 
.A1(n_1319),
.A2(n_1213),
.B(n_257),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1289),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1319),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1314),
.A2(n_1318),
.B(n_1309),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1278),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1268),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1286),
.B(n_45),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1271),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1313),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1292),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1294),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1260),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1297),
.B(n_124),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1300),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1286),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1305),
.A2(n_47),
.B1(n_127),
.B2(n_130),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1294),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1299),
.B(n_353),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1294),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1320),
.A2(n_133),
.B(n_139),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1286),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1274),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1275),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1252),
.Y(n_1360)
);

CKINVDCx8_ASAP7_75t_R g1361 ( 
.A(n_1256),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1279),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1274),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1307),
.B(n_141),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1274),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1297),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1247),
.B(n_346),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1264),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1251),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1287),
.Y(n_1370)
);

NOR2x1_ASAP7_75t_R g1371 ( 
.A(n_1281),
.B(n_145),
.Y(n_1371)
);

INVx11_ASAP7_75t_L g1372 ( 
.A(n_1281),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1275),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1261),
.B(n_151),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1266),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1316),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1284),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_1298),
.Y(n_1378)
);

OA21x2_ASAP7_75t_L g1379 ( 
.A1(n_1308),
.A2(n_153),
.B(n_155),
.Y(n_1379)
);

AO21x1_ASAP7_75t_SL g1380 ( 
.A1(n_1282),
.A2(n_157),
.B(n_158),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1253),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1266),
.Y(n_1382)
);

NAND2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1265),
.B(n_159),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1272),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1258),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1270),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1269),
.A2(n_345),
.B(n_164),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1270),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1301),
.B(n_160),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1295),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1265),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1350),
.B(n_1315),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1335),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1322),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_R g1395 ( 
.A(n_1377),
.B(n_1317),
.Y(n_1395)
);

INVxp67_ASAP7_75t_L g1396 ( 
.A(n_1360),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1335),
.B(n_1303),
.Y(n_1397)
);

CKINVDCx8_ASAP7_75t_R g1398 ( 
.A(n_1377),
.Y(n_1398)
);

XNOR2xp5_ASAP7_75t_L g1399 ( 
.A(n_1325),
.B(n_1290),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1341),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1361),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1350),
.B(n_1288),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1369),
.Y(n_1403)
);

XNOR2xp5_ASAP7_75t_L g1404 ( 
.A(n_1343),
.B(n_1246),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1363),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_1368),
.Y(n_1406)
);

INVxp67_ASAP7_75t_L g1407 ( 
.A(n_1358),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1350),
.B(n_1263),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1336),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1349),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1323),
.B(n_1296),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1382),
.B(n_1245),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1382),
.B(n_1366),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1346),
.B(n_1312),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1323),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1346),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1359),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1338),
.Y(n_1418)
);

OR2x6_ASAP7_75t_L g1419 ( 
.A(n_1349),
.B(n_1293),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1342),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1372),
.B(n_1262),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1348),
.B(n_1291),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1329),
.B(n_1249),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1329),
.B(n_1250),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1343),
.B(n_1259),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1361),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1365),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1374),
.B(n_1310),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_1367),
.Y(n_1429)
);

NAND2xp33_ASAP7_75t_R g1430 ( 
.A(n_1349),
.B(n_1283),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_R g1431 ( 
.A(n_1329),
.B(n_176),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1344),
.Y(n_1432)
);

XOR2xp5_ASAP7_75t_L g1433 ( 
.A(n_1354),
.B(n_1277),
.Y(n_1433)
);

XOR2xp5_ASAP7_75t_L g1434 ( 
.A(n_1354),
.B(n_1277),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1374),
.B(n_1330),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1351),
.B(n_1276),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1328),
.Y(n_1437)
);

INVxp67_ASAP7_75t_L g1438 ( 
.A(n_1367),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_R g1439 ( 
.A(n_1372),
.B(n_178),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1328),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1331),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1375),
.B(n_181),
.Y(n_1442)
);

OR2x6_ASAP7_75t_L g1443 ( 
.A(n_1383),
.B(n_189),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_R g1444 ( 
.A(n_1378),
.B(n_1391),
.Y(n_1444)
);

BUFx10_ASAP7_75t_L g1445 ( 
.A(n_1371),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1331),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1386),
.B(n_191),
.Y(n_1447)
);

NAND2xp33_ASAP7_75t_R g1448 ( 
.A(n_1340),
.B(n_192),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1388),
.B(n_1345),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1389),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1357),
.B(n_193),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1345),
.B(n_197),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1364),
.B(n_200),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1364),
.B(n_205),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1359),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1383),
.Y(n_1456)
);

NAND2xp33_ASAP7_75t_SL g1457 ( 
.A(n_1389),
.B(n_207),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1334),
.Y(n_1458)
);

OR2x6_ASAP7_75t_L g1459 ( 
.A(n_1387),
.B(n_208),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_R g1460 ( 
.A(n_1362),
.B(n_209),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1352),
.B(n_212),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1394),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1409),
.Y(n_1463)
);

AOI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1457),
.A2(n_1390),
.B1(n_1327),
.B2(n_1355),
.C(n_1353),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1435),
.B(n_1340),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1450),
.B(n_1327),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1400),
.B(n_1340),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1396),
.B(n_1334),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1418),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1420),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1393),
.B(n_1380),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1415),
.B(n_1380),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1428),
.B(n_1339),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1432),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1429),
.B(n_1373),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1456),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1433),
.A2(n_1362),
.B1(n_1356),
.B2(n_1379),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1433),
.A2(n_1362),
.B1(n_1356),
.B2(n_1379),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1416),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1437),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1405),
.B(n_1403),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1440),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1406),
.B(n_1339),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1458),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1414),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1455),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1427),
.B(n_1373),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1399),
.A2(n_1353),
.B1(n_1355),
.B2(n_1347),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1444),
.B(n_1347),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1438),
.B(n_1417),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1407),
.B(n_1324),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1441),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1446),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1425),
.A2(n_1410),
.B1(n_1454),
.B2(n_1395),
.Y(n_1494)
);

NAND2x1_ASAP7_75t_L g1495 ( 
.A(n_1419),
.B(n_1381),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1449),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1417),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1424),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1412),
.B(n_1321),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1443),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1422),
.B(n_1321),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1419),
.B(n_1321),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1404),
.B(n_1376),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1423),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1404),
.B(n_1324),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1436),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1426),
.B(n_1376),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1451),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1413),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1411),
.B(n_1385),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1392),
.B(n_1385),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1401),
.B(n_1384),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1452),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1397),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1434),
.B(n_1370),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1421),
.B(n_1384),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1399),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1498),
.B(n_1443),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1504),
.B(n_1402),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1504),
.B(n_1408),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1479),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1480),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1482),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1498),
.B(n_1381),
.Y(n_1524)
);

OAI31xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1466),
.A2(n_1461),
.A3(n_1430),
.B(n_1434),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1462),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1463),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1516),
.B(n_1453),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1490),
.B(n_1326),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1497),
.B(n_1370),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1502),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1470),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1486),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1474),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1469),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1486),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1484),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1490),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1510),
.B(n_1459),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1475),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1466),
.A2(n_1459),
.B1(n_1356),
.B2(n_1379),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1465),
.B(n_1333),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1494),
.A2(n_1398),
.B1(n_1447),
.B2(n_1442),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1492),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1475),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1500),
.A2(n_1448),
.B1(n_1445),
.B2(n_1337),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1468),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1485),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1503),
.B(n_1333),
.Y(n_1549)
);

INVx4_ASAP7_75t_L g1550 ( 
.A(n_1500),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1493),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1502),
.A2(n_1332),
.B(n_1326),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1467),
.B(n_1337),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1483),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1521),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1521),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1524),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1518),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1524),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1533),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1536),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1538),
.B(n_1481),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1530),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1538),
.B(n_1512),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1529),
.B(n_1540),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1543),
.B(n_1476),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1530),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1529),
.B(n_1501),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1522),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1518),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1520),
.B(n_1507),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1520),
.B(n_1511),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1519),
.B(n_1472),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1519),
.B(n_1489),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1522),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1531),
.B(n_1515),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1523),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1545),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1518),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1528),
.B(n_1554),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1527),
.Y(n_1581)
);

AO221x2_ASAP7_75t_L g1582 ( 
.A1(n_1566),
.A2(n_1517),
.B1(n_1525),
.B2(n_1526),
.C(n_1532),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1564),
.B(n_1528),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1564),
.B(n_1527),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1576),
.A2(n_1500),
.B1(n_1546),
.B2(n_1515),
.Y(n_1585)
);

OAI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1579),
.A2(n_1500),
.B1(n_1478),
.B2(n_1477),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1581),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1578),
.Y(n_1588)
);

NOR4xp25_ASAP7_75t_SL g1589 ( 
.A(n_1579),
.B(n_1508),
.C(n_1534),
.D(n_1548),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1576),
.B(n_1523),
.Y(n_1590)
);

NOR2x1_ASAP7_75t_L g1591 ( 
.A(n_1560),
.B(n_1550),
.Y(n_1591)
);

AOI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1574),
.A2(n_1514),
.B1(n_1539),
.B2(n_1494),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1561),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1571),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1574),
.A2(n_1539),
.B1(n_1541),
.B2(n_1471),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1561),
.Y(n_1596)
);

AO221x1_ASAP7_75t_L g1597 ( 
.A1(n_1558),
.A2(n_1547),
.B1(n_1537),
.B2(n_1535),
.C(n_1509),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1558),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1562),
.B(n_1537),
.Y(n_1599)
);

AO221x2_ASAP7_75t_L g1600 ( 
.A1(n_1557),
.A2(n_1550),
.B1(n_1501),
.B2(n_1513),
.C(n_1476),
.Y(n_1600)
);

INVxp33_ASAP7_75t_SL g1601 ( 
.A(n_1562),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_L g1602 ( 
.A(n_1558),
.B(n_1550),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1580),
.B(n_1473),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1583),
.B(n_1570),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1588),
.Y(n_1605)
);

NAND2xp33_ASAP7_75t_L g1606 ( 
.A(n_1593),
.B(n_1570),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1587),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1594),
.B(n_1570),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1590),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1584),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1599),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1597),
.Y(n_1612)
);

AO21x1_ASAP7_75t_L g1613 ( 
.A1(n_1586),
.A2(n_1568),
.B(n_1557),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1596),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1603),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1601),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1598),
.B(n_1573),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1592),
.B(n_1572),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1582),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1582),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1589),
.B(n_1580),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1600),
.B(n_1568),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1600),
.B(n_1573),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1619),
.A2(n_1585),
.B1(n_1464),
.B2(n_1595),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1604),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1605),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1607),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1620),
.B(n_1559),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1610),
.Y(n_1629)
);

NAND4xp25_ASAP7_75t_L g1630 ( 
.A(n_1616),
.B(n_1591),
.C(n_1602),
.D(n_1464),
.Y(n_1630)
);

AOI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1612),
.A2(n_1613),
.B1(n_1621),
.B2(n_1622),
.C(n_1618),
.Y(n_1631)
);

OAI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1621),
.A2(n_1495),
.B(n_1559),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1615),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1609),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1626),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1627),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1633),
.B(n_1611),
.Y(n_1637)
);

NOR2x1_ASAP7_75t_L g1638 ( 
.A(n_1630),
.B(n_1614),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1628),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1625),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1634),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1629),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1624),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_SL g1644 ( 
.A1(n_1632),
.A2(n_1622),
.B1(n_1631),
.B2(n_1623),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1642),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1637),
.Y(n_1646)
);

INVx5_ASAP7_75t_SL g1647 ( 
.A(n_1640),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1638),
.Y(n_1648)
);

BUFx4_ASAP7_75t_SL g1649 ( 
.A(n_1635),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1639),
.B(n_1624),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1636),
.B(n_1614),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1643),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1636),
.Y(n_1653)
);

NAND4xp25_ASAP7_75t_L g1654 ( 
.A(n_1651),
.B(n_1644),
.C(n_1641),
.D(n_1617),
.Y(n_1654)
);

OAI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1648),
.A2(n_1606),
.B(n_1608),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1650),
.A2(n_1645),
.B(n_1653),
.Y(n_1656)
);

NOR2x1_ASAP7_75t_L g1657 ( 
.A(n_1646),
.B(n_1608),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1647),
.B(n_1572),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1652),
.A2(n_1488),
.B1(n_1553),
.B2(n_1577),
.C(n_1569),
.Y(n_1659)
);

NOR4xp25_ASAP7_75t_L g1660 ( 
.A(n_1649),
.B(n_1575),
.C(n_1555),
.D(n_1556),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_SL g1661 ( 
.A(n_1647),
.B(n_1571),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1653),
.Y(n_1662)
);

AOI221x1_ASAP7_75t_L g1663 ( 
.A1(n_1651),
.A2(n_1499),
.B1(n_1439),
.B2(n_1544),
.C(n_1551),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1662),
.Y(n_1664)
);

AOI322xp5_ASAP7_75t_L g1665 ( 
.A1(n_1659),
.A2(n_1657),
.A3(n_1661),
.B1(n_1658),
.B2(n_1656),
.C1(n_1654),
.C2(n_1660),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1655),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1663),
.A2(n_1506),
.B1(n_1553),
.B2(n_1488),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1661),
.A2(n_1565),
.B1(n_1499),
.B2(n_1563),
.Y(n_1668)
);

AOI321xp33_ASAP7_75t_L g1669 ( 
.A1(n_1656),
.A2(n_1487),
.A3(n_1505),
.B1(n_1549),
.B2(n_1565),
.C(n_1496),
.Y(n_1669)
);

OAI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1660),
.A2(n_1551),
.B1(n_1544),
.B2(n_1567),
.C(n_1563),
.Y(n_1670)
);

NAND3xp33_ASAP7_75t_L g1671 ( 
.A(n_1665),
.B(n_1552),
.C(n_1567),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1664),
.Y(n_1672)
);

OAI211xp5_ASAP7_75t_L g1673 ( 
.A1(n_1666),
.A2(n_1431),
.B(n_1460),
.C(n_1552),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1669),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1668),
.Y(n_1675)
);

XNOR2x1_ASAP7_75t_L g1676 ( 
.A(n_1667),
.B(n_1549),
.Y(n_1676)
);

INVxp67_ASAP7_75t_SL g1677 ( 
.A(n_1670),
.Y(n_1677)
);

AND4x1_ASAP7_75t_L g1678 ( 
.A(n_1666),
.B(n_1542),
.C(n_219),
.D(n_222),
.Y(n_1678)
);

NAND4xp75_ASAP7_75t_L g1679 ( 
.A(n_1666),
.B(n_1552),
.C(n_1542),
.D(n_230),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_R g1680 ( 
.A(n_1672),
.B(n_216),
.Y(n_1680)
);

NAND2xp33_ASAP7_75t_SL g1681 ( 
.A(n_1674),
.B(n_1491),
.Y(n_1681)
);

NAND2xp33_ASAP7_75t_SL g1682 ( 
.A(n_1675),
.B(n_1337),
.Y(n_1682)
);

NAND2xp33_ASAP7_75t_SL g1683 ( 
.A(n_1671),
.B(n_223),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_R g1684 ( 
.A(n_1677),
.B(n_231),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1678),
.B(n_232),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_R g1686 ( 
.A(n_1679),
.B(n_243),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_R g1687 ( 
.A(n_1673),
.B(n_245),
.Y(n_1687)
);

A2O1A1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1683),
.A2(n_1681),
.B(n_1685),
.C(n_1682),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1684),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1680),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_SL g1691 ( 
.A(n_1686),
.B(n_1676),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1687),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1683),
.B(n_247),
.Y(n_1693)
);

CKINVDCx20_ASAP7_75t_R g1694 ( 
.A(n_1684),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1688),
.A2(n_1332),
.B(n_262),
.Y(n_1695)
);

INVx5_ASAP7_75t_L g1696 ( 
.A(n_1694),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1693),
.A2(n_248),
.B(n_265),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1692),
.A2(n_1690),
.B1(n_1689),
.B2(n_1691),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1691),
.A2(n_267),
.B1(n_270),
.B2(n_272),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1689),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1696),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1696),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1700),
.Y(n_1703)
);

OA21x2_ASAP7_75t_L g1704 ( 
.A1(n_1698),
.A2(n_275),
.B(n_276),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1697),
.Y(n_1705)
);

AOI31xp33_ASAP7_75t_L g1706 ( 
.A1(n_1702),
.A2(n_1695),
.A3(n_1699),
.B(n_281),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1705),
.A2(n_278),
.B1(n_279),
.B2(n_282),
.Y(n_1707)
);

AOI31xp33_ASAP7_75t_L g1708 ( 
.A1(n_1701),
.A2(n_283),
.A3(n_284),
.B(n_285),
.Y(n_1708)
);

XNOR2xp5_ASAP7_75t_L g1709 ( 
.A(n_1707),
.B(n_1704),
.Y(n_1709)
);

NAND4xp75_ASAP7_75t_L g1710 ( 
.A(n_1706),
.B(n_1704),
.C(n_1703),
.D(n_296),
.Y(n_1710)
);

XNOR2xp5_ASAP7_75t_L g1711 ( 
.A(n_1708),
.B(n_342),
.Y(n_1711)
);

AOI321xp33_ASAP7_75t_L g1712 ( 
.A1(n_1710),
.A2(n_289),
.A3(n_295),
.B1(n_297),
.B2(n_298),
.C(n_300),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1709),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1713),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1712),
.Y(n_1715)
);

CKINVDCx20_ASAP7_75t_R g1716 ( 
.A(n_1713),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1714),
.A2(n_1711),
.B1(n_303),
.B2(n_304),
.C(n_305),
.Y(n_1717)
);

OAI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1717),
.A2(n_1716),
.B1(n_1715),
.B2(n_308),
.Y(n_1718)
);


endmodule