module fake_aes_8990_n_722 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_722);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_722;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_L g81 ( .A(n_47), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_44), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_64), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_73), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_79), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_55), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_21), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_20), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_63), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_12), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_36), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_26), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_9), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_56), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_27), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_5), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_43), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_49), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_9), .Y(n_99) );
BUFx3_ASAP7_75t_L g100 ( .A(n_17), .Y(n_100) );
INVxp33_ASAP7_75t_L g101 ( .A(n_21), .Y(n_101) );
INVxp33_ASAP7_75t_L g102 ( .A(n_58), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_51), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_80), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_13), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_4), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_38), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_65), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_8), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_16), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_48), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_26), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_35), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_74), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_50), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_33), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_77), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_71), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_37), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_7), .Y(n_120) );
INVxp33_ASAP7_75t_L g121 ( .A(n_27), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_6), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_8), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_19), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_62), .Y(n_125) );
INVxp33_ASAP7_75t_L g126 ( .A(n_54), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_20), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_42), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_40), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_1), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_87), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_99), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_99), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_99), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_125), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_83), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_125), .Y(n_137) );
BUFx8_ASAP7_75t_L g138 ( .A(n_125), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_101), .B(n_0), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_121), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_83), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_100), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_84), .B(n_2), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_100), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_100), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_93), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_83), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_88), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_85), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_85), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_86), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_88), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_87), .B(n_3), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_95), .B(n_6), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_88), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_86), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_109), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_90), .A2(n_7), .B1(n_10), .B2(n_11), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_84), .Y(n_160) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_108), .B(n_78), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_95), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_109), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_109), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_110), .Y(n_165) );
NAND2xp33_ASAP7_75t_SL g166 ( .A(n_81), .B(n_10), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_97), .B(n_11), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_108), .B(n_12), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_110), .Y(n_169) );
AND2x6_ASAP7_75t_L g170 ( .A(n_97), .B(n_39), .Y(n_170) );
XNOR2xp5_ASAP7_75t_L g171 ( .A(n_92), .B(n_13), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_98), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_114), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_110), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
INVx2_ASAP7_75t_SL g176 ( .A(n_138), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_131), .B(n_102), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_144), .B(n_126), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_136), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_162), .A2(n_123), .B1(n_106), .B2(n_96), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_170), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_136), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
AND2x6_ASAP7_75t_L g188 ( .A(n_143), .B(n_115), .Y(n_188) );
INVx5_ASAP7_75t_L g189 ( .A(n_170), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_134), .B(n_130), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_136), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_160), .B(n_94), .Y(n_192) );
NAND2x1p5_ASAP7_75t_L g193 ( .A(n_143), .B(n_130), .Y(n_193) );
INVxp67_ASAP7_75t_L g194 ( .A(n_139), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_134), .B(n_122), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_134), .B(n_122), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_136), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_136), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_172), .B(n_94), .Y(n_199) );
INVx8_ASAP7_75t_L g200 ( .A(n_170), .Y(n_200) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_161), .B(n_129), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_172), .B(n_91), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_157), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_136), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_161), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_141), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_141), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_157), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_134), .B(n_123), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_141), .Y(n_210) );
BUFx2_ASAP7_75t_L g211 ( .A(n_138), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_141), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_141), .Y(n_213) );
NAND2x1p5_ASAP7_75t_L g214 ( .A(n_161), .B(n_112), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_172), .B(n_112), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_138), .B(n_89), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_141), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_152), .B(n_129), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_138), .B(n_128), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_152), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_166), .A2(n_106), .B1(n_127), .B2(n_124), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_152), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_171), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_152), .B(n_157), .Y(n_224) );
NAND3x1_ASAP7_75t_L g225 ( .A(n_173), .B(n_96), .C(n_127), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_132), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_132), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_152), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_133), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_152), .Y(n_230) );
AND2x6_ASAP7_75t_L g231 ( .A(n_148), .B(n_128), .Y(n_231) );
AND2x6_ASAP7_75t_L g232 ( .A(n_148), .B(n_113), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_133), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_142), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_142), .B(n_113), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_170), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_149), .B(n_124), .Y(n_237) );
AO22x2_ASAP7_75t_L g238 ( .A1(n_140), .A2(n_82), .B1(n_118), .B2(n_117), .Y(n_238) );
BUFx4f_ASAP7_75t_L g239 ( .A(n_170), .Y(n_239) );
INVxp67_ASAP7_75t_L g240 ( .A(n_168), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_145), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_145), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_146), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_176), .B(n_211), .Y(n_244) );
BUFx2_ASAP7_75t_L g245 ( .A(n_188), .Y(n_245) );
CKINVDCx16_ASAP7_75t_R g246 ( .A(n_180), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_175), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_178), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_177), .B(n_154), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_230), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_190), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_211), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_223), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_176), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_201), .A2(n_140), .B1(n_173), .B2(n_119), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_205), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_193), .A2(n_155), .B(n_154), .C(n_159), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_194), .B(n_167), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_179), .A2(n_146), .B(n_135), .C(n_137), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_205), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_180), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_183), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_184), .B(n_155), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_185), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_201), .A2(n_170), .B1(n_148), .B2(n_120), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_188), .B(n_147), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_187), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_188), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_192), .B(n_82), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_202), .B(n_170), .Y(n_270) );
NAND2x1p5_ASAP7_75t_L g271 ( .A(n_184), .B(n_98), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_195), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_195), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_203), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_188), .B(n_147), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_230), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_200), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_199), .B(n_170), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_208), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_240), .B(n_149), .Y(n_280) );
AND2x2_ASAP7_75t_SL g281 ( .A(n_239), .B(n_103), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_193), .B(n_171), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_226), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_188), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_227), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_188), .B(n_149), .Y(n_286) );
BUFx3_ASAP7_75t_L g287 ( .A(n_200), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_215), .B(n_149), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_200), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_196), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_229), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_238), .A2(n_120), .B1(n_159), .B2(n_135), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_215), .B(n_163), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_230), .Y(n_294) );
AND2x4_ASAP7_75t_SL g295 ( .A(n_184), .B(n_103), .Y(n_295) );
INVxp67_ASAP7_75t_L g296 ( .A(n_196), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_237), .B(n_105), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_233), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_221), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_234), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_241), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_237), .B(n_174), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_182), .Y(n_303) );
BUFx4f_ASAP7_75t_L g304 ( .A(n_200), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_190), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_230), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_236), .B(n_104), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_190), .Y(n_308) );
BUFx4f_ASAP7_75t_L g309 ( .A(n_236), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_214), .A2(n_104), .B1(n_107), .B2(n_111), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_216), .B(n_107), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_230), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_220), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_214), .A2(n_135), .B1(n_137), .B2(n_165), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_237), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_220), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_242), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_247), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_261), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_266), .A2(n_238), .B1(n_209), .B2(n_231), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_304), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_266), .A2(n_238), .B1(n_209), .B2(n_231), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_304), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_283), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_252), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_266), .A2(n_238), .B1(n_225), .B2(n_219), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_268), .A2(n_239), .B1(n_225), .B2(n_236), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_249), .B(n_209), .Y(n_328) );
INVxp67_ASAP7_75t_L g329 ( .A(n_282), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_315), .Y(n_330) );
BUFx8_ASAP7_75t_L g331 ( .A(n_245), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_251), .Y(n_332) );
INVx4_ASAP7_75t_L g333 ( .A(n_304), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_246), .Y(n_334) );
OAI21xp33_ASAP7_75t_L g335 ( .A1(n_303), .A2(n_235), .B(n_243), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_253), .Y(n_336) );
INVx5_ASAP7_75t_L g337 ( .A(n_252), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_296), .B(n_239), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_282), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_252), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_303), .B(n_236), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_278), .A2(n_189), .B(n_236), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_252), .Y(n_343) );
AND3x2_ASAP7_75t_L g344 ( .A(n_275), .B(n_111), .C(n_116), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_275), .A2(n_232), .B1(n_231), .B2(n_189), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_252), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_277), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_272), .B(n_231), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_275), .A2(n_232), .B1(n_231), .B2(n_189), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_245), .Y(n_350) );
INVx4_ASAP7_75t_L g351 ( .A(n_268), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_277), .Y(n_352) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_299), .A2(n_164), .B1(n_153), .B2(n_174), .C1(n_169), .C2(n_165), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_247), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_295), .Y(n_355) );
INVxp67_ASAP7_75t_SL g356 ( .A(n_284), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_270), .A2(n_189), .B(n_224), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_273), .B(n_189), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_287), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_253), .Y(n_360) );
INVx4_ASAP7_75t_L g361 ( .A(n_287), .Y(n_361) );
CKINVDCx8_ASAP7_75t_R g362 ( .A(n_256), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_255), .A2(n_299), .B1(n_258), .B2(n_281), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_251), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_290), .B(n_231), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_263), .A2(n_224), .B(n_218), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_289), .B(n_232), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_254), .B(n_115), .Y(n_368) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_289), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_256), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_248), .Y(n_371) );
A2O1A1Ixp33_ASAP7_75t_L g372 ( .A1(n_283), .A2(n_137), .B(n_218), .C(n_164), .Y(n_372) );
NAND2xp33_ASAP7_75t_L g373 ( .A(n_271), .B(n_232), .Y(n_373) );
NOR2x1_ASAP7_75t_L g374 ( .A(n_373), .B(n_286), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g375 ( .A1(n_326), .A2(n_260), .B1(n_310), .B2(n_305), .Y(n_375) );
AOI21xp33_ASAP7_75t_L g376 ( .A1(n_336), .A2(n_257), .B(n_269), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_337), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_355), .B(n_254), .Y(n_378) );
INVx2_ASAP7_75t_SL g379 ( .A(n_337), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_370), .Y(n_380) );
AO31x2_ASAP7_75t_L g381 ( .A1(n_324), .A2(n_259), .A3(n_314), .B(n_285), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_337), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_336), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_318), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_328), .B(n_292), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_318), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_354), .B(n_293), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_333), .B(n_251), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_324), .Y(n_389) );
AO31x2_ASAP7_75t_L g390 ( .A1(n_354), .A2(n_317), .A3(n_285), .B(n_291), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_319), .B(n_297), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_371), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_371), .B(n_293), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_358), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_332), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_358), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_329), .B(n_297), .Y(n_397) );
A2O1A1Ixp33_ASAP7_75t_L g398 ( .A1(n_335), .A2(n_311), .B(n_317), .C(n_291), .Y(n_398) );
OAI221xp5_ASAP7_75t_L g399 ( .A1(n_363), .A2(n_280), .B1(n_265), .B2(n_260), .C(n_305), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_348), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_339), .A2(n_297), .B1(n_281), .B2(n_308), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_320), .A2(n_264), .B1(n_248), .B2(n_274), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_353), .B(n_302), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_322), .A2(n_308), .B1(n_305), .B2(n_302), .Y(n_404) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_360), .A2(n_308), .B1(n_271), .B2(n_298), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_360), .B(n_288), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_341), .A2(n_302), .B1(n_298), .B2(n_300), .Y(n_407) );
OAI321xp33_ASAP7_75t_L g408 ( .A1(n_375), .A2(n_327), .A3(n_345), .B1(n_349), .B2(n_116), .C(n_117), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_403), .A2(n_355), .B1(n_350), .B2(n_362), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_405), .A2(n_350), .B1(n_362), .B2(n_337), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_402), .A2(n_373), .B1(n_370), .B2(n_344), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_384), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_387), .B(n_262), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_384), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_407), .A2(n_337), .B1(n_271), .B2(n_274), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_376), .A2(n_338), .B1(n_334), .B2(n_330), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_399), .A2(n_338), .B1(n_334), .B2(n_331), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_392), .B(n_262), .Y(n_418) );
OAI211xp5_ASAP7_75t_L g419 ( .A1(n_401), .A2(n_169), .B(n_153), .C(n_163), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_387), .B(n_346), .Y(n_420) );
AOI33xp33_ASAP7_75t_L g421 ( .A1(n_404), .A2(n_156), .A3(n_158), .B1(n_118), .B2(n_364), .B3(n_264), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_384), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_392), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_402), .A2(n_300), .B1(n_301), .B2(n_372), .C(n_279), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_386), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_406), .A2(n_351), .B1(n_333), .B2(n_365), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_406), .A2(n_331), .B1(n_368), .B2(n_301), .Y(n_427) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_380), .A2(n_351), .B1(n_333), .B2(n_361), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_385), .A2(n_331), .B1(n_279), .B2(n_267), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_393), .A2(n_267), .B1(n_367), .B2(n_361), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_386), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_393), .A2(n_232), .B1(n_295), .B2(n_356), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_386), .B(n_346), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_398), .A2(n_351), .B1(n_361), .B2(n_340), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_390), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_397), .B(n_367), .Y(n_436) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_412), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_411), .A2(n_389), .B1(n_391), .B2(n_379), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_435), .B(n_390), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_425), .Y(n_440) );
OAI31xp33_ASAP7_75t_L g441 ( .A1(n_409), .A2(n_397), .A3(n_391), .B(n_396), .Y(n_441) );
OAI211xp5_ASAP7_75t_L g442 ( .A1(n_411), .A2(n_383), .B(n_156), .C(n_158), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_425), .Y(n_443) );
OAI33xp33_ASAP7_75t_L g444 ( .A1(n_428), .A2(n_396), .A3(n_394), .B1(n_389), .B2(n_400), .B3(n_378), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_435), .B(n_390), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_431), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_423), .B(n_390), .Y(n_447) );
OA21x2_ASAP7_75t_L g448 ( .A1(n_424), .A2(n_400), .B(n_394), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_431), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_423), .B(n_390), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_420), .B(n_390), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_417), .A2(n_388), .B1(n_377), .B2(n_379), .Y(n_452) );
OAI33xp33_ASAP7_75t_L g453 ( .A1(n_410), .A2(n_395), .A3(n_228), .B1(n_212), .B2(n_217), .B3(n_210), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_412), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_414), .Y(n_455) );
BUFx3_ASAP7_75t_L g456 ( .A(n_420), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_414), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_413), .B(n_382), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_422), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_416), .A2(n_395), .B1(n_388), .B2(n_366), .C(n_377), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_429), .A2(n_388), .B1(n_374), .B2(n_395), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_436), .A2(n_388), .B1(n_374), .B2(n_382), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_413), .B(n_382), .Y(n_463) );
NAND4xp25_ASAP7_75t_SL g464 ( .A(n_427), .B(n_14), .C(n_15), .D(n_17), .Y(n_464) );
BUFx2_ASAP7_75t_L g465 ( .A(n_422), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_419), .A2(n_382), .B1(n_307), .B2(n_367), .C(n_343), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_418), .B(n_381), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_432), .A2(n_325), .B1(n_340), .B2(n_343), .Y(n_468) );
AOI211xp5_ASAP7_75t_L g469 ( .A1(n_408), .A2(n_244), .B(n_191), .C(n_181), .Y(n_469) );
OAI31xp33_ASAP7_75t_SL g470 ( .A1(n_426), .A2(n_381), .A3(n_19), .B(n_22), .Y(n_470) );
AOI222xp33_ASAP7_75t_SL g471 ( .A1(n_415), .A2(n_18), .B1(n_22), .B2(n_23), .C1(n_24), .C2(n_25), .Y(n_471) );
OAI211xp5_ASAP7_75t_SL g472 ( .A1(n_421), .A2(n_222), .B(n_228), .C(n_186), .Y(n_472) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_434), .A2(n_186), .B(n_198), .Y(n_473) );
OAI21xp33_ASAP7_75t_L g474 ( .A1(n_432), .A2(n_198), .B(n_210), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_447), .B(n_420), .Y(n_475) );
OAI221xp5_ASAP7_75t_L g476 ( .A1(n_470), .A2(n_430), .B1(n_418), .B2(n_433), .C(n_340), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_438), .A2(n_420), .B1(n_433), .B2(n_232), .Y(n_477) );
AOI211x1_ASAP7_75t_L g478 ( .A1(n_464), .A2(n_18), .B(n_23), .C(n_24), .Y(n_478) );
NAND2x1_ASAP7_75t_L g479 ( .A(n_447), .B(n_325), .Y(n_479) );
NAND4xp25_ASAP7_75t_L g480 ( .A(n_441), .B(n_212), .C(n_217), .D(n_25), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_467), .B(n_381), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_442), .A2(n_357), .B(n_343), .Y(n_482) );
OAI31xp33_ASAP7_75t_L g483 ( .A1(n_472), .A2(n_325), .A3(n_222), .B(n_342), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_465), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_465), .Y(n_485) );
OAI21xp33_ASAP7_75t_L g486 ( .A1(n_447), .A2(n_181), .B(n_197), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_450), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_439), .B(n_381), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_450), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_450), .B(n_369), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_459), .Y(n_491) );
AOI221xp5_ASAP7_75t_L g492 ( .A1(n_444), .A2(n_222), .B1(n_191), .B2(n_181), .C(n_213), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_467), .B(n_381), .Y(n_493) );
AOI31xp67_ASAP7_75t_L g494 ( .A1(n_459), .A2(n_294), .A3(n_250), .B(n_276), .Y(n_494) );
AOI33xp33_ASAP7_75t_L g495 ( .A1(n_461), .A2(n_313), .A3(n_316), .B1(n_306), .B2(n_312), .B3(n_250), .Y(n_495) );
AND2x2_ASAP7_75t_SL g496 ( .A(n_451), .B(n_323), .Y(n_496) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_460), .A2(n_181), .B1(n_204), .B2(n_206), .C(n_207), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_439), .B(n_381), .Y(n_498) );
OAI221xp5_ASAP7_75t_L g499 ( .A1(n_452), .A2(n_181), .B1(n_191), .B2(n_197), .C(n_204), .Y(n_499) );
BUFx2_ASAP7_75t_L g500 ( .A(n_451), .Y(n_500) );
OAI222xp33_ASAP7_75t_L g501 ( .A1(n_451), .A2(n_28), .B1(n_29), .B2(n_30), .C1(n_31), .C2(n_32), .Y(n_501) );
INVxp33_ASAP7_75t_L g502 ( .A(n_458), .Y(n_502) );
OAI31xp33_ASAP7_75t_L g503 ( .A1(n_458), .A2(n_294), .A3(n_276), .B(n_306), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_445), .B(n_34), .Y(n_504) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_437), .A2(n_312), .B(n_316), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_463), .B(n_369), .Y(n_506) );
OAI221xp5_ASAP7_75t_L g507 ( .A1(n_462), .A2(n_191), .B1(n_197), .B2(n_204), .C(n_206), .Y(n_507) );
INVxp67_ASAP7_75t_SL g508 ( .A(n_445), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_471), .A2(n_359), .B1(n_352), .B2(n_347), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_440), .B(n_41), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_463), .B(n_369), .Y(n_511) );
BUFx2_ASAP7_75t_L g512 ( .A(n_454), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_440), .B(n_45), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_443), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_454), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_456), .Y(n_516) );
INVx4_ASAP7_75t_L g517 ( .A(n_456), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_443), .B(n_207), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_446), .B(n_369), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_446), .B(n_46), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_449), .B(n_52), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_449), .B(n_53), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_455), .B(n_57), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_457), .B(n_59), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_448), .A2(n_369), .B1(n_359), .B2(n_352), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_457), .B(n_359), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_473), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_514), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_487), .B(n_448), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_508), .B(n_448), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_514), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_515), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_512), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_512), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_487), .B(n_489), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_489), .B(n_448), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_484), .Y(n_537) );
NOR3xp33_ASAP7_75t_L g538 ( .A(n_480), .B(n_453), .C(n_469), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_500), .B(n_473), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_500), .B(n_60), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_485), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_475), .B(n_473), .Y(n_542) );
AOI21xp33_ASAP7_75t_L g543 ( .A1(n_479), .A2(n_468), .B(n_474), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_491), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_475), .B(n_204), .Y(n_545) );
AOI31xp33_ASAP7_75t_L g546 ( .A1(n_502), .A2(n_466), .A3(n_66), .B(n_67), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_481), .B(n_206), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_485), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_488), .B(n_61), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_491), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_488), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_478), .B(n_206), .C(n_213), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_493), .B(n_206), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_505), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_498), .B(n_68), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_505), .Y(n_556) );
INVx2_ASAP7_75t_SL g557 ( .A(n_479), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_498), .B(n_207), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_516), .B(n_207), .Y(n_559) );
AND3x1_ASAP7_75t_L g560 ( .A(n_509), .B(n_69), .C(n_70), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_496), .B(n_197), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_517), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_504), .B(n_191), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_517), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_517), .B(n_72), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_490), .B(n_197), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_519), .B(n_204), .Y(n_567) );
OAI211xp5_ASAP7_75t_SL g568 ( .A1(n_509), .A2(n_313), .B(n_76), .C(n_75), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_518), .Y(n_569) );
OAI221xp5_ASAP7_75t_SL g570 ( .A1(n_477), .A2(n_213), .B1(n_347), .B2(n_352), .C(n_359), .Y(n_570) );
OAI33xp33_ASAP7_75t_L g571 ( .A1(n_506), .A2(n_213), .A3(n_347), .B1(n_352), .B2(n_359), .B3(n_321), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_496), .B(n_213), .Y(n_572) );
BUFx2_ASAP7_75t_L g573 ( .A(n_496), .Y(n_573) );
BUFx2_ASAP7_75t_L g574 ( .A(n_505), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_511), .B(n_352), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_505), .Y(n_576) );
INVx3_ASAP7_75t_L g577 ( .A(n_527), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_526), .B(n_518), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_527), .B(n_347), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_478), .B(n_347), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_494), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_525), .Y(n_582) );
BUFx2_ASAP7_75t_L g583 ( .A(n_510), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_525), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_510), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_494), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_495), .B(n_321), .C(n_323), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_551), .B(n_520), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_528), .Y(n_589) );
NAND4xp25_ASAP7_75t_L g590 ( .A(n_538), .B(n_476), .C(n_492), .D(n_497), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_551), .B(n_486), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_531), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_532), .B(n_513), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_583), .A2(n_510), .B1(n_521), .B2(n_522), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_531), .Y(n_595) );
AOI31xp33_ASAP7_75t_L g596 ( .A1(n_560), .A2(n_513), .A3(n_520), .B(n_522), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_542), .B(n_521), .Y(n_597) );
AND2x2_ASAP7_75t_SL g598 ( .A(n_583), .B(n_524), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_542), .B(n_524), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_564), .Y(n_600) );
BUFx2_ASAP7_75t_L g601 ( .A(n_564), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_532), .B(n_523), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_537), .B(n_483), .C(n_482), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_533), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_535), .B(n_523), .Y(n_605) );
OAI21x1_ASAP7_75t_SL g606 ( .A1(n_562), .A2(n_501), .B(n_499), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_533), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_571), .A2(n_507), .B(n_503), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_534), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g610 ( .A1(n_546), .A2(n_309), .B(n_321), .Y(n_610) );
AOI211xp5_ASAP7_75t_L g611 ( .A1(n_552), .A2(n_321), .B(n_323), .C(n_309), .Y(n_611) );
INVxp67_ASAP7_75t_SL g612 ( .A(n_541), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_535), .B(n_309), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_557), .B(n_321), .Y(n_614) );
XNOR2xp5_ASAP7_75t_L g615 ( .A(n_562), .B(n_323), .Y(n_615) );
AOI211x1_ASAP7_75t_SL g616 ( .A1(n_568), .A2(n_323), .B(n_580), .C(n_543), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_534), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_569), .B(n_529), .Y(n_618) );
NOR3xp33_ASAP7_75t_L g619 ( .A(n_565), .B(n_553), .C(n_547), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_540), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_578), .B(n_548), .Y(n_621) );
INVxp33_ASAP7_75t_SL g622 ( .A(n_573), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_549), .A2(n_555), .B1(n_585), .B2(n_582), .Y(n_623) );
AND2x2_ASAP7_75t_SL g624 ( .A(n_573), .B(n_540), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_569), .B(n_529), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_585), .B(n_555), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_544), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_536), .B(n_578), .Y(n_628) );
AND3x2_ASAP7_75t_L g629 ( .A(n_540), .B(n_574), .C(n_555), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_550), .Y(n_630) );
NAND2xp5_ASAP7_75t_R g631 ( .A(n_557), .B(n_549), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_536), .B(n_539), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_558), .B(n_530), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_549), .B(n_545), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_539), .B(n_584), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_621), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_624), .B(n_574), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_612), .B(n_530), .Y(n_638) );
AND2x4_ASAP7_75t_L g639 ( .A(n_601), .B(n_577), .Y(n_639) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_629), .A2(n_587), .B(n_577), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_622), .B(n_577), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_589), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_596), .A2(n_570), .B(n_554), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_635), .B(n_584), .Y(n_644) );
XNOR2xp5_ASAP7_75t_L g645 ( .A(n_624), .B(n_545), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_598), .A2(n_554), .B1(n_556), .B2(n_576), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_592), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_595), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_604), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_607), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_635), .B(n_582), .Y(n_651) );
INVx4_ASAP7_75t_SL g652 ( .A(n_615), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_622), .B(n_558), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_609), .Y(n_654) );
NOR3xp33_ASAP7_75t_L g655 ( .A(n_590), .B(n_603), .C(n_610), .Y(n_655) );
AOI321xp33_ASAP7_75t_L g656 ( .A1(n_623), .A2(n_561), .A3(n_572), .B1(n_579), .B2(n_563), .C(n_575), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_617), .Y(n_657) );
INVx4_ASAP7_75t_L g658 ( .A(n_629), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_SL g659 ( .A1(n_600), .A2(n_556), .B(n_576), .C(n_575), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_598), .B(n_579), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_628), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g662 ( .A1(n_608), .A2(n_561), .B(n_572), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_618), .Y(n_663) );
AOI311xp33_ASAP7_75t_L g664 ( .A1(n_626), .A2(n_567), .A3(n_559), .B(n_586), .C(n_581), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_625), .A2(n_581), .B1(n_586), .B2(n_559), .C(n_566), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_633), .B(n_566), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_605), .B(n_597), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_606), .A2(n_611), .B(n_619), .C(n_593), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_623), .A2(n_594), .B1(n_620), .B2(n_626), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_627), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g671 ( .A1(n_634), .A2(n_591), .B1(n_631), .B2(n_602), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_588), .A2(n_597), .B1(n_599), .B2(n_591), .Y(n_672) );
INVxp67_ASAP7_75t_L g673 ( .A(n_630), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_599), .Y(n_674) );
AOI222xp33_ASAP7_75t_L g675 ( .A1(n_613), .A2(n_159), .B1(n_635), .B2(n_624), .C1(n_598), .C2(n_551), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_614), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_613), .B(n_614), .Y(n_677) );
OAI211xp5_ASAP7_75t_L g678 ( .A1(n_616), .A2(n_623), .B(n_601), .C(n_594), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_614), .B(n_635), .Y(n_679) );
XNOR2x1_ASAP7_75t_L g680 ( .A(n_629), .B(n_171), .Y(n_680) );
INVxp67_ASAP7_75t_L g681 ( .A(n_601), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_632), .B(n_635), .Y(n_682) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_596), .A2(n_546), .B(n_538), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_632), .B(n_635), .Y(n_684) );
XNOR2xp5_ASAP7_75t_L g685 ( .A(n_624), .B(n_380), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_685), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_638), .B(n_672), .Y(n_687) );
OAI211xp5_ASAP7_75t_L g688 ( .A1(n_683), .A2(n_655), .B(n_675), .C(n_668), .Y(n_688) );
AO221x1_ASAP7_75t_L g689 ( .A1(n_671), .A2(n_646), .B1(n_669), .B2(n_681), .C(n_658), .Y(n_689) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_685), .B(n_658), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_674), .Y(n_691) );
O2A1O1Ixp33_ASAP7_75t_L g692 ( .A1(n_678), .A2(n_659), .B(n_640), .C(n_637), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g693 ( .A1(n_680), .A2(n_662), .B(n_638), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_680), .B(n_664), .C(n_643), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_654), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_657), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_684), .B(n_682), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_637), .A2(n_660), .B1(n_641), .B2(n_679), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_660), .A2(n_677), .B1(n_641), .B2(n_636), .Y(n_699) );
INVx1_ASAP7_75t_SL g700 ( .A(n_690), .Y(n_700) );
NOR5xp2_ASAP7_75t_L g701 ( .A(n_694), .B(n_673), .C(n_670), .D(n_652), .E(n_661), .Y(n_701) );
OAI221xp5_ASAP7_75t_SL g702 ( .A1(n_688), .A2(n_692), .B1(n_686), .B2(n_699), .C(n_698), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_688), .B(n_665), .C(n_659), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_695), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_693), .B(n_663), .Y(n_705) );
OAI211xp5_ASAP7_75t_SL g706 ( .A1(n_689), .A2(n_656), .B(n_651), .C(n_644), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_687), .A2(n_639), .B(n_645), .Y(n_707) );
OA22x2_ASAP7_75t_L g708 ( .A1(n_700), .A2(n_691), .B1(n_697), .B2(n_696), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_702), .A2(n_667), .B1(n_682), .B2(n_684), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_706), .A2(n_652), .B1(n_639), .B2(n_653), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_703), .A2(n_652), .B1(n_653), .B2(n_650), .Y(n_711) );
AND2x4_ASAP7_75t_L g712 ( .A(n_707), .B(n_705), .Y(n_712) );
NOR2xp67_ASAP7_75t_L g713 ( .A(n_710), .B(n_704), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_708), .Y(n_714) );
XOR2xp5_ASAP7_75t_L g715 ( .A(n_712), .B(n_666), .Y(n_715) );
NOR2x1_ASAP7_75t_L g716 ( .A(n_714), .B(n_709), .Y(n_716) );
AOI222xp33_ASAP7_75t_L g717 ( .A1(n_713), .A2(n_701), .B1(n_711), .B2(n_649), .C1(n_647), .C2(n_648), .Y(n_717) );
OAI21xp33_ASAP7_75t_L g718 ( .A1(n_716), .A2(n_715), .B(n_676), .Y(n_718) );
XNOR2x1_ASAP7_75t_L g719 ( .A(n_717), .B(n_676), .Y(n_719) );
AND2x2_ASAP7_75t_SL g720 ( .A(n_718), .B(n_642), .Y(n_720) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_720), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_720), .B(n_719), .Y(n_722) );
endmodule