module fake_aes_9314_n_30 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
AND2x2_ASAP7_75t_L g13 ( .A(n_9), .B(n_11), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_7), .B(n_1), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_3), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_3), .B(n_1), .Y(n_18) );
NAND2x1p5_ASAP7_75t_L g19 ( .A(n_18), .B(n_0), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_16), .B(n_0), .Y(n_20) );
AOI21xp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_13), .B(n_14), .Y(n_21) );
OA21x2_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_15), .B(n_13), .Y(n_22) );
AND2x4_ASAP7_75t_L g23 ( .A(n_22), .B(n_18), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AOI221xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_23), .B1(n_19), .B2(n_16), .C(n_17), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_2), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_25), .B(n_2), .Y(n_28) );
OAI221xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_17), .B1(n_8), .B2(n_10), .C(n_12), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_27), .B1(n_17), .B2(n_5), .Y(n_30) );
endmodule