module real_jpeg_18059_n_4 (n_3, n_1, n_0, n_2, n_4);

input n_3;
input n_1;
input n_0;
input n_2;

output n_4;

wire n_5;
wire n_8;
wire n_12;
wire n_11;
wire n_13;
wire n_6;
wire n_7;
wire n_10;
wire n_9;

INVx1_ASAP7_75t_SL g7 ( 
.A(n_0),
.Y(n_7)
);

INVx2_ASAP7_75t_R g5 ( 
.A(n_1),
.Y(n_5)
);

OAI322xp33_ASAP7_75t_L g4 ( 
.A1(n_2),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_4)
);

INVx2_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

INVx2_ASAP7_75t_SL g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_12),
.Y(n_10)
);

BUFx12f_ASAP7_75t_SL g12 ( 
.A(n_13),
.Y(n_12)
);


endmodule