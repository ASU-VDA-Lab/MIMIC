module fake_jpeg_23335_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_7),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_19),
.Y(n_22)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_8),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_10),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_0),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_15),
.B1(n_11),
.B2(n_8),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_30),
.B1(n_34),
.B2(n_22),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_15),
.B1(n_11),
.B2(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_35),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_20),
.B1(n_18),
.B2(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_24),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_40),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_44),
.B1(n_37),
.B2(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_24),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_47),
.A2(n_32),
.B(n_29),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_44),
.C(n_41),
.Y(n_48)
);

OAI321xp33_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_49),
.A3(n_45),
.B1(n_36),
.B2(n_37),
.C(n_5),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_51),
.Y(n_52)
);

A2O1A1O1Ixp25_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_1),
.B(n_2),
.C(n_3),
.D(n_6),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_7),
.Y(n_54)
);


endmodule