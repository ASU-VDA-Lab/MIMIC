module fake_aes_1233_n_43 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_43);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_43;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_33;
wire n_30;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_SL g11 ( .A(n_1), .B(n_0), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_3), .Y(n_12) );
CKINVDCx16_ASAP7_75t_R g13 ( .A(n_1), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_2), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_10), .B(n_2), .Y(n_16) );
NAND2xp33_ASAP7_75t_SL g17 ( .A(n_9), .B(n_4), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_13), .B(n_0), .Y(n_18) );
NOR2xp33_ASAP7_75t_R g19 ( .A(n_12), .B(n_3), .Y(n_19) );
AOI22xp33_ASAP7_75t_L g20 ( .A1(n_15), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_13), .B(n_9), .Y(n_21) );
INVx1_ASAP7_75t_SL g22 ( .A(n_14), .Y(n_22) );
BUFx12f_ASAP7_75t_L g23 ( .A(n_16), .Y(n_23) );
INVx3_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_15), .Y(n_25) );
OAI22xp33_ASAP7_75t_SL g26 ( .A1(n_18), .A2(n_11), .B1(n_17), .B2(n_7), .Y(n_26) );
INVx3_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
A2O1A1Ixp33_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_21), .B(n_16), .C(n_22), .Y(n_28) );
NAND3xp33_ASAP7_75t_L g29 ( .A(n_25), .B(n_20), .C(n_16), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_22), .B1(n_17), .B2(n_11), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_28), .B(n_27), .Y(n_31) );
OAI33xp33_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_26), .A3(n_19), .B1(n_24), .B2(n_27), .B3(n_8), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
NOR2xp33_ASAP7_75t_R g35 ( .A(n_32), .B(n_24), .Y(n_35) );
INVx1_ASAP7_75t_SL g36 ( .A(n_35), .Y(n_36) );
NAND2xp5_ASAP7_75t_L g37 ( .A(n_34), .B(n_24), .Y(n_37) );
INVx2_ASAP7_75t_L g38 ( .A(n_33), .Y(n_38) );
OR3x2_ASAP7_75t_L g39 ( .A(n_36), .B(n_33), .C(n_26), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_38), .Y(n_40) );
NAND3xp33_ASAP7_75t_SL g41 ( .A(n_37), .B(n_30), .C(n_6), .Y(n_41) );
OR2x6_ASAP7_75t_L g42 ( .A(n_40), .B(n_5), .Y(n_42) );
AOI22xp33_ASAP7_75t_L g43 ( .A1(n_42), .A2(n_39), .B1(n_41), .B2(n_32), .Y(n_43) );
endmodule