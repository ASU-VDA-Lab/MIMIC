module fake_jpeg_15048_n_187 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_34),
.B(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_32),
.Y(n_51)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_50),
.Y(n_64)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx9p33_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_70),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_67),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_23),
.B(n_19),
.C(n_17),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_63),
.B(n_66),
.C(n_73),
.Y(n_104)
);

OR2x2_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_21),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_18),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_72),
.Y(n_88)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_44),
.B(n_26),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_22),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_79),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_33),
.B1(n_40),
.B2(n_35),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_58),
.B1(n_39),
.B2(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_30),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_31),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_43),
.B(n_24),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_73),
.Y(n_116)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_100),
.B1(n_103),
.B2(n_74),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_97),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_42),
.C(n_41),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_77),
.C(n_93),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_20),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_101),
.Y(n_123)
);

AO22x1_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_41),
.B1(n_38),
.B2(n_43),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_16),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_61),
.A2(n_39),
.B1(n_29),
.B2(n_31),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_111),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_63),
.Y(n_110)
);

AOI221xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_26),
.B1(n_16),
.B2(n_27),
.C(n_23),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_73),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_84),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_116),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_76),
.Y(n_114)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_66),
.C(n_27),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_120),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_43),
.C(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_90),
.B(n_20),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_71),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_68),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_96),
.A3(n_100),
.B1(n_104),
.B2(n_90),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_130),
.B1(n_115),
.B2(n_117),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_100),
.B1(n_95),
.B2(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_131),
.B(n_115),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_32),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_134),
.C(n_108),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_105),
.A2(n_102),
.B(n_30),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_137),
.A2(n_139),
.B(n_140),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_29),
.B(n_19),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_79),
.B(n_2),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_150),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_123),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_149),
.C(n_151),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_133),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_129),
.B(n_109),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_109),
.C(n_107),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_21),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_153),
.C(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_107),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_160),
.C(n_163),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_130),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_161),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_146),
.B1(n_131),
.B2(n_17),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_124),
.C(n_140),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_137),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_126),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_167),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_146),
.C(n_112),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_32),
.C(n_135),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_87),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_162),
.A2(n_157),
.B(n_13),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_170),
.A2(n_8),
.B(n_14),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_162),
.B1(n_135),
.B2(n_74),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_172),
.A2(n_166),
.B(n_169),
.C(n_1),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_178),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_10),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_171),
.A2(n_80),
.B1(n_4),
.B2(n_1),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_4),
.C(n_5),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_176),
.A2(n_175),
.B(n_5),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_181),
.B(n_7),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_184),
.C(n_12),
.Y(n_185)
);

NOR2xp67_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_10),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_185),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_14),
.Y(n_187)
);


endmodule