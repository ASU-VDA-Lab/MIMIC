module real_aes_17023_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_103;
wire n_166;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
AND2x4_ASAP7_75t_L g111 ( .A(n_0), .B(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_1), .A2(n_3), .B1(n_151), .B2(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_2), .A2(n_43), .B1(n_158), .B2(n_271), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_4), .A2(n_24), .B1(n_252), .B2(n_271), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_5), .A2(n_17), .B1(n_148), .B2(n_207), .Y(n_206) );
AOI22x1_ASAP7_75t_SL g496 ( .A1(n_6), .A2(n_75), .B1(n_497), .B2(n_498), .Y(n_496) );
INVxp67_ASAP7_75t_SL g498 ( .A(n_6), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_7), .A2(n_60), .B1(n_189), .B2(n_254), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_8), .A2(n_18), .B1(n_158), .B2(n_193), .Y(n_544) );
INVx1_ASAP7_75t_L g112 ( .A(n_9), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_10), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_11), .A2(n_102), .B1(n_118), .B2(n_870), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_12), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_13), .A2(n_19), .B1(n_188), .B2(n_191), .Y(n_187) );
BUFx2_ASAP7_75t_L g115 ( .A(n_14), .Y(n_115) );
OR2x2_ASAP7_75t_L g127 ( .A(n_14), .B(n_38), .Y(n_127) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_15), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_16), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_20), .A2(n_99), .B1(n_148), .B2(n_151), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_21), .A2(n_39), .B1(n_203), .B2(n_204), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_22), .B(n_149), .Y(n_222) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_23), .A2(n_57), .B(n_167), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_25), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_26), .Y(n_607) );
INVx4_ASAP7_75t_R g538 ( .A(n_27), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_28), .B(n_155), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_29), .A2(n_47), .B1(n_175), .B2(n_178), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_30), .A2(n_53), .B1(n_148), .B2(n_178), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_31), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_32), .B(n_203), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_33), .Y(n_235) );
INVx1_ASAP7_75t_L g572 ( .A(n_34), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_35), .B(n_271), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_SL g617 ( .A1(n_36), .A2(n_154), .B(n_158), .C(n_618), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_37), .A2(n_54), .B1(n_158), .B2(n_178), .Y(n_605) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_38), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_40), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_41), .A2(n_87), .B1(n_158), .B2(n_251), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_42), .A2(n_46), .B1(n_158), .B2(n_193), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_44), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_45), .A2(n_58), .B1(n_148), .B2(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g581 ( .A(n_48), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_49), .B(n_158), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_50), .Y(n_554) );
INVx2_ASAP7_75t_L g507 ( .A(n_51), .Y(n_507) );
INVx1_ASAP7_75t_L g107 ( .A(n_52), .Y(n_107) );
BUFx3_ASAP7_75t_L g862 ( .A(n_52), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_55), .A2(n_88), .B1(n_158), .B2(n_178), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_56), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_59), .B(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_61), .A2(n_76), .B1(n_157), .B2(n_175), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_62), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_63), .A2(n_78), .B1(n_158), .B2(n_193), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_64), .A2(n_97), .B1(n_148), .B2(n_191), .Y(n_232) );
AND2x4_ASAP7_75t_L g144 ( .A(n_65), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g167 ( .A(n_66), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_67), .A2(n_90), .B1(n_175), .B2(n_178), .Y(n_568) );
AO22x1_ASAP7_75t_L g522 ( .A1(n_68), .A2(n_77), .B1(n_204), .B2(n_523), .Y(n_522) );
OAI22x1_ASAP7_75t_SL g852 ( .A1(n_69), .A2(n_72), .B1(n_853), .B2(n_854), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g853 ( .A(n_69), .Y(n_853) );
INVx1_ASAP7_75t_L g145 ( .A(n_70), .Y(n_145) );
AND2x2_ASAP7_75t_L g620 ( .A(n_71), .B(n_228), .Y(n_620) );
INVx1_ASAP7_75t_L g854 ( .A(n_72), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_73), .B(n_254), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_74), .Y(n_613) );
INVx1_ASAP7_75t_L g497 ( .A(n_75), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_79), .B(n_271), .Y(n_555) );
INVx2_ASAP7_75t_L g155 ( .A(n_80), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_81), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_82), .B(n_228), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_83), .A2(n_98), .B1(n_178), .B2(n_254), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_84), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_85), .B(n_165), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_86), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_89), .B(n_228), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_91), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_92), .B(n_228), .Y(n_551) );
INVx1_ASAP7_75t_L g110 ( .A(n_93), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_93), .B(n_125), .Y(n_124) );
NAND2xp33_ASAP7_75t_L g225 ( .A(n_94), .B(n_149), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_95), .A2(n_195), .B(n_254), .C(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g540 ( .A(n_96), .B(n_541), .Y(n_540) );
NAND2xp33_ASAP7_75t_L g559 ( .A(n_100), .B(n_176), .Y(n_559) );
CKINVDCx10_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx11_ASAP7_75t_R g873 ( .A(n_103), .Y(n_873) );
OR2x6_ASAP7_75t_L g103 ( .A(n_104), .B(n_113), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NOR2x1p5_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g125 ( .A(n_107), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_109), .Y(n_849) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g512 ( .A(n_110), .Y(n_512) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVxp33_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
OR2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_128), .Y(n_118) );
AOI21xp33_ASAP7_75t_L g129 ( .A1(n_119), .A2(n_130), .B(n_500), .Y(n_129) );
NOR2x1_ASAP7_75t_R g119 ( .A(n_120), .B(n_121), .Y(n_119) );
BUFx2_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx4_ASAP7_75t_L g502 ( .A(n_123), .Y(n_502) );
AND2x6_ASAP7_75t_SL g123 ( .A(n_124), .B(n_126), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_126), .B(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2x1_ASAP7_75t_L g861 ( .A(n_127), .B(n_862), .Y(n_861) );
OAI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_503), .B(n_508), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B1(n_496), .B2(n_499), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OA22x2_ASAP7_75t_L g509 ( .A1(n_132), .A2(n_510), .B1(n_513), .B2(n_848), .Y(n_509) );
AND3x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_393), .C(n_471), .Y(n_132) );
NOR2x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_336), .Y(n_133) );
NAND3xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_283), .C(n_306), .Y(n_134) );
AOI221x1_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_213), .B1(n_236), .B2(n_245), .C(n_258), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_183), .Y(n_136) );
AND2x4_ASAP7_75t_L g373 ( .A(n_137), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_171), .Y(n_138) );
INVx2_ASAP7_75t_L g332 ( .A(n_139), .Y(n_332) );
INVx1_ASAP7_75t_L g359 ( .A(n_139), .Y(n_359) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g239 ( .A(n_140), .Y(n_239) );
AND2x4_ASAP7_75t_L g310 ( .A(n_140), .B(n_240), .Y(n_310) );
AO31x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_146), .A3(n_162), .B(n_168), .Y(n_140) );
AO31x2_ASAP7_75t_L g230 ( .A1(n_141), .A2(n_196), .A3(n_231), .B(n_234), .Y(n_230) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_142), .A2(n_533), .B(n_536), .Y(n_532) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AO31x2_ASAP7_75t_L g185 ( .A1(n_143), .A2(n_186), .A3(n_196), .B(n_198), .Y(n_185) );
AO31x2_ASAP7_75t_L g200 ( .A1(n_143), .A2(n_201), .A3(n_209), .B(n_211), .Y(n_200) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_143), .A2(n_269), .A3(n_273), .B(n_274), .Y(n_268) );
AO31x2_ASAP7_75t_L g542 ( .A1(n_143), .A2(n_170), .A3(n_543), .B(n_546), .Y(n_542) );
BUFx10_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
INVx1_ASAP7_75t_L g529 ( .A(n_144), .Y(n_529) );
BUFx10_ASAP7_75t_L g563 ( .A(n_144), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_153), .B1(n_156), .B2(n_159), .Y(n_146) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_149), .Y(n_523) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g152 ( .A(n_150), .Y(n_152) );
INVx3_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_150), .Y(n_176) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
INVx1_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
INVx1_ASAP7_75t_L g205 ( .A(n_150), .Y(n_205) );
INVx1_ASAP7_75t_L g208 ( .A(n_150), .Y(n_208) );
INVx2_ASAP7_75t_L g252 ( .A(n_150), .Y(n_252) );
INVx1_ASAP7_75t_L g254 ( .A(n_150), .Y(n_254) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_150), .Y(n_271) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_152), .B(n_615), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g173 ( .A1(n_153), .A2(n_159), .B1(n_174), .B2(n_177), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_153), .A2(n_187), .B1(n_192), .B2(n_194), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_153), .A2(n_159), .B1(n_202), .B2(n_206), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_153), .A2(n_224), .B(n_225), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_153), .A2(n_194), .B1(n_232), .B2(n_233), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_153), .A2(n_250), .B1(n_253), .B2(n_255), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_153), .A2(n_159), .B1(n_270), .B2(n_272), .Y(n_269) );
OAI22x1_ASAP7_75t_L g543 ( .A1(n_153), .A2(n_255), .B1(n_544), .B2(n_545), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_153), .A2(n_255), .B1(n_568), .B2(n_569), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_153), .A2(n_525), .B1(n_604), .B2(n_605), .Y(n_603) );
INVx6_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
O2A1O1Ixp5_ASAP7_75t_L g220 ( .A1(n_154), .A2(n_193), .B(n_221), .C(n_222), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_154), .A2(n_522), .B(n_524), .C(n_528), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_154), .A2(n_559), .B(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_154), .B(n_522), .Y(n_634) );
BUFx8_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
INVx1_ASAP7_75t_L g195 ( .A(n_155), .Y(n_195) );
INVx1_ASAP7_75t_L g580 ( .A(n_155), .Y(n_580) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
INVx4_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g525 ( .A(n_160), .Y(n_525) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g557 ( .A(n_161), .Y(n_557) );
AO31x2_ASAP7_75t_L g172 ( .A1(n_162), .A2(n_173), .A3(n_179), .B(n_181), .Y(n_172) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_162), .A2(n_532), .B(n_540), .Y(n_531) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_SL g198 ( .A(n_164), .B(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_164), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g170 ( .A(n_165), .Y(n_170) );
INVx2_ASAP7_75t_L g197 ( .A(n_165), .Y(n_197) );
OAI21xp33_ASAP7_75t_L g528 ( .A1(n_165), .A2(n_527), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_166), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_170), .B(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g392 ( .A(n_171), .Y(n_392) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g240 ( .A(n_172), .Y(n_240) );
AND2x4_ASAP7_75t_L g281 ( .A(n_172), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g301 ( .A(n_172), .B(n_200), .Y(n_301) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_172), .Y(n_353) );
INVx1_ASAP7_75t_L g446 ( .A(n_172), .Y(n_446) );
AND2x2_ASAP7_75t_L g492 ( .A(n_172), .B(n_185), .Y(n_492) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g203 ( .A(n_176), .Y(n_203) );
OAI22xp33_ASAP7_75t_L g537 ( .A1(n_176), .A2(n_208), .B1(n_538), .B2(n_539), .Y(n_537) );
INVx2_ASAP7_75t_L g570 ( .A(n_178), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_178), .B(n_579), .Y(n_578) );
AO31x2_ASAP7_75t_L g248 ( .A1(n_179), .A2(n_209), .A3(n_249), .B(n_256), .Y(n_248) );
AO31x2_ASAP7_75t_L g566 ( .A1(n_179), .A2(n_196), .A3(n_567), .B(n_571), .Y(n_566) );
INVx2_ASAP7_75t_SL g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_SL g226 ( .A(n_180), .Y(n_226) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_184), .B(n_358), .Y(n_357) );
NAND2x1_ASAP7_75t_L g362 ( .A(n_184), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g486 ( .A(n_184), .B(n_384), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_184), .B(n_440), .Y(n_490) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_200), .Y(n_184) );
INVx4_ASAP7_75t_SL g242 ( .A(n_185), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_185), .B(n_244), .Y(n_294) );
BUFx2_ASAP7_75t_L g378 ( .A(n_185), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_185), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_190), .B(n_535), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g553 ( .A1(n_193), .A2(n_554), .B(n_555), .C(n_556), .Y(n_553) );
INVx1_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g255 ( .A(n_195), .Y(n_255) );
AOI21x1_ASAP7_75t_L g609 ( .A1(n_196), .A2(n_610), .B(n_620), .Y(n_609) );
BUFx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g541 ( .A(n_197), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_197), .B(n_547), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_197), .B(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_197), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g244 ( .A(n_200), .Y(n_244) );
INVx2_ASAP7_75t_L g282 ( .A(n_200), .Y(n_282) );
AND2x2_ASAP7_75t_L g284 ( .A(n_200), .B(n_239), .Y(n_284) );
INVx1_ASAP7_75t_L g309 ( .A(n_200), .Y(n_309) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_200), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_200), .B(n_392), .Y(n_423) );
OAI21xp33_ASAP7_75t_SL g576 ( .A1(n_204), .A2(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
BUFx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_210), .B(n_212), .Y(n_211) );
INVx2_ASAP7_75t_SL g218 ( .A(n_210), .Y(n_218) );
INVx4_ASAP7_75t_L g228 ( .A(n_210), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_210), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_210), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g585 ( .A(n_210), .B(n_563), .Y(n_585) );
INVxp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVxp67_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g467 ( .A(n_215), .B(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_229), .Y(n_215) );
AND2x4_ASAP7_75t_L g262 ( .A(n_216), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g324 ( .A(n_216), .B(n_267), .Y(n_324) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g410 ( .A(n_217), .Y(n_410) );
OAI21x1_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_227), .Y(n_217) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_218), .A2(n_219), .B(n_227), .Y(n_297) );
OAI21x1_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_223), .B(n_226), .Y(n_219) );
INVx2_ASAP7_75t_L g273 ( .A(n_228), .Y(n_273) );
NOR2x1_ASAP7_75t_L g561 ( .A(n_228), .B(n_562), .Y(n_561) );
AND2x4_ASAP7_75t_L g322 ( .A(n_229), .B(n_248), .Y(n_322) );
INVx3_ASAP7_75t_L g345 ( .A(n_229), .Y(n_345) );
INVx2_ASAP7_75t_L g366 ( .A(n_229), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_229), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_229), .B(n_266), .Y(n_460) );
INVx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g247 ( .A(n_230), .B(n_248), .Y(n_247) );
BUFx2_ASAP7_75t_L g261 ( .A(n_230), .Y(n_261) );
AND2x2_ASAP7_75t_L g339 ( .A(n_230), .B(n_263), .Y(n_339) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_241), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx3_ASAP7_75t_L g317 ( .A(n_239), .Y(n_317) );
AND2x2_ASAP7_75t_L g352 ( .A(n_239), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g421 ( .A(n_239), .B(n_242), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_240), .B(n_242), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_241), .B(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g280 ( .A(n_242), .Y(n_280) );
AND2x2_ASAP7_75t_L g308 ( .A(n_242), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g326 ( .A(n_242), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g368 ( .A(n_242), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_242), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g429 ( .A(n_242), .Y(n_429) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_247), .B(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_SL g303 ( .A(n_247), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g382 ( .A(n_247), .B(n_265), .Y(n_382) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_247), .Y(n_417) );
INVx2_ASAP7_75t_L g434 ( .A(n_247), .Y(n_434) );
INVx2_ASAP7_75t_L g263 ( .A(n_248), .Y(n_263) );
OR2x2_ASAP7_75t_L g314 ( .A(n_248), .B(n_305), .Y(n_314) );
INVx1_ASAP7_75t_L g335 ( .A(n_248), .Y(n_335) );
BUFx2_ASAP7_75t_L g350 ( .A(n_248), .Y(n_350) );
OR2x2_ASAP7_75t_L g419 ( .A(n_248), .B(n_268), .Y(n_419) );
INVx2_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_252), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_255), .B(n_537), .Y(n_536) );
AOI21xp5_ASAP7_75t_SL g258 ( .A1(n_259), .A2(n_264), .B(n_277), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g385 ( .A1(n_259), .A2(n_341), .B(n_386), .C(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g285 ( .A(n_260), .B(n_286), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_260), .A2(n_319), .B1(n_485), .B2(n_486), .Y(n_484) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g276 ( .A(n_262), .Y(n_276) );
AND2x4_ASAP7_75t_L g404 ( .A(n_262), .B(n_313), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_262), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_276), .Y(n_264) );
INVx1_ASAP7_75t_L g286 ( .A(n_265), .Y(n_286) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x4_ASAP7_75t_L g304 ( .A(n_266), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_267), .B(n_297), .Y(n_347) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g296 ( .A(n_268), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g313 ( .A(n_268), .Y(n_313) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_268), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_271), .B(n_613), .Y(n_612) );
AO31x2_ASAP7_75t_L g602 ( .A1(n_273), .A2(n_563), .A3(n_603), .B(n_606), .Y(n_602) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
AND2x2_ASAP7_75t_L g299 ( .A(n_279), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_280), .B(n_359), .Y(n_398) );
INVx2_ASAP7_75t_L g290 ( .A(n_281), .Y(n_290) );
AND2x2_ASAP7_75t_L g367 ( .A(n_281), .B(n_368), .Y(n_367) );
NAND2x1p5_ASAP7_75t_L g412 ( .A(n_281), .B(n_331), .Y(n_412) );
AND2x2_ASAP7_75t_L g449 ( .A(n_281), .B(n_421), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B(n_287), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_295), .B1(n_298), .B2(n_302), .Y(n_287) );
NOR2x1_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g493 ( .A(n_290), .Y(n_493) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g333 ( .A(n_296), .Y(n_333) );
AND2x2_ASAP7_75t_L g360 ( .A(n_296), .B(n_345), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_296), .B(n_339), .Y(n_430) );
AND2x4_ASAP7_75t_L g476 ( .A(n_296), .B(n_322), .Y(n_476) );
INVx1_ASAP7_75t_L g305 ( .A(n_297), .Y(n_305) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_L g482 ( .A(n_300), .B(n_378), .Y(n_482) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g415 ( .A(n_301), .B(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g443 ( .A(n_301), .B(n_317), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_302), .B(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g424 ( .A(n_304), .B(n_425), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_311), .B1(n_315), .B2(n_319), .C(n_325), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_L g341 ( .A(n_308), .Y(n_341) );
AND2x2_ASAP7_75t_L g465 ( .A(n_308), .B(n_331), .Y(n_465) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_309), .Y(n_329) );
INVx3_ASAP7_75t_L g327 ( .A(n_310), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_310), .B(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g399 ( .A(n_310), .B(n_400), .Y(n_399) );
NOR2xp67_ASAP7_75t_SL g311 ( .A(n_312), .B(n_314), .Y(n_311) );
AND2x2_ASAP7_75t_L g338 ( .A(n_312), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_312), .B(n_345), .Y(n_407) );
AOI322xp5_ASAP7_75t_L g413 ( .A1(n_312), .A2(n_399), .A3(n_414), .B1(n_417), .B2(n_418), .C1(n_420), .C2(n_424), .Y(n_413) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g355 ( .A(n_313), .B(n_322), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_314), .B(n_366), .Y(n_365) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_314), .B(n_464), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_315), .A2(n_457), .B1(n_461), .B2(n_465), .Y(n_456) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx4_ASAP7_75t_L g440 ( .A(n_317), .Y(n_440) );
OR2x2_ASAP7_75t_L g470 ( .A(n_317), .B(n_445), .Y(n_470) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g483 ( .A(n_322), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_323), .B(n_349), .Y(n_370) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI211x1_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B(n_333), .C(n_334), .Y(n_325) );
INVx2_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g390 ( .A(n_331), .Y(n_390) );
NAND2x1_ASAP7_75t_L g481 ( .A(n_331), .B(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g387 ( .A(n_332), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g452 ( .A(n_334), .Y(n_452) );
BUFx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_354), .C(n_369), .Y(n_336) );
OAI211xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B(n_342), .C(n_352), .Y(n_337) );
INVx1_ASAP7_75t_L g351 ( .A(n_338), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_339), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g409 ( .A(n_339), .B(n_410), .Y(n_409) );
NAND2xp33_ASAP7_75t_L g432 ( .A(n_339), .B(n_380), .Y(n_432) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_351), .Y(n_342) );
INVx1_ASAP7_75t_L g478 ( .A(n_343), .Y(n_478) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_344), .B(n_348), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx2_ASAP7_75t_L g425 ( .A(n_345), .Y(n_425) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g380 ( .A(n_347), .Y(n_380) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_347), .Y(n_455) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_360), .B2(n_361), .C(n_364), .Y(n_354) );
INVxp67_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g416 ( .A(n_359), .Y(n_416) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g402 ( .A(n_366), .Y(n_402) );
NOR2x1p5_ASAP7_75t_L g418 ( .A(n_366), .B(n_419), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_367), .A2(n_406), .B(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g374 ( .A(n_368), .Y(n_374) );
AOI211xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B(n_375), .C(n_385), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .B1(n_381), .B2(n_383), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g464 ( .A(n_388), .Y(n_464) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
NOR3xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_426), .C(n_447), .Y(n_393) );
NAND3xp33_ASAP7_75t_SL g394 ( .A(n_395), .B(n_405), .C(n_413), .Y(n_394) );
OAI21xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_399), .B(n_401), .Y(n_395) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
AND2x2_ASAP7_75t_L g495 ( .A(n_402), .B(n_463), .Y(n_495) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g441 ( .A1(n_404), .A2(n_442), .B(n_444), .Y(n_441) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
OR2x2_ASAP7_75t_L g433 ( .A(n_410), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g468 ( .A(n_419), .Y(n_468) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_422), .Y(n_485) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g428 ( .A(n_423), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g438 ( .A(n_423), .Y(n_438) );
OAI221xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_430), .B1(n_431), .B2(n_435), .C(n_441), .Y(n_426) );
OAI21xp5_ASAP7_75t_L g472 ( .A1(n_427), .A2(n_473), .B(n_477), .Y(n_472) );
BUFx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI32xp33_ASAP7_75t_L g466 ( .A1(n_429), .A2(n_440), .A3(n_467), .B1(n_468), .B2(n_469), .Y(n_466) );
AND2x2_ASAP7_75t_SL g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_442), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI211xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_450), .B(n_456), .C(n_466), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NOR3xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_479), .C(n_487), .Y(n_471) );
INVxp33_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI21xp33_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_483), .B(n_484), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_491), .B(n_494), .Y(n_487) );
INVxp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_SL g491 ( .A(n_492), .B(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_496), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx12f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_507), .B(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g867 ( .A(n_507), .Y(n_867) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_850), .B(n_855), .C(n_863), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g855 ( .A1(n_509), .A2(n_852), .B(n_856), .Y(n_855) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx8_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g860 ( .A(n_512), .B(n_861), .Y(n_860) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_747), .Y(n_513) );
AND3x1_ASAP7_75t_L g514 ( .A(n_515), .B(n_665), .C(n_724), .Y(n_514) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_564), .B1(n_586), .B2(n_637), .C(n_640), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_548), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .Y(n_518) );
INVx2_ASAP7_75t_L g597 ( .A(n_519), .Y(n_597) );
AND2x2_ASAP7_75t_L g652 ( .A(n_519), .B(n_596), .Y(n_652) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g745 ( .A(n_520), .B(n_680), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_520), .B(n_542), .Y(n_809) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g633 ( .A(n_524), .Y(n_633) );
OAI21x1_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B(n_527), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_525), .A2(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g635 ( .A(n_528), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_529), .A2(n_611), .B(n_617), .Y(n_610) );
INVx2_ASAP7_75t_L g684 ( .A(n_530), .Y(n_684) );
OR2x2_ASAP7_75t_L g773 ( .A(n_530), .B(n_690), .Y(n_773) );
OR2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_542), .Y(n_530) );
INVx1_ASAP7_75t_L g590 ( .A(n_531), .Y(n_590) );
INVx2_ASAP7_75t_L g675 ( .A(n_531), .Y(n_675) );
AND2x2_ASAP7_75t_L g699 ( .A(n_531), .B(n_542), .Y(n_699) );
AND2x4_ASAP7_75t_L g712 ( .A(n_531), .B(n_632), .Y(n_712) );
AND2x2_ASAP7_75t_L g729 ( .A(n_531), .B(n_593), .Y(n_729) );
AND2x2_ASAP7_75t_L g739 ( .A(n_531), .B(n_631), .Y(n_739) );
AND2x2_ASAP7_75t_L g767 ( .A(n_531), .B(n_550), .Y(n_767) );
INVx2_ASAP7_75t_L g596 ( .A(n_542), .Y(n_596) );
AND2x2_ASAP7_75t_L g636 ( .A(n_542), .B(n_550), .Y(n_636) );
INVx2_ASAP7_75t_L g680 ( .A(n_542), .Y(n_680) );
AND2x2_ASAP7_75t_L g812 ( .A(n_542), .B(n_675), .Y(n_812) );
AND3x1_ASAP7_75t_L g648 ( .A(n_548), .B(n_590), .C(n_649), .Y(n_648) );
NAND2x1p5_ASAP7_75t_L g664 ( .A(n_548), .B(n_652), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_548), .B(n_812), .Y(n_829) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx2_ASAP7_75t_L g733 ( .A(n_549), .Y(n_733) );
AND2x2_ASAP7_75t_L g842 ( .A(n_549), .B(n_624), .Y(n_842) );
BUFx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g593 ( .A(n_550), .Y(n_593) );
AND2x2_ASAP7_75t_L g595 ( .A(n_550), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g681 ( .A(n_550), .Y(n_681) );
NAND2x1p5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
OAI21x1_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_558), .B(n_561), .Y(n_552) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g708 ( .A(n_565), .B(n_709), .Y(n_708) );
AND2x4_ASAP7_75t_L g815 ( .A(n_565), .B(n_705), .Y(n_815) );
AND2x2_ASAP7_75t_L g822 ( .A(n_565), .B(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_573), .Y(n_565) );
INVx1_ASAP7_75t_L g639 ( .A(n_566), .Y(n_639) );
INVx1_ASAP7_75t_L g657 ( .A(n_566), .Y(n_657) );
OR2x2_ASAP7_75t_L g661 ( .A(n_566), .B(n_602), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_566), .B(n_602), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_566), .B(n_626), .Y(n_687) );
INVx1_ASAP7_75t_L g759 ( .A(n_566), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_566), .B(n_608), .Y(n_818) );
OR2x2_ASAP7_75t_L g656 ( .A(n_573), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_573), .B(n_624), .Y(n_663) );
INVx3_ASAP7_75t_L g671 ( .A(n_573), .Y(n_671) );
NAND2x1p5_ASAP7_75t_SL g696 ( .A(n_573), .B(n_670), .Y(n_696) );
BUFx2_ASAP7_75t_L g718 ( .A(n_573), .Y(n_718) );
INVx1_ASAP7_75t_L g723 ( .A(n_573), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_573), .B(n_759), .Y(n_776) );
AND2x4_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_582), .B(n_585), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
BUFx4f_ASAP7_75t_L g616 ( .A(n_580), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_621), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_594), .B(n_598), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g654 ( .A(n_590), .Y(n_654) );
INVx1_ASAP7_75t_L g746 ( .A(n_590), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_591), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g782 ( .A(n_591), .B(n_699), .Y(n_782) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g794 ( .A(n_592), .B(n_712), .Y(n_794) );
BUFx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g698 ( .A(n_593), .B(n_631), .Y(n_698) );
AND2x2_ASAP7_75t_L g738 ( .A(n_593), .B(n_680), .Y(n_738) );
AND2x4_ASAP7_75t_SL g594 ( .A(n_595), .B(n_597), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_595), .B(n_674), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_595), .B(n_712), .Y(n_721) );
AND2x2_ASAP7_75t_L g761 ( .A(n_595), .B(n_754), .Y(n_761) );
INVx1_ASAP7_75t_L g778 ( .A(n_596), .Y(n_778) );
OAI322xp33_ASAP7_75t_L g640 ( .A1(n_597), .A2(n_641), .A3(n_647), .B1(n_650), .B2(n_655), .C1(n_659), .C2(n_664), .Y(n_640) );
AOI32xp33_ASAP7_75t_L g731 ( .A1(n_597), .A2(n_691), .A3(n_732), .B1(n_734), .B2(n_736), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_597), .B(n_800), .Y(n_799) );
AND2x2_ASAP7_75t_L g819 ( .A(n_597), .B(n_738), .Y(n_819) );
INVxp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g658 ( .A(n_601), .Y(n_658) );
AND2x2_ASAP7_75t_L g722 ( .A(n_601), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g796 ( .A(n_601), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_601), .B(n_758), .Y(n_797) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_608), .Y(n_601) );
INVx2_ASAP7_75t_SL g626 ( .A(n_602), .Y(n_626) );
BUFx2_ASAP7_75t_L g644 ( .A(n_602), .Y(n_644) );
INVx2_ASAP7_75t_L g670 ( .A(n_608), .Y(n_670) );
OR2x2_ASAP7_75t_L g706 ( .A(n_608), .B(n_626), .Y(n_706) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g624 ( .A(n_609), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_614), .B(n_616), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_627), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g823 ( .A(n_623), .Y(n_823) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_624), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_624), .B(n_671), .Y(n_686) );
INVxp67_ASAP7_75t_L g693 ( .A(n_624), .Y(n_693) );
OR2x2_ASAP7_75t_L g763 ( .A(n_625), .B(n_670), .Y(n_763) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_636), .Y(n_628) );
AND2x2_ASAP7_75t_L g683 ( .A(n_629), .B(n_684), .Y(n_683) );
NOR2x1_ASAP7_75t_L g846 ( .A(n_629), .B(n_681), .Y(n_846) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g754 ( .A(n_630), .Y(n_754) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g674 ( .A(n_631), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g779 ( .A(n_632), .B(n_675), .Y(n_779) );
AOI21x1_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_635), .Y(n_632) );
INVx2_ASAP7_75t_L g715 ( .A(n_636), .Y(n_715) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g646 ( .A(n_639), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_645), .Y(n_641) );
INVx1_ASAP7_75t_L g719 ( .A(n_642), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_642), .B(n_758), .Y(n_827) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_643), .B(n_776), .Y(n_775) );
AND2x4_ASAP7_75t_L g786 ( .A(n_643), .B(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g695 ( .A(n_646), .B(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_646), .B(n_704), .Y(n_703) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g691 ( .A(n_656), .Y(n_691) );
INVx1_ASAP7_75t_L g787 ( .A(n_656), .Y(n_787) );
INVx1_ASAP7_75t_L g837 ( .A(n_656), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_660), .B(n_710), .Y(n_742) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g727 ( .A(n_661), .Y(n_727) );
OR2x2_ASAP7_75t_L g735 ( .A(n_661), .B(n_696), .Y(n_735) );
OR2x2_ASAP7_75t_L g803 ( .A(n_661), .B(n_710), .Y(n_803) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g751 ( .A(n_663), .B(n_668), .Y(n_751) );
INVx1_ASAP7_75t_L g834 ( .A(n_664), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_700), .Y(n_665) );
OAI321xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_672), .A3(n_676), .B1(n_682), .B2(n_685), .C(n_688), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_667), .B(n_773), .Y(n_772) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g710 ( .A(n_670), .Y(n_710) );
AND2x4_ASAP7_75t_L g758 ( .A(n_671), .B(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g762 ( .A(n_671), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_673), .B(n_841), .Y(n_840) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI211xp5_ASAP7_75t_L g768 ( .A1(n_677), .A2(n_769), .B(n_772), .C(n_774), .Y(n_768) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g766 ( .A(n_679), .Y(n_766) );
INVx1_ASAP7_75t_L g800 ( .A(n_679), .Y(n_800) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g690 ( .A(n_681), .Y(n_690) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g689 ( .A(n_684), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_685), .B(n_751), .Y(n_750) );
OR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_686), .Y(n_790) );
AOI32xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .A3(n_692), .B1(n_694), .B2(n_697), .Y(n_688) );
OR2x2_ASAP7_75t_L g844 ( .A(n_690), .B(n_745), .Y(n_844) );
AND2x2_ASAP7_75t_L g725 ( .A(n_692), .B(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g770 ( .A(n_693), .B(n_771), .Y(n_770) );
NAND2x1_ASAP7_75t_L g836 ( .A(n_693), .B(n_837), .Y(n_836) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
AND2x2_ASAP7_75t_L g816 ( .A(n_698), .B(n_812), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_699), .B(n_754), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_699), .A2(n_726), .B1(n_822), .B2(n_824), .Y(n_821) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B1(n_707), .B2(n_711), .C(n_713), .Y(n_700) );
INVxp67_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g757 ( .A(n_705), .B(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g847 ( .A(n_709), .B(n_726), .Y(n_847) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx3_ASAP7_75t_L g717 ( .A(n_712), .Y(n_717) );
AND2x2_ASAP7_75t_L g824 ( .A(n_712), .B(n_766), .Y(n_824) );
AOI32xp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_718), .A3(n_719), .B1(n_720), .B2(n_722), .Y(n_713) );
NOR2xp33_ASAP7_75t_SL g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x4_ASAP7_75t_L g726 ( .A(n_723), .B(n_727), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_728), .B(n_730), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g740 ( .A1(n_726), .A2(n_741), .B(n_743), .Y(n_740) );
OAI21xp33_ASAP7_75t_L g839 ( .A1(n_726), .A2(n_840), .B(n_843), .Y(n_839) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_740), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
AND2x2_ASAP7_75t_L g838 ( .A(n_739), .B(n_800), .Y(n_838) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx3_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
NOR4xp75_ASAP7_75t_L g747 ( .A(n_748), .B(n_780), .C(n_804), .D(n_830), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_768), .Y(n_748) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_752), .B(n_755), .Y(n_749) );
INVx2_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
OAI22xp33_ASAP7_75t_L g792 ( .A1(n_753), .A2(n_793), .B1(n_795), .B2(n_797), .Y(n_792) );
OAI22xp33_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_760), .B1(n_762), .B2(n_764), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_756), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g771 ( .A(n_758), .Y(n_771) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
OAI21xp33_ASAP7_75t_L g845 ( .A1(n_765), .A2(n_846), .B(n_847), .Y(n_845) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AOI21xp33_ASAP7_75t_L g798 ( .A1(n_773), .A2(n_799), .B(n_801), .Y(n_798) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_777), .Y(n_774) );
OR2x2_ASAP7_75t_L g795 ( .A(n_776), .B(n_796), .Y(n_795) );
BUFx2_ASAP7_75t_L g791 ( .A(n_777), .Y(n_791) );
AND2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
OAI21xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_783), .B(n_788), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVxp67_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
AOI211xp5_ASAP7_75t_SL g788 ( .A1(n_789), .A2(n_791), .B(n_792), .C(n_798), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVxp67_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g813 ( .A(n_795), .Y(n_813) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND2x1_ASAP7_75t_SL g804 ( .A(n_805), .B(n_820), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_814), .Y(n_805) );
OAI21xp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_810), .B(n_813), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B1(n_817), .B2(n_819), .Y(n_814) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
AND2x2_ASAP7_75t_L g820 ( .A(n_821), .B(n_825), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_822), .A2(n_834), .B1(n_835), .B2(n_838), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_826), .B(n_828), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_845), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_839), .Y(n_832) );
INVxp67_ASAP7_75t_SL g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_SL g863 ( .A(n_856), .B(n_864), .Y(n_863) );
BUFx10_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g869 ( .A(n_862), .Y(n_869) );
INVx1_ASAP7_75t_SL g864 ( .A(n_865), .Y(n_864) );
BUFx12f_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
AND2x6_ASAP7_75t_SL g866 ( .A(n_867), .B(n_868), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_871), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_872), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g872 ( .A(n_873), .Y(n_872) );
endmodule