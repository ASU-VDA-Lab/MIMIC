module fake_jpeg_3184_n_388 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_388);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_388;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_26),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

NAND2x1_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_0),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_52),
.B(n_85),
.Y(n_143)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_26),
.B(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_68),
.B(n_92),
.Y(n_127)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_SL g74 ( 
.A1(n_25),
.A2(n_1),
.B(n_2),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_74),
.A2(n_16),
.B(n_42),
.Y(n_121)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_83),
.B(n_84),
.Y(n_146)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_89),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_90),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_35),
.B(n_2),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_91),
.B(n_24),
.Y(n_148)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_93),
.B(n_94),
.Y(n_136)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_95),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_32),
.B1(n_24),
.B2(n_43),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_96),
.A2(n_97),
.B1(n_112),
.B2(n_29),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_16),
.B1(n_43),
.B2(n_42),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_72),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_16),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_67),
.Y(n_153)
);

CKINVDCx12_ASAP7_75t_R g120 ( 
.A(n_80),
.Y(n_120)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_121),
.B(n_144),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_79),
.A2(n_35),
.B(n_22),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_46),
.B1(n_31),
.B2(n_47),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_130),
.A2(n_44),
.B1(n_41),
.B2(n_20),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_48),
.A2(n_47),
.B1(n_28),
.B2(n_32),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_139),
.A2(n_27),
.B1(n_47),
.B2(n_63),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_88),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_141),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_90),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_95),
.B(n_28),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_55),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_56),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_148),
.B(n_27),
.Y(n_154)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_151),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_152),
.A2(n_162),
.B1(n_178),
.B2(n_168),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_153),
.B(n_165),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_154),
.B(n_158),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_155),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_108),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_161),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_66),
.B1(n_59),
.B2(n_19),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_164),
.A2(n_175),
.B1(n_188),
.B2(n_122),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_2),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_124),
.A2(n_46),
.B1(n_31),
.B2(n_29),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_168),
.A2(n_130),
.B(n_128),
.C(n_137),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_114),
.B(n_3),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_169),
.B(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_105),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_171),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_174),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_143),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_46),
.B1(n_31),
.B2(n_29),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_186),
.Y(n_217)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_22),
.B1(n_19),
.B2(n_44),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_101),
.A2(n_22),
.B1(n_19),
.B2(n_44),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_174),
.B1(n_117),
.B2(n_156),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_102),
.B(n_3),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_184),
.B(n_187),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_97),
.A2(n_22),
.B1(n_19),
.B2(n_41),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_102),
.B(n_4),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_129),
.A2(n_22),
.B1(n_19),
.B2(n_41),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_103),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_189),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_110),
.B(n_22),
.C(n_5),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_191),
.A3(n_169),
.B1(n_153),
.B2(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_107),
.B(n_4),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_170),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_195),
.A2(n_203),
.B1(n_171),
.B2(n_176),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_156),
.A2(n_147),
.B1(n_104),
.B2(n_131),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_198),
.A2(n_202),
.B1(n_209),
.B2(n_178),
.Y(n_232)
);

AOI32xp33_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_111),
.A3(n_137),
.B1(n_122),
.B2(n_98),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_200),
.B(n_111),
.Y(n_252)
);

NOR2x1_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_224),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_164),
.A2(n_107),
.B1(n_118),
.B2(n_133),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_116),
.B1(n_123),
.B2(n_142),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_150),
.A2(n_133),
.B1(n_118),
.B2(n_146),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_223),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_162),
.A2(n_146),
.B(n_103),
.C(n_105),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_219),
.B(n_109),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_168),
.A2(n_98),
.B(n_117),
.C(n_109),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_227),
.Y(n_229)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_216),
.A2(n_191),
.B1(n_187),
.B2(n_184),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_230),
.A2(n_237),
.B1(n_197),
.B2(n_219),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_234),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g283 ( 
.A1(n_232),
.A2(n_258),
.B(n_212),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_190),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_236),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_217),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_163),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_221),
.A2(n_152),
.B1(n_142),
.B2(n_134),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_247),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_183),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_177),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_241),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_242),
.A2(n_252),
.B(n_199),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_159),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_257),
.C(n_220),
.Y(n_279)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

INVx13_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_226),
.B(n_167),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_250),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_213),
.B(n_116),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_249),
.Y(n_286)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_186),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_193),
.B(n_161),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_217),
.Y(n_273)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_253),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_180),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_254),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_255),
.Y(n_266)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_256),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_197),
.B(n_209),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_211),
.A2(n_151),
.B1(n_157),
.B2(n_134),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_251),
.B1(n_229),
.B2(n_231),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_260),
.A2(n_264),
.B1(n_272),
.B2(n_258),
.Y(n_300)
);

AND2x6_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_200),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_267),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_198),
.B1(n_202),
.B2(n_219),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_246),
.A2(n_201),
.B1(n_227),
.B2(n_222),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_271),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_232),
.A2(n_201),
.B1(n_227),
.B2(n_222),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_229),
.A2(n_196),
.B1(n_160),
.B2(n_182),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_273),
.B(n_207),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_274),
.A2(n_283),
.B(n_256),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_250),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_280),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_279),
.B(n_253),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_240),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_205),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_215),
.B(n_237),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_230),
.A2(n_196),
.B1(n_214),
.B2(n_199),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_282),
.A2(n_228),
.B1(n_238),
.B2(n_249),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_276),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_292),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_233),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_289),
.C(n_290),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_243),
.C(n_257),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_245),
.C(n_234),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_276),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_294),
.B(n_298),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_236),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_295),
.B(n_259),
.Y(n_331)
);

AOI221xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_247),
.B1(n_254),
.B2(n_241),
.C(n_239),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_296),
.A2(n_300),
.B1(n_264),
.B2(n_263),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_299),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_301),
.A2(n_303),
.B(n_281),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_310),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_268),
.A2(n_215),
.B(n_255),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_265),
.B(n_255),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_306),
.C(n_307),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_273),
.A2(n_214),
.B1(n_218),
.B2(n_166),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_286),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_210),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_210),
.C(n_207),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_308),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_294),
.B(n_268),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_212),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_297),
.A2(n_267),
.B1(n_264),
.B2(n_262),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_315),
.A2(n_317),
.B1(n_319),
.B2(n_323),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_318),
.Y(n_343)
);

OA22x2_ASAP7_75t_L g318 ( 
.A1(n_297),
.A2(n_301),
.B1(n_300),
.B2(n_309),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_291),
.A2(n_262),
.B1(n_282),
.B2(n_275),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_293),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_331),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_290),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_326),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_287),
.A2(n_286),
.B1(n_272),
.B2(n_284),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_302),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_284),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_311),
.Y(n_344)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

FAx1_ASAP7_75t_SL g332 ( 
.A(n_313),
.B(n_292),
.CI(n_293),
.CON(n_332),
.SN(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_304),
.C(n_307),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_336),
.C(n_340),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_325),
.C(n_312),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_315),
.A2(n_310),
.B1(n_271),
.B2(n_305),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_346),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_274),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_341),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_325),
.B(n_298),
.C(n_303),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_283),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_320),
.C(n_319),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_336),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_283),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_345),
.B(n_318),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_L g346 ( 
.A1(n_314),
.A2(n_277),
.B1(n_270),
.B2(n_278),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_353),
.Y(n_356)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_335),
.Y(n_350)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_350),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_343),
.A2(n_316),
.B(n_314),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_351),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_333),
.A2(n_327),
.B(n_328),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_354),
.B(n_332),
.C(n_330),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_327),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_324),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_342),
.C(n_344),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_358),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_341),
.C(n_339),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_360),
.B(n_347),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_362),
.B(n_352),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_359),
.A2(n_352),
.B1(n_351),
.B2(n_348),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_364),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_361),
.B(n_354),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_365),
.A2(n_371),
.B(n_10),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_366),
.B(n_149),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_359),
.A2(n_285),
.B(n_266),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_368),
.A2(n_5),
.B(n_8),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_362),
.A2(n_214),
.B1(n_285),
.B2(n_212),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_356),
.A2(n_285),
.B1(n_131),
.B2(n_99),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_358),
.A2(n_192),
.B(n_99),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_149),
.C(n_125),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_374),
.B(n_376),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_366),
.B(n_10),
.C(n_12),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_375),
.B(n_370),
.C(n_369),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_379),
.A2(n_380),
.B(n_381),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_372),
.B(n_14),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_377),
.B(n_10),
.C(n_13),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_378),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_382),
.A2(n_383),
.B(n_13),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_373),
.C(n_374),
.Y(n_383)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_385),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_384),
.Y(n_387)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_387),
.Y(n_388)
);


endmodule