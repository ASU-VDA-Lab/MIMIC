module fake_jpeg_22845_n_206 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_22),
.Y(n_37)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_35),
.B1(n_23),
.B2(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_27),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_23),
.B1(n_24),
.B2(n_15),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_33),
.B1(n_35),
.B2(n_34),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_15),
.B1(n_23),
.B2(n_24),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_47),
.B1(n_49),
.B2(n_13),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_45),
.B1(n_27),
.B2(n_29),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_32),
.C(n_36),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_28),
.C(n_36),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_16),
.B1(n_21),
.B2(n_17),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_26),
.B1(n_17),
.B2(n_21),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_50),
.B(n_52),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_46),
.B1(n_38),
.B2(n_32),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_52),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_43),
.C(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_36),
.B(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_67),
.B1(n_69),
.B2(n_38),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_66),
.B1(n_42),
.B2(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_65),
.Y(n_78)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_39),
.A2(n_29),
.B1(n_27),
.B2(n_32),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_29),
.B(n_27),
.C(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_29),
.B1(n_13),
.B2(n_14),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_85),
.B1(n_53),
.B2(n_38),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_43),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_73),
.Y(n_99)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_61),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_84),
.B1(n_66),
.B2(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_86),
.Y(n_100)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_59),
.B1(n_69),
.B2(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_101),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_90),
.B(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_54),
.Y(n_91)
);

BUFx24_ASAP7_75t_SL g92 ( 
.A(n_81),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_67),
.B(n_60),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_93),
.A2(n_98),
.B(n_31),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_87),
.B1(n_83),
.B2(n_46),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_14),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_85),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_108),
.B(n_99),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_73),
.B(n_71),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_114),
.B1(n_91),
.B2(n_105),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_113),
.Y(n_131)
);

NOR3xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_83),
.C(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_90),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_75),
.B1(n_70),
.B2(n_82),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_88),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_70),
.B1(n_65),
.B2(n_79),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_88),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_44),
.B1(n_51),
.B2(n_22),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_125),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_115),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_89),
.C(n_101),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_118),
.A3(n_121),
.B1(n_117),
.B2(n_113),
.C1(n_106),
.C2(n_111),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_128),
.B1(n_130),
.B2(n_133),
.Y(n_141)
);

OA21x2_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_99),
.B(n_94),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_137),
.Y(n_144)
);

OAI22x1_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_99),
.B1(n_51),
.B2(n_44),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_19),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_99),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_20),
.B(n_19),
.C(n_25),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_138),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_140),
.B1(n_109),
.B2(n_119),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_110),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_133),
.A2(n_120),
.B1(n_107),
.B2(n_122),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_124),
.B1(n_134),
.B2(n_135),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_106),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_150),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_106),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_121),
.C(n_119),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_153),
.C(n_155),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_51),
.C(n_31),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_51),
.C(n_31),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_142),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_165),
.Y(n_175)
);

AOI321xp33_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_130),
.A3(n_132),
.B1(n_140),
.B2(n_139),
.C(n_131),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_SL g168 ( 
.A(n_162),
.B(n_167),
.C(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_44),
.C(n_138),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_153),
.C(n_143),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_44),
.B1(n_25),
.B2(n_22),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_166),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_169),
.C(n_178),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_144),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_5),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_163),
.B(n_151),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_172),
.B(n_5),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_154),
.C(n_145),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_178),
.C(n_164),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_123),
.Y(n_177)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_7),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_183),
.C(n_187),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_166),
.B1(n_159),
.B2(n_162),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_10),
.B1(n_12),
.B2(n_3),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_176),
.B(n_8),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_182),
.B(n_186),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_8),
.C(n_11),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_9),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_175),
.C(n_171),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_188),
.B(n_10),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_187),
.A2(n_170),
.B(n_2),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_191),
.B(n_12),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_184),
.A2(n_9),
.B(n_11),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_9),
.C(n_11),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_194),
.C(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

AOI21x1_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_197),
.B(n_198),
.Y(n_202)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_12),
.C(n_2),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_190),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_192),
.C(n_2),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_202),
.B1(n_1),
.B2(n_4),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_1),
.C(n_4),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_204),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_4),
.Y(n_206)
);


endmodule