module fake_netlist_1_7810_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx2_ASAP7_75t_SL g11 ( .A(n_10), .Y(n_11) );
NOR2xp33_ASAP7_75t_R g12 ( .A(n_9), .B(n_8), .Y(n_12) );
NAND3xp33_ASAP7_75t_L g13 ( .A(n_1), .B(n_6), .C(n_7), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_2), .B(n_6), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
A2O1A1Ixp33_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_0), .B(n_1), .C(n_2), .Y(n_19) );
AOI22xp33_ASAP7_75t_L g20 ( .A1(n_16), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_11), .A2(n_3), .B(n_4), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_14), .B(n_4), .Y(n_22) );
NAND3xp33_ASAP7_75t_SL g23 ( .A(n_20), .B(n_12), .C(n_15), .Y(n_23) );
XOR2x2_ASAP7_75t_SL g24 ( .A(n_22), .B(n_15), .Y(n_24) );
INVxp67_ASAP7_75t_L g25 ( .A(n_18), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_21), .A2(n_17), .B1(n_11), .B2(n_13), .Y(n_26) );
NOR2x1_ASAP7_75t_L g27 ( .A(n_23), .B(n_19), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_20), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_26), .B(n_17), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
OAI221xp5_ASAP7_75t_L g31 ( .A1(n_27), .A2(n_23), .B1(n_24), .B2(n_13), .C(n_12), .Y(n_31) );
NAND3xp33_ASAP7_75t_SL g32 ( .A(n_31), .B(n_28), .C(n_24), .Y(n_32) );
OAI22xp5_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_28), .B1(n_4), .B2(n_7), .Y(n_33) );
BUFx2_ASAP7_75t_L g34 ( .A(n_33), .Y(n_34) );
BUFx2_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
AOI22x1_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_5), .B1(n_10), .B2(n_36), .Y(n_37) );
AOI22xp33_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_34), .B1(n_35), .B2(n_32), .Y(n_38) );
endmodule