module fake_jpeg_2997_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_12),
.B(n_3),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_27),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_3),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_18),
.B1(n_10),
.B2(n_15),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_22),
.B(n_21),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_11),
.B(n_19),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_9),
.B(n_25),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_15),
.B1(n_13),
.B2(n_19),
.Y(n_32)
);

OA21x2_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_23),
.B(n_6),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_16),
.B1(n_9),
.B2(n_7),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_23),
.B1(n_6),
.B2(n_7),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_25),
.B1(n_20),
.B2(n_27),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_48),
.B1(n_33),
.B2(n_32),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_45),
.B1(n_46),
.B2(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_50),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_5),
.B1(n_23),
.B2(n_37),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_45),
.B(n_48),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_42),
.B(n_45),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_32),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_56),
.B(n_63),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.Y(n_71)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

AOI322xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_66),
.A3(n_60),
.B1(n_54),
.B2(n_38),
.C1(n_57),
.C2(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_74),
.Y(n_75)
);

AOI21x1_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_57),
.B(n_60),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_38),
.B1(n_47),
.B2(n_50),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_34),
.Y(n_78)
);


endmodule