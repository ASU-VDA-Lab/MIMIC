module real_jpeg_15534_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_23),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_1),
.Y(n_147)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_1),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g367 ( 
.A(n_1),
.Y(n_367)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_1),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_2),
.A2(n_10),
.B1(n_150),
.B2(n_154),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_2),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_2),
.B(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_2),
.B(n_296),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_2),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_2),
.B(n_78),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_2),
.B(n_425),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_2),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_2),
.B(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_3),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g372 ( 
.A(n_3),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_4),
.B(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_4),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_4),
.B(n_167),
.Y(n_166)
);

AND2x4_ASAP7_75t_SL g181 ( 
.A(n_4),
.B(n_177),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_4),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_4),
.B(n_237),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_4),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_4),
.B(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_5),
.A2(n_20),
.B(n_22),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_31),
.Y(n_30)
);

AND2x4_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_6),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_6),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g204 ( 
.A(n_6),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_6),
.B(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_7),
.Y(n_119)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_7),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_7),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_7),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_8),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_8),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_8),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_8),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_8),
.B(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_8),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_8),
.B(n_339),
.Y(n_338)
);

NAND2x1_ASAP7_75t_L g137 ( 
.A(n_9),
.B(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_9),
.Y(n_159)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_9),
.B(n_78),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g188 ( 
.A(n_9),
.B(n_184),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_9),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_9),
.B(n_177),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_9),
.B(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_9),
.B(n_440),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_10),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_10),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_10),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_10),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_10),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_10),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_10),
.B(n_334),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_10),
.Y(n_379)
);

BUFx4f_ASAP7_75t_L g143 ( 
.A(n_11),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_11),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_11),
.Y(n_202)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_11),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_12),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_12),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_12),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_12),
.B(n_223),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_12),
.B(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_12),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_12),
.B(n_240),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_12),
.B(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_13),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_13),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_13),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_14),
.Y(n_238)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_14),
.Y(n_304)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_14),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_15),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_15),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_15),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_15),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_15),
.B(n_301),
.Y(n_467)
);

BUFx2_ASAP7_75t_R g487 ( 
.A(n_15),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_16),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_17),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_17),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_17),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_17),
.B(n_174),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_17),
.B(n_301),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_17),
.B(n_150),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_17),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_17),
.B(n_455),
.Y(n_454)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_18),
.Y(n_175)
);

BUFx8_ASAP7_75t_L g214 ( 
.A(n_18),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_569),
.B(n_577),
.C(n_579),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_126),
.B(n_568),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2x1_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_79),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_27),
.B(n_79),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_59),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_48),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_29),
.B(n_48),
.C(n_59),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_35),
.C(n_41),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_30),
.A2(n_35),
.B1(n_53),
.B2(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_SL g571 ( 
.A(n_30),
.B(n_50),
.C(n_55),
.Y(n_571)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_33),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_34),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_35),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_69),
.C(n_76),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_35),
.A2(n_63),
.B1(n_76),
.B2(n_77),
.Y(n_121)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_50),
.A2(n_54),
.B1(n_573),
.B2(n_577),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_116),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_52),
.B(n_199),
.Y(n_198)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.C(n_68),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_60),
.A2(n_61),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_64),
.B(n_68),
.Y(n_125)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2x2_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_76),
.A2(n_77),
.B1(n_115),
.B2(n_327),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_111),
.C(n_115),
.Y(n_110)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_78),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_122),
.C(n_123),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_80),
.B(n_543),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_110),
.C(n_120),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_81),
.B(n_541),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_99),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_100),
.C(n_104),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_89),
.C(n_95),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_83),
.A2(n_84),
.B1(n_89),
.B2(n_90),
.Y(n_532)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_88),
.Y(n_395)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2x1_ASAP7_75t_L g531 ( 
.A(n_95),
.B(n_532),
.Y(n_531)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_103),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_109),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_109),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_110),
.B(n_120),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_SL g535 ( 
.A(n_111),
.B(n_536),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_115),
.A2(n_198),
.B1(n_208),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_115),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_115),
.B(n_208),
.C(n_318),
.Y(n_537)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_122),
.B(n_123),
.Y(n_543)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI21x1_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_525),
.B(n_563),
.Y(n_126)
);

AO21x2_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_356),
.B(n_522),
.Y(n_127)
);

NOR2xp67_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_312),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_268),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_130),
.B(n_268),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_193),
.Y(n_130)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_131),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_170),
.C(n_185),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_133),
.B(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_148),
.C(n_156),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_134),
.B(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_140),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g533 ( 
.A(n_135),
.B(n_262),
.C(n_349),
.Y(n_533)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_137),
.B(n_141),
.C(n_144),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_137),
.B(n_262),
.Y(n_346)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_139),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_143),
.Y(n_494)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_147),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_148),
.A2(n_149),
.B1(n_156),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_149),
.A2(n_375),
.B(n_378),
.Y(n_374)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_156),
.Y(n_406)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_162),
.C(n_166),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_158),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_157),
.A2(n_158),
.B1(n_166),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g347 ( 
.A(n_158),
.B(n_198),
.C(n_204),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_162),
.B(n_282),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_165),
.Y(n_247)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_166),
.Y(n_283)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_169),
.Y(n_365)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_169),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_170),
.A2(n_185),
.B1(n_186),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_170),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_180),
.C(n_182),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_171),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.C(n_176),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_172),
.A2(n_176),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_172),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_172),
.B(n_420),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_173),
.B(n_384),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_176),
.Y(n_386)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_178),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_308),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_182),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_192),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_188),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_188),
.B(n_362),
.C(n_368),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_188),
.A2(n_258),
.B1(n_368),
.B2(n_369),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_189),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_192),
.B(n_257),
.C(n_258),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_228),
.B1(n_266),
.B2(n_267),
.Y(n_193)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_194),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_209),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_195),
.B(n_210),
.C(n_216),
.Y(n_352)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_203),
.B1(n_204),
.B2(n_208),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_198),
.Y(n_208)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_202),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_203),
.A2(n_204),
.B1(n_215),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_211),
.C(n_215),
.Y(n_210)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_207),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_216),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_217),
.B(n_222),
.C(n_225),
.Y(n_329)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_255),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_229),
.B(n_256),
.C(n_259),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.C(n_248),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_230),
.B(n_233),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.C(n_244),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_234),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_239),
.A2(n_244),
.B1(n_245),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_244),
.B(n_394),
.C(n_396),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_244),
.A2(n_245),
.B1(n_394),
.B2(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_246),
.Y(n_423)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_251),
.C(n_254),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_260),
.B(n_265),
.C(n_351),
.Y(n_350)
);

XNOR2x1_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_262),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_266),
.B(n_354),
.C(n_355),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_274),
.C(n_277),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_270),
.A2(n_271),
.B1(n_274),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_274),
.Y(n_413)
);

XOR2x2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_278),
.B(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_305),
.C(n_309),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_279),
.B(n_408),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.C(n_294),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_281),
.B(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_284),
.B(n_294),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_291),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_285),
.B(n_291),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_290),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_299),
.C(n_300),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_295),
.A2(n_299),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_295),
.Y(n_390)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_299),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_299),
.B(n_464),
.C(n_466),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_299),
.A2(n_391),
.B1(n_466),
.B2(n_467),
.Y(n_477)
);

XOR2x1_ASAP7_75t_L g388 ( 
.A(n_300),
.B(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_306),
.B(n_309),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_312),
.A2(n_523),
.B(n_524),
.Y(n_522)
);

AND2x2_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_353),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_313),
.B(n_353),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_314),
.B(n_316),
.C(n_343),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_343),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_328),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_317),
.B(n_329),
.C(n_330),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_326),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_331),
.B(n_333),
.C(n_338),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_338),
.Y(n_332)
);

INVx8_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2x1_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_352),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_350),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_345),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.Y(n_345)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_346),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_347),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_350),
.B(n_556),
.C(n_557),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_352),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_518),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_409),
.C(n_414),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_401),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_359),
.B(n_401),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_387),
.C(n_399),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_360),
.B(n_516),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_373),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_374),
.C(n_383),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_362),
.B(n_508),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_366),
.Y(n_362)
);

XNOR2x1_ASAP7_75t_SL g453 ( 
.A(n_363),
.B(n_366),
.Y(n_453)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_363),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_363),
.A2(n_471),
.B1(n_472),
.B2(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_383),
.Y(n_373)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_385),
.B(n_421),
.C(n_424),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_387),
.B(n_399),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_392),
.C(n_397),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_388),
.B(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_393),
.B(n_398),
.Y(n_503)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

XOR2x2_ASAP7_75t_SL g447 ( 
.A(n_396),
.B(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_407),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_403),
.B(n_404),
.C(n_407),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_410),
.Y(n_520)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_411),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_415),
.A2(n_513),
.B(n_517),
.Y(n_414)
);

AOI21x1_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_499),
.B(n_512),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_458),
.B(n_498),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_444),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_418),
.B(n_444),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_428),
.C(n_435),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_419),
.B(n_461),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_424),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx6_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_428),
.A2(n_429),
.B1(n_435),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_434),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_430),
.B(n_434),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

AO22x1_ASAP7_75t_SL g435 ( 
.A1(n_436),
.A2(n_439),
.B1(n_442),
.B2(n_443),
.Y(n_435)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_436),
.Y(n_442)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_439),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_442),
.Y(n_451)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_440),
.Y(n_474)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_443),
.B(n_491),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_450),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_446),
.B(n_447),
.C(n_450),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

MAJx2_ASAP7_75t_L g510 ( 
.A(n_451),
.B(n_453),
.C(n_454),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_468),
.B(n_497),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_463),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_460),
.B(n_463),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_464),
.A2(n_465),
.B1(n_476),
.B2(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_469),
.A2(n_478),
.B(n_496),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_475),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_470),
.B(n_475),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_472),
.Y(n_470)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_472),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_479),
.A2(n_490),
.B(n_495),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_488),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_488),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_481),
.B(n_487),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_487),
.B(n_492),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_500),
.B(n_511),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_511),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_502),
.B1(n_504),
.B2(n_505),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_501),
.B(n_506),
.C(n_510),
.Y(n_514)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_507),
.B1(n_509),
.B2(n_510),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_514),
.B(n_515),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_520),
.C(n_521),
.Y(n_518)
);

NOR3xp33_ASAP7_75t_SL g525 ( 
.A(n_526),
.B(n_544),
.C(n_558),
.Y(n_525)
);

OAI21x1_ASAP7_75t_SL g563 ( 
.A1(n_526),
.A2(n_564),
.B(n_567),
.Y(n_563)
);

NOR2x1_ASAP7_75t_R g526 ( 
.A(n_527),
.B(n_542),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_527),
.B(n_542),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_534),
.C(n_539),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_528),
.B(n_547),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_531),
.C(n_533),
.Y(n_528)
);

INVxp33_ASAP7_75t_SL g529 ( 
.A(n_530),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_530),
.B(n_552),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_531),
.B(n_533),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_534),
.A2(n_539),
.B1(n_540),
.B2(n_548),
.Y(n_547)
);

INVxp33_ASAP7_75t_SL g548 ( 
.A(n_534),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_537),
.C(n_538),
.Y(n_534)
);

XNOR2x2_ASAP7_75t_L g553 ( 
.A(n_535),
.B(n_554),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_537),
.B(n_538),
.Y(n_554)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

AOI21x1_ASAP7_75t_L g564 ( 
.A1(n_545),
.A2(n_565),
.B(n_566),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_549),
.Y(n_545)
);

NOR2xp67_ASAP7_75t_SL g566 ( 
.A(n_546),
.B(n_549),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_550),
.B(n_553),
.C(n_555),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_550),
.A2(n_551),
.B1(n_553),
.B2(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_553),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_555),
.B(n_561),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_560),
.Y(n_558)
);

NOR2x1_ASAP7_75t_L g565 ( 
.A(n_559),
.B(n_560),
.Y(n_565)
);

NOR2xp67_ASAP7_75t_R g569 ( 
.A(n_570),
.B(n_578),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_570),
.B(n_578),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_571),
.B(n_572),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_573),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_575),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_580),
.Y(n_579)
);


endmodule