module fake_jpeg_4716_n_25 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_25);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_25;

wire n_21;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_24;
wire n_17;
wire n_15;

OR2x2_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_10),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_8),
.B(n_1),
.Y(n_15)
);

AO22x1_ASAP7_75t_SL g16 ( 
.A1(n_5),
.A2(n_2),
.B1(n_13),
.B2(n_6),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_11),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_3),
.B(n_7),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_0),
.A2(n_4),
.B(n_12),
.Y(n_19)
);

AO22x1_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_0),
.B1(n_4),
.B2(n_19),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_21),
.C(n_22),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_15),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_15),
.B1(n_18),
.B2(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_20),
.Y(n_25)
);


endmodule