module real_jpeg_20766_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_255;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_0),
.A2(n_69),
.B1(n_73),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_0),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_0),
.A2(n_56),
.B1(n_57),
.B2(n_109),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_109),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_109),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_2),
.A2(n_69),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_2),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_2),
.A2(n_56),
.B1(n_57),
.B2(n_74),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_74),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_74),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_3),
.A2(n_36),
.B1(n_69),
.B2(n_73),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_3),
.A2(n_36),
.B1(n_56),
.B2(n_57),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_3),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_4),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_4),
.B(n_71),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_4),
.A2(n_14),
.B(n_29),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_124),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_4),
.A2(n_82),
.B1(n_101),
.B2(n_197),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_4),
.B(n_170),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_4),
.B(n_56),
.Y(n_221)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_4),
.A2(n_56),
.B(n_221),
.Y(n_225)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_6),
.A2(n_69),
.B1(n_73),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_6),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_135),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_135),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_135),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_28),
.Y(n_31)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_7),
.Y(n_101)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_9),
.A2(n_30),
.B1(n_56),
.B2(n_57),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_9),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_11),
.A2(n_47),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_47),
.Y(n_126)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_13),
.A2(n_56),
.B1(n_57),
.B2(n_68),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_14),
.A2(n_39),
.B(n_43),
.C(n_44),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_39),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_15),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_138),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_19),
.B(n_111),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_89),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_78),
.B2(n_79),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_24),
.B(n_37),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_32),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_25),
.A2(n_101),
.B(n_126),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_27),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_28),
.B(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_31),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_31),
.A2(n_35),
.B(n_100),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_32),
.A2(n_82),
.B(n_184),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_34),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_34),
.A2(n_82),
.B1(n_181),
.B2(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_35),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_38),
.A2(n_48),
.B(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_38),
.A2(n_85),
.B(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_38),
.A2(n_44),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_38),
.A2(n_44),
.B1(n_192),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_38),
.A2(n_44),
.B1(n_212),
.B2(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_38),
.A2(n_228),
.B(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_40),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

AOI32xp33_ASAP7_75t_L g220 ( 
.A1(n_39),
.A2(n_54),
.A3(n_57),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_40),
.A2(n_45),
.B(n_124),
.C(n_188),
.Y(n_187)
);

NAND2xp33_ASAP7_75t_SL g222 ( 
.A(n_40),
.B(n_53),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_44),
.A2(n_46),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_44),
.B(n_124),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_64),
.B1(n_65),
.B2(n_77),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_55),
.B(n_58),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_53),
.B(n_56),
.C(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_63),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_52),
.B(n_104),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_52),
.A2(n_60),
.B1(n_129),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_52),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_52),
.A2(n_60),
.B1(n_169),
.B2(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_56),
.Y(n_61)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_68),
.Y(n_122)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_57),
.A2(n_70),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_59),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_59),
.A2(n_128),
.B(n_130),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_59),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_72),
.B(n_75),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_72),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_66),
.A2(n_108),
.B1(n_110),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_67),
.A2(n_71),
.B1(n_123),
.B2(n_134),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.C(n_71),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_69),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g123 ( 
.A(n_69),
.B(n_124),
.CON(n_123),
.SN(n_123)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_71),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_84),
.B2(n_88),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_82),
.A2(n_98),
.B1(n_101),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_87),
.B(n_148),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_102),
.C(n_106),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_91),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_101),
.B(n_124),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_106),
.B1(n_107),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_118),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_112),
.A2(n_116),
.B1(n_117),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_112),
.Y(n_257)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_118),
.A2(n_119),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_127),
.C(n_131),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_125),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_131),
.B1(n_132),
.B2(n_155),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_127),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_172),
.B(n_252),
.C(n_258),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_157),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_140),
.B(n_157),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_153),
.B2(n_156),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_143),
.B(n_144),
.C(n_156),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.C(n_152),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_151),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_152),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_158),
.B(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_167),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_166),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_167),
.B(n_238),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_251),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_246),
.B(n_250),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_233),
.B(n_245),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_215),
.B(n_232),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_204),
.B(n_214),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_193),
.B(n_203),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_185),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_185),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_187),
.B(n_189),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_198),
.B(n_202),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_196),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_205),
.B(n_206),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_213),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_217),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_223),
.B1(n_230),
.B2(n_231),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_218),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_223),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_226),
.B1(n_227),
.B2(n_229),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_224),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_229),
.C(n_230),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_234),
.B(n_235),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_240),
.B2(n_241),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_242),
.C(n_244),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_247),
.B(n_248),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_254),
.Y(n_258)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);


endmodule