module fake_jpeg_22033_n_150 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_150);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_0),
.CON(n_37),
.SN(n_37)
);

NOR3xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_17),
.C(n_16),
.Y(n_61)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_42),
.B1(n_18),
.B2(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_40),
.A2(n_32),
.B1(n_15),
.B2(n_19),
.Y(n_70)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_44),
.Y(n_52)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_23),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_24),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_55),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_29),
.B1(n_18),
.B2(n_30),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_32),
.B1(n_21),
.B2(n_5),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_59),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

CKINVDCx6p67_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_25),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_42),
.B1(n_37),
.B2(n_31),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_66),
.B1(n_70),
.B2(n_6),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_31),
.B1(n_30),
.B2(n_15),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_17),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_73),
.B(n_84),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_2),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_87),
.C(n_94),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_57),
.B1(n_62),
.B2(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_3),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_13),
.B(n_7),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_69),
.B(n_10),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_6),
.C(n_7),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_91),
.Y(n_105)
);

CKINVDCx12_ASAP7_75t_R g90 ( 
.A(n_48),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_9),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_9),
.C(n_10),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_65),
.B(n_58),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_100),
.B(n_111),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_73),
.B(n_92),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_87),
.B1(n_76),
.B2(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_51),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_108),
.Y(n_118)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_53),
.A3(n_51),
.B1(n_68),
.B2(n_56),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_77),
.Y(n_109)
);

OR2x2_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_79),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_80),
.C(n_83),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_115),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_110),
.C(n_95),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_75),
.B1(n_74),
.B2(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NOR4xp25_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_74),
.C(n_78),
.D(n_93),
.Y(n_121)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_99),
.CI(n_101),
.CON(n_130),
.SN(n_130)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_104),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_108),
.B1(n_103),
.B2(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_133),
.B(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_118),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_78),
.B(n_97),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_118),
.B1(n_116),
.B2(n_115),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_132),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_133),
.A2(n_114),
.B(n_112),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_138),
.B(n_127),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_139),
.B(n_141),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_143),
.B(n_145),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_135),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_144),
.A3(n_120),
.B1(n_117),
.B2(n_85),
.C1(n_78),
.C2(n_106),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_78),
.C(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_149),
.Y(n_150)
);


endmodule