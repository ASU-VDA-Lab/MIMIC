module fake_netlist_1_5124_n_520 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_520);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_520;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_45), .Y(n_76) );
INVxp67_ASAP7_75t_SL g77 ( .A(n_19), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_1), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_69), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_16), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_72), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_35), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_28), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_26), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_16), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_70), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_40), .Y(n_87) );
OR2x2_ASAP7_75t_L g88 ( .A(n_3), .B(n_56), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_9), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_4), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_14), .Y(n_91) );
INVx3_ASAP7_75t_L g92 ( .A(n_38), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_64), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_74), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_4), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_52), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_31), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_55), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_73), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_20), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_71), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_43), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_8), .Y(n_103) );
NOR2xp67_ASAP7_75t_L g104 ( .A(n_12), .B(n_33), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_17), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_8), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_54), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_11), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_39), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_41), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_92), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_92), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_76), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_85), .B(n_0), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_92), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_97), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_85), .B(n_0), .Y(n_117) );
INVxp67_ASAP7_75t_L g118 ( .A(n_89), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_76), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_81), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_81), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_89), .B(n_1), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_96), .B(n_2), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_97), .Y(n_124) );
INVx5_ASAP7_75t_L g125 ( .A(n_101), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_83), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_98), .B(n_2), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
BUFx12f_ASAP7_75t_L g130 ( .A(n_93), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_101), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_110), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_84), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_122), .B(n_90), .Y(n_134) );
AND2x6_ASAP7_75t_L g135 ( .A(n_122), .B(n_86), .Y(n_135) );
INVxp67_ASAP7_75t_SL g136 ( .A(n_118), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_111), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_130), .Y(n_138) );
INVx4_ASAP7_75t_L g139 ( .A(n_125), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_118), .B(n_102), .Y(n_140) );
OR2x2_ASAP7_75t_L g141 ( .A(n_113), .B(n_80), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_130), .B(n_82), .Y(n_142) );
INVx6_ASAP7_75t_L g143 ( .A(n_111), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_122), .B(n_113), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_130), .B(n_100), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_119), .B(n_93), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_111), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_111), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_119), .B(n_109), .Y(n_150) );
INVx1_ASAP7_75t_SL g151 ( .A(n_122), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_111), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_111), .Y(n_153) );
NOR2x1p5_ASAP7_75t_L g154 ( .A(n_114), .B(n_80), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_120), .B(n_90), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_112), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_122), .B(n_103), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_120), .B(n_109), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_137), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_140), .B(n_121), .Y(n_160) );
OR2x6_ASAP7_75t_L g161 ( .A(n_144), .B(n_114), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_156), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_156), .Y(n_163) );
INVx2_ASAP7_75t_SL g164 ( .A(n_144), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_147), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_135), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_147), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_136), .B(n_121), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_134), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_135), .Y(n_174) );
INVx5_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_138), .Y(n_176) );
NAND3xp33_ASAP7_75t_L g177 ( .A(n_134), .B(n_133), .C(n_128), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_157), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_142), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_141), .B(n_128), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_157), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_141), .B(n_129), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_157), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_158), .B(n_129), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_135), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_145), .B(n_133), .Y(n_187) );
OR2x6_ASAP7_75t_L g188 ( .A(n_157), .B(n_117), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_135), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_155), .B(n_132), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_188), .A2(n_135), .B1(n_154), .B2(n_151), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_180), .B(n_146), .Y(n_193) );
INVx5_ASAP7_75t_L g194 ( .A(n_174), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_181), .B(n_135), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_SL g196 ( .A1(n_185), .A2(n_149), .B(n_148), .C(n_153), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_188), .A2(n_135), .B1(n_155), .B2(n_154), .Y(n_197) );
BUFx2_ASAP7_75t_SL g198 ( .A(n_174), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_160), .A2(n_126), .B(n_132), .C(n_123), .Y(n_199) );
INVx1_ASAP7_75t_SL g200 ( .A(n_161), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_162), .Y(n_201) );
NAND2x1p5_ASAP7_75t_L g202 ( .A(n_174), .B(n_126), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_163), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_163), .Y(n_204) );
INVx1_ASAP7_75t_SL g205 ( .A(n_161), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_183), .B(n_150), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_183), .B(n_78), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_189), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_174), .B(n_126), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_188), .B(n_126), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_177), .A2(n_153), .B(n_152), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_188), .B(n_132), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_188), .B(n_132), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_186), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_186), .Y(n_215) );
INVx4_ASAP7_75t_L g216 ( .A(n_189), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_189), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_186), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_161), .B(n_117), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_169), .Y(n_220) );
INVx2_ASAP7_75t_SL g221 ( .A(n_167), .Y(n_221) );
BUFx2_ASAP7_75t_SL g222 ( .A(n_167), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_191), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_207), .A2(n_161), .B1(n_164), .B2(n_173), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_191), .B(n_187), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_191), .Y(n_226) );
BUFx2_ASAP7_75t_L g227 ( .A(n_202), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_204), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_200), .A2(n_161), .B1(n_164), .B2(n_184), .Y(n_229) );
BUFx4f_ASAP7_75t_SL g230 ( .A(n_216), .Y(n_230) );
OAI211xp5_ASAP7_75t_L g231 ( .A1(n_197), .A2(n_127), .B(n_190), .C(n_171), .Y(n_231) );
OAI21x1_ASAP7_75t_L g232 ( .A1(n_211), .A2(n_148), .B(n_149), .Y(n_232) );
INVx8_ASAP7_75t_L g233 ( .A(n_194), .Y(n_233) );
INVx1_ASAP7_75t_SL g234 ( .A(n_200), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_194), .Y(n_235) );
NAND2xp33_ASAP7_75t_L g236 ( .A(n_194), .B(n_186), .Y(n_236) );
AO31x2_ASAP7_75t_L g237 ( .A1(n_199), .A2(n_124), .A3(n_116), .B(n_115), .Y(n_237) );
OAI222xp33_ASAP7_75t_L g238 ( .A1(n_205), .A2(n_88), .B1(n_108), .B2(n_103), .C1(n_176), .C2(n_94), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_204), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_204), .B(n_169), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_219), .A2(n_177), .B1(n_184), .B2(n_179), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_201), .Y(n_242) );
OAI22xp33_ASAP7_75t_L g243 ( .A1(n_219), .A2(n_79), .B1(n_99), .B2(n_108), .Y(n_243) );
OAI222xp33_ASAP7_75t_L g244 ( .A1(n_205), .A2(n_88), .B1(n_77), .B2(n_95), .C1(n_91), .C2(n_105), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_201), .B(n_182), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_193), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_203), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_202), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_243), .A2(n_197), .B1(n_213), .B2(n_212), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_228), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_225), .A2(n_195), .B1(n_203), .B2(n_192), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_243), .A2(n_212), .B1(n_213), .B2(n_195), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_228), .Y(n_253) );
NAND2xp33_ASAP7_75t_SL g254 ( .A(n_248), .B(n_212), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_224), .A2(n_213), .B1(n_206), .B2(n_209), .Y(n_255) );
AOI221xp5_ASAP7_75t_L g256 ( .A1(n_238), .A2(n_206), .B1(n_220), .B2(n_210), .C(n_173), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_248), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_246), .A2(n_209), .B1(n_220), .B2(n_210), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_223), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_223), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_227), .B(n_194), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_223), .B(n_209), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_225), .A2(n_168), .B1(n_222), .B2(n_209), .Y(n_263) );
AOI222xp33_ASAP7_75t_L g264 ( .A1(n_238), .A2(n_106), .B1(n_168), .B2(n_182), .C1(n_172), .C2(n_179), .Y(n_264) );
OAI211xp5_ASAP7_75t_SL g265 ( .A1(n_231), .A2(n_107), .B(n_87), .C(n_86), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_242), .A2(n_172), .B1(n_221), .B2(n_222), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_226), .B(n_202), .Y(n_267) );
AOI221xp5_ASAP7_75t_L g268 ( .A1(n_244), .A2(n_196), .B1(n_116), .B2(n_124), .C(n_115), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_242), .A2(n_221), .B1(n_198), .B2(n_216), .Y(n_269) );
NOR3xp33_ASAP7_75t_SL g270 ( .A(n_256), .B(n_244), .C(n_231), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_261), .B(n_226), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_264), .A2(n_247), .B1(n_245), .B2(n_241), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_254), .A2(n_241), .B1(n_229), .B2(n_227), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_252), .A2(n_247), .B1(n_245), .B2(n_230), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_250), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_249), .B(n_245), .Y(n_276) );
OAI211xp5_ASAP7_75t_L g277 ( .A1(n_258), .A2(n_104), .B(n_124), .C(n_116), .Y(n_277) );
OAI21xp33_ASAP7_75t_L g278 ( .A1(n_265), .A2(n_87), .B(n_110), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_263), .A2(n_239), .B1(n_226), .B2(n_240), .Y(n_279) );
OAI31xp33_ASAP7_75t_L g280 ( .A1(n_251), .A2(n_202), .A3(n_234), .B(n_240), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_259), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_250), .B(n_239), .Y(n_282) );
OAI221xp5_ASAP7_75t_L g283 ( .A1(n_255), .A2(n_234), .B1(n_239), .B2(n_112), .C(n_115), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_259), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_263), .A2(n_230), .B1(n_233), .B2(n_221), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_253), .Y(n_286) );
OAI22xp33_ASAP7_75t_L g287 ( .A1(n_257), .A2(n_233), .B1(n_235), .B2(n_194), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_261), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_253), .B(n_237), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_262), .B(n_216), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_281), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_272), .A2(n_270), .B1(n_274), .B2(n_273), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_281), .B(n_260), .Y(n_293) );
AOI33xp33_ASAP7_75t_L g294 ( .A1(n_272), .A2(n_112), .A3(n_268), .B1(n_262), .B2(n_266), .B3(n_260), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_284), .B(n_267), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_284), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_282), .B(n_267), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_282), .B(n_237), .Y(n_298) );
NAND4xp25_ASAP7_75t_SL g299 ( .A(n_285), .B(n_269), .C(n_261), .D(n_6), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_276), .A2(n_233), .B1(n_235), .B2(n_236), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_288), .B(n_3), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_289), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_288), .B(n_237), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_275), .B(n_237), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_286), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_271), .B(n_237), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_288), .B(n_237), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_271), .Y(n_308) );
AOI33xp33_ASAP7_75t_L g309 ( .A1(n_287), .A2(n_152), .A3(n_6), .B1(n_7), .B2(n_9), .B3(n_10), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_271), .B(n_237), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_280), .Y(n_311) );
INVx5_ASAP7_75t_L g312 ( .A(n_279), .Y(n_312) );
AND2x4_ASAP7_75t_SL g313 ( .A(n_290), .B(n_216), .Y(n_313) );
INVxp67_ASAP7_75t_L g314 ( .A(n_290), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_283), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_277), .Y(n_316) );
OAI22xp33_ASAP7_75t_L g317 ( .A1(n_278), .A2(n_233), .B1(n_235), .B2(n_194), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_275), .B(n_232), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_281), .B(n_5), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_281), .B(n_5), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_302), .B(n_131), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_302), .B(n_306), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_291), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_303), .B(n_131), .Y(n_324) );
OAI22xp33_ASAP7_75t_L g325 ( .A1(n_292), .A2(n_233), .B1(n_194), .B2(n_217), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_296), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_296), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_302), .B(n_131), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_291), .B(n_131), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_306), .B(n_131), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_299), .A2(n_233), .B1(n_198), .B2(n_232), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_311), .B(n_131), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_297), .B(n_7), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_301), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_297), .B(n_10), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_295), .B(n_11), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_298), .B(n_131), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_305), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_298), .B(n_232), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_295), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_319), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_299), .A2(n_218), .B1(n_215), .B2(n_214), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_303), .B(n_12), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_292), .A2(n_218), .B1(n_215), .B2(n_214), .Y(n_344) );
NOR3xp33_ASAP7_75t_L g345 ( .A(n_309), .B(n_218), .C(n_215), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_305), .B(n_13), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_303), .B(n_57), .Y(n_347) );
NAND3xp33_ASAP7_75t_SL g348 ( .A(n_294), .B(n_13), .C(n_14), .Y(n_348) );
NAND2x1p5_ASAP7_75t_L g349 ( .A(n_319), .B(n_217), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_303), .B(n_15), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_314), .B(n_15), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_293), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_296), .B(n_59), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_314), .B(n_17), .Y(n_354) );
NOR3xp33_ASAP7_75t_SL g355 ( .A(n_316), .B(n_18), .C(n_19), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_310), .B(n_18), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_293), .Y(n_357) );
NAND3xp33_ASAP7_75t_SL g358 ( .A(n_315), .B(n_211), .C(n_22), .Y(n_358) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_317), .A2(n_217), .B(n_208), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_293), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_293), .B(n_21), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_310), .B(n_125), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_307), .B(n_125), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_338), .Y(n_365) );
OAI31xp33_ASAP7_75t_L g366 ( .A1(n_325), .A2(n_311), .A3(n_316), .B(n_313), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_322), .B(n_307), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_326), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_340), .B(n_304), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_322), .B(n_312), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_339), .B(n_312), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_334), .B(n_308), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_339), .B(n_312), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_330), .B(n_312), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_330), .B(n_312), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_357), .B(n_312), .Y(n_376) );
NOR3xp33_ASAP7_75t_L g377 ( .A(n_348), .B(n_315), .C(n_311), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_357), .B(n_312), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_356), .B(n_304), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_356), .B(n_320), .Y(n_380) );
XNOR2xp5_ASAP7_75t_L g381 ( .A(n_343), .B(n_313), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_323), .B(n_318), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_362), .B(n_311), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_327), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_337), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_344), .A2(n_308), .B1(n_318), .B2(n_313), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_341), .B(n_300), .Y(n_387) );
INVx1_ASAP7_75t_SL g388 ( .A(n_336), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_337), .Y(n_389) );
OAI21xp33_ASAP7_75t_L g390 ( .A1(n_355), .A2(n_178), .B(n_159), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_321), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_343), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_352), .B(n_23), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_321), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_360), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_328), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_324), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_329), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_324), .B(n_24), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_329), .B(n_25), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_324), .B(n_27), .Y(n_401) );
OAI31xp33_ASAP7_75t_L g402 ( .A1(n_350), .A2(n_218), .A3(n_215), .B(n_214), .Y(n_402) );
AOI322xp5_ASAP7_75t_L g403 ( .A1(n_350), .A2(n_125), .A3(n_214), .B1(n_32), .B2(n_34), .C1(n_36), .C2(n_37), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_333), .B(n_29), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_328), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_335), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_363), .B(n_364), .Y(n_407) );
NAND4xp25_ASAP7_75t_L g408 ( .A(n_354), .B(n_351), .C(n_346), .D(n_358), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_364), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_353), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_353), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_353), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_347), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_367), .B(n_347), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_408), .B(n_332), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_365), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_365), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_395), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_367), .B(n_397), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_395), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_377), .A2(n_347), .B1(n_332), .B2(n_345), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_388), .A2(n_363), .B1(n_361), .B2(n_349), .C(n_331), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_382), .Y(n_423) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_404), .B(n_342), .C(n_359), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_383), .B(n_349), .Y(n_425) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_399), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_382), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_385), .B(n_389), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_385), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_409), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_409), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_397), .B(n_30), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_407), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_407), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_392), .B(n_42), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_384), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_381), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_369), .B(n_44), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_384), .Y(n_439) );
OAI221xp5_ASAP7_75t_L g440 ( .A1(n_366), .A2(n_125), .B1(n_143), .B2(n_208), .C(n_217), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_379), .B(n_46), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_398), .B(n_47), .Y(n_442) );
XOR2x2_ASAP7_75t_L g443 ( .A(n_381), .B(n_48), .Y(n_443) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_372), .B(n_125), .C(n_208), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_398), .B(n_49), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_370), .B(n_50), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_396), .B(n_405), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_396), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_405), .B(n_51), .Y(n_449) );
AOI32xp33_ASAP7_75t_L g450 ( .A1(n_413), .A2(n_53), .A3(n_58), .B1(n_60), .B2(n_61), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_391), .B(n_62), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_386), .B(n_125), .Y(n_452) );
OAI21xp5_ASAP7_75t_SL g453 ( .A1(n_402), .A2(n_217), .B(n_208), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_368), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_380), .B(n_406), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_413), .B(n_217), .Y(n_456) );
XNOR2xp5_ASAP7_75t_L g457 ( .A(n_387), .B(n_63), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_391), .B(n_65), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_370), .B(n_66), .Y(n_459) );
XOR2xp5_ASAP7_75t_L g460 ( .A(n_371), .B(n_67), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_393), .A2(n_178), .B(n_165), .C(n_170), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_393), .B(n_208), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_394), .B(n_68), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_394), .Y(n_464) );
OAI221xp5_ASAP7_75t_L g465 ( .A1(n_403), .A2(n_143), .B1(n_170), .B2(n_165), .C(n_159), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_376), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_399), .B(n_159), .Y(n_467) );
AOI322xp5_ASAP7_75t_L g468 ( .A1(n_373), .A2(n_75), .A3(n_165), .B1(n_166), .B2(n_170), .C1(n_175), .C2(n_139), .Y(n_468) );
NAND4xp75_ASAP7_75t_L g469 ( .A(n_401), .B(n_166), .C(n_175), .D(n_139), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_410), .Y(n_470) );
OAI21xp33_ASAP7_75t_SL g471 ( .A1(n_373), .A2(n_166), .B(n_175), .Y(n_471) );
OAI21xp5_ASAP7_75t_SL g472 ( .A1(n_401), .A2(n_175), .B(n_374), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_410), .B(n_175), .Y(n_473) );
OAI21xp33_ASAP7_75t_L g474 ( .A1(n_374), .A2(n_175), .B(n_375), .Y(n_474) );
OAI21xp33_ASAP7_75t_L g475 ( .A1(n_375), .A2(n_376), .B(n_378), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_SL g476 ( .A1(n_411), .A2(n_412), .B(n_378), .C(n_400), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_411), .B(n_412), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_400), .B(n_390), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_365), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_367), .B(n_371), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_423), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_437), .A2(n_472), .B1(n_421), .B2(n_460), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_415), .B(n_421), .C(n_422), .Y(n_483) );
NAND3xp33_ASAP7_75t_SL g484 ( .A(n_450), .B(n_453), .C(n_422), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_480), .B(n_419), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_415), .A2(n_452), .B1(n_427), .B2(n_475), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_455), .B(n_428), .Y(n_487) );
OAI21xp33_ASAP7_75t_SL g488 ( .A1(n_480), .A2(n_462), .B(n_452), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_433), .B(n_434), .Y(n_489) );
AOI221xp5_ASAP7_75t_SL g490 ( .A1(n_440), .A2(n_474), .B1(n_414), .B2(n_466), .C(n_447), .Y(n_490) );
INVx2_ASAP7_75t_SL g491 ( .A(n_426), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_426), .A2(n_478), .B1(n_440), .B2(n_466), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_431), .A2(n_430), .B1(n_477), .B2(n_429), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_448), .B(n_457), .Y(n_494) );
OAI21xp33_ASAP7_75t_SL g495 ( .A1(n_462), .A2(n_432), .B(n_467), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_471), .A2(n_443), .B(n_467), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_476), .A2(n_461), .B(n_456), .Y(n_497) );
AOI221xp5_ASAP7_75t_L g498 ( .A1(n_483), .A2(n_476), .B1(n_470), .B2(n_418), .C(n_420), .Y(n_498) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_484), .B(n_469), .Y(n_499) );
OAI21xp33_ASAP7_75t_L g500 ( .A1(n_488), .A2(n_425), .B(n_477), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_481), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_493), .Y(n_502) );
AOI211xp5_ASAP7_75t_L g503 ( .A1(n_482), .A2(n_424), .B(n_426), .C(n_465), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_490), .A2(n_424), .B1(n_426), .B2(n_417), .Y(n_504) );
AOI211xp5_ASAP7_75t_L g505 ( .A1(n_495), .A2(n_446), .B(n_459), .C(n_444), .Y(n_505) );
XNOR2xp5_ASAP7_75t_L g506 ( .A(n_486), .B(n_464), .Y(n_506) );
NOR4xp75_ASAP7_75t_L g507 ( .A(n_500), .B(n_496), .C(n_492), .D(n_491), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g508 ( .A(n_499), .B(n_497), .C(n_494), .D(n_468), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_503), .A2(n_489), .B1(n_487), .B2(n_485), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_504), .A2(n_502), .B1(n_505), .B2(n_506), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_501), .B(n_489), .Y(n_511) );
OAI221xp5_ASAP7_75t_L g512 ( .A1(n_508), .A2(n_498), .B1(n_441), .B2(n_438), .C(n_442), .Y(n_512) );
AND4x1_ASAP7_75t_L g513 ( .A(n_510), .B(n_435), .C(n_445), .D(n_449), .Y(n_513) );
OAI221xp5_ASAP7_75t_L g514 ( .A1(n_509), .A2(n_416), .B1(n_479), .B2(n_439), .C(n_436), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_513), .Y(n_515) );
XNOR2xp5_ASAP7_75t_L g516 ( .A(n_512), .B(n_507), .Y(n_516) );
OAI22xp33_ASAP7_75t_SL g517 ( .A1(n_516), .A2(n_514), .B1(n_511), .B2(n_451), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_517), .B(n_515), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_518), .A2(n_463), .B(n_458), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_519), .A2(n_473), .B(n_454), .Y(n_520) );
endmodule