module fake_aes_395_n_27 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_27);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
BUFx2_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
AOI22xp5_ASAP7_75t_L g15 ( .A1(n_11), .A2(n_0), .B1(n_5), .B2(n_6), .Y(n_15) );
AOI21x1_ASAP7_75t_L g16 ( .A1(n_12), .A2(n_8), .B(n_0), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_2), .B(n_1), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_10), .Y(n_18) );
OR2x6_ASAP7_75t_L g19 ( .A(n_1), .B(n_4), .Y(n_19) );
AOI21xp5_ASAP7_75t_L g20 ( .A1(n_14), .A2(n_3), .B(n_9), .Y(n_20) );
A2O1A1Ixp33_ASAP7_75t_L g21 ( .A1(n_18), .A2(n_2), .B(n_13), .C(n_15), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_21), .B(n_19), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_20), .Y(n_23) );
INVx2_ASAP7_75t_SL g24 ( .A(n_23), .Y(n_24) );
NAND2x1p5_ASAP7_75t_L g25 ( .A(n_24), .B(n_17), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_25), .B(n_24), .Y(n_26) );
OAI21xp5_ASAP7_75t_SL g27 ( .A1(n_26), .A2(n_16), .B(n_19), .Y(n_27) );
endmodule