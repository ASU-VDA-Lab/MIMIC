module real_aes_10588_n_360 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_1966, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_360);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_1966;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_360;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_1929;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_501;
wire n_488;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1940;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1914;
wire n_724;
wire n_1648;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_1638;
wire n_1072;
wire n_495;
wire n_370;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_367;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1855;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_1226;
wire n_1617;
wire n_525;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1691;
wire n_640;
wire n_1931;
wire n_1176;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1584;
wire n_1277;
wire n_1049;
wire n_1950;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_1025;
wire n_532;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_729;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g1903 ( .A1(n_0), .A2(n_174), .B1(n_1400), .B2(n_1904), .C(n_1905), .Y(n_1903) );
AOI221xp5_ASAP7_75t_L g1935 ( .A1(n_0), .A2(n_359), .B1(n_608), .B2(n_1165), .C(n_1936), .Y(n_1935) );
INVxp67_ASAP7_75t_SL g1208 ( .A(n_1), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_1), .A2(n_347), .B1(n_784), .B2(n_1235), .Y(n_1234) );
OA22x2_ASAP7_75t_L g727 ( .A1(n_2), .A2(n_728), .B1(n_802), .B2(n_803), .Y(n_727) );
INVxp67_ASAP7_75t_SL g803 ( .A(n_2), .Y(n_803) );
INVx1_ASAP7_75t_L g1474 ( .A(n_3), .Y(n_1474) );
INVx1_ASAP7_75t_L g1714 ( .A(n_4), .Y(n_1714) );
INVx1_ASAP7_75t_L g1573 ( .A(n_5), .Y(n_1573) );
INVxp33_ASAP7_75t_L g1228 ( .A(n_6), .Y(n_1228) );
AOI21xp33_ASAP7_75t_L g1244 ( .A1(n_6), .A2(n_600), .B(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g994 ( .A(n_7), .Y(n_994) );
AOI221xp5_ASAP7_75t_SL g1016 ( .A1(n_7), .A2(n_135), .B1(n_610), .B2(n_770), .C(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g1216 ( .A(n_8), .Y(n_1216) );
INVx1_ASAP7_75t_L g987 ( .A(n_9), .Y(n_987) );
AOI221xp5_ASAP7_75t_L g1025 ( .A1(n_9), .A2(n_239), .B1(n_766), .B2(n_1026), .C(n_1027), .Y(n_1025) );
AOI22xp33_ASAP7_75t_SL g936 ( .A1(n_10), .A2(n_160), .B1(n_937), .B2(n_939), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_10), .A2(n_57), .B1(n_588), .B2(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g1278 ( .A(n_11), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_12), .A2(n_298), .B1(n_1114), .B2(n_1115), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_12), .A2(n_332), .B1(n_784), .B2(n_889), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1330 ( .A1(n_13), .A2(n_65), .B1(n_667), .B2(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g1354 ( .A(n_13), .Y(n_1354) );
XNOR2x2_ASAP7_75t_L g929 ( .A(n_14), .B(n_930), .Y(n_929) );
AO221x2_ASAP7_75t_L g1712 ( .A1(n_14), .A2(n_272), .B1(n_1669), .B2(n_1691), .C(n_1713), .Y(n_1712) );
INVxp33_ASAP7_75t_L g1226 ( .A(n_15), .Y(n_1226) );
NAND2xp33_ASAP7_75t_SL g1242 ( .A(n_15), .B(n_1243), .Y(n_1242) );
AOI22xp33_ASAP7_75t_SL g941 ( .A1(n_16), .A2(n_57), .B1(n_716), .B2(n_942), .Y(n_941) );
AOI21xp33_ASAP7_75t_L g965 ( .A1(n_16), .A2(n_465), .B(n_698), .Y(n_965) );
CKINVDCx16_ASAP7_75t_R g1723 ( .A(n_17), .Y(n_1723) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_18), .A2(n_249), .B1(n_731), .B2(n_732), .Y(n_730) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_18), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g673 ( .A(n_19), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g1268 ( .A1(n_20), .A2(n_299), .B1(n_883), .B2(n_1262), .Y(n_1268) );
INVxp67_ASAP7_75t_SL g1303 ( .A(n_20), .Y(n_1303) );
INVxp33_ASAP7_75t_L g1482 ( .A(n_21), .Y(n_1482) );
AOI221xp5_ASAP7_75t_L g1528 ( .A1(n_21), .A2(n_77), .B1(n_1067), .B2(n_1529), .C(n_1530), .Y(n_1528) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_22), .A2(n_69), .B1(n_585), .B2(n_587), .C(n_590), .Y(n_584) );
INVx1_ASAP7_75t_L g641 ( .A(n_22), .Y(n_641) );
INVx1_ASAP7_75t_L g956 ( .A(n_23), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_23), .A2(n_309), .B1(n_588), .B2(n_698), .Y(n_967) );
OAI221xp5_ASAP7_75t_L g1221 ( .A1(n_24), .A2(n_326), .B1(n_738), .B2(n_989), .C(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1246 ( .A(n_24), .Y(n_1246) );
AOI221xp5_ASAP7_75t_L g1310 ( .A1(n_25), .A2(n_355), .B1(n_469), .B2(n_1311), .C(n_1313), .Y(n_1310) );
INVx1_ASAP7_75t_L g1342 ( .A(n_25), .Y(n_1342) );
OAI22xp5_ASAP7_75t_L g1378 ( .A1(n_26), .A2(n_349), .B1(n_427), .B2(n_1074), .Y(n_1378) );
INVxp67_ASAP7_75t_SL g1418 ( .A(n_26), .Y(n_1418) );
INVx1_ASAP7_75t_L g1613 ( .A(n_27), .Y(n_1613) );
AOI22xp33_ASAP7_75t_L g1641 ( .A1(n_27), .A2(n_56), .B1(n_1642), .B2(n_1643), .Y(n_1641) );
INVx1_ASAP7_75t_L g1141 ( .A(n_28), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_29), .A2(n_168), .B1(n_1115), .B2(n_1120), .Y(n_1119) );
INVxp67_ASAP7_75t_L g1133 ( .A(n_29), .Y(n_1133) );
INVxp33_ASAP7_75t_L g1603 ( .A(n_30), .Y(n_1603) );
AOI22xp33_ASAP7_75t_L g1633 ( .A1(n_30), .A2(n_81), .B1(n_588), .B2(n_898), .Y(n_1633) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_31), .A2(n_346), .B1(n_1240), .B2(n_1504), .Y(n_1503) );
INVxp67_ASAP7_75t_SL g1541 ( .A(n_31), .Y(n_1541) );
OAI211xp5_ASAP7_75t_SL g1259 ( .A1(n_32), .A2(n_482), .B(n_1260), .C(n_1271), .Y(n_1259) );
AOI221xp5_ASAP7_75t_L g1298 ( .A1(n_32), .A2(n_200), .B1(n_942), .B2(n_1299), .C(n_1301), .Y(n_1298) );
INVx1_ASAP7_75t_L g617 ( .A(n_33), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g988 ( .A1(n_34), .A2(n_314), .B1(n_737), .B2(n_738), .C(n_989), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_34), .A2(n_314), .B1(n_776), .B2(n_777), .Y(n_1024) );
INVx1_ASAP7_75t_L g366 ( .A(n_35), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_36), .A2(n_317), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
AOI221xp5_ASAP7_75t_L g1086 ( .A1(n_36), .A2(n_155), .B1(n_465), .B2(n_688), .C(n_1087), .Y(n_1086) );
OAI221xp5_ASAP7_75t_L g1609 ( .A1(n_37), .A2(n_206), .B1(n_520), .B2(n_531), .C(n_737), .Y(n_1609) );
OAI33xp33_ASAP7_75t_L g1636 ( .A1(n_37), .A2(n_206), .A3(n_473), .B1(n_677), .B2(n_778), .B3(n_1966), .Y(n_1636) );
OAI221xp5_ASAP7_75t_L g736 ( .A1(n_38), .A2(n_70), .B1(n_520), .B2(n_737), .C(n_738), .Y(n_736) );
OAI222xp33_ASAP7_75t_L g775 ( .A1(n_38), .A2(n_70), .B1(n_236), .B2(n_616), .C1(n_776), .C2(n_777), .Y(n_775) );
INVx1_ASAP7_75t_L g1219 ( .A(n_39), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g1566 ( .A1(n_40), .A2(n_64), .B1(n_427), .B2(n_1567), .Y(n_1566) );
OAI221xp5_ASAP7_75t_L g1586 ( .A1(n_40), .A2(n_64), .B1(n_738), .B2(n_989), .C(n_1222), .Y(n_1586) );
AOI21xp33_ASAP7_75t_L g687 ( .A1(n_41), .A2(n_688), .B(n_690), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_41), .A2(n_87), .B1(n_514), .B2(n_553), .C(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g1382 ( .A(n_42), .Y(n_1382) );
OAI221xp5_ASAP7_75t_L g1398 ( .A1(n_42), .A2(n_302), .B1(n_1399), .B2(n_1400), .C(n_1401), .Y(n_1398) );
INVx1_ASAP7_75t_L g1489 ( .A(n_43), .Y(n_1489) );
CKINVDCx5p33_ASAP7_75t_R g1008 ( .A(n_44), .Y(n_1008) );
INVxp33_ASAP7_75t_SL g1110 ( .A(n_45), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_45), .A2(n_156), .B1(n_441), .B2(n_790), .Y(n_1130) );
AOI22xp33_ASAP7_75t_SL g1261 ( .A1(n_46), .A2(n_105), .B1(n_765), .B2(n_1262), .Y(n_1261) );
AOI22xp33_ASAP7_75t_SL g1285 ( .A1(n_46), .A2(n_180), .B1(n_1117), .B2(n_1286), .Y(n_1285) );
AOI221xp5_ASAP7_75t_L g1269 ( .A1(n_47), .A2(n_215), .B1(n_446), .B2(n_765), .C(n_1270), .Y(n_1269) );
OAI21xp33_ASAP7_75t_SL g1283 ( .A1(n_47), .A2(n_732), .B(n_1284), .Y(n_1283) );
OAI222xp33_ASAP7_75t_L g894 ( .A1(n_48), .A2(n_177), .B1(n_279), .B2(n_895), .C1(n_897), .C2(n_899), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_48), .A2(n_177), .B1(n_925), .B2(n_926), .C(n_927), .Y(n_924) );
CKINVDCx16_ASAP7_75t_R g1368 ( .A(n_49), .Y(n_1368) );
INVx1_ASAP7_75t_L g1069 ( .A(n_50), .Y(n_1069) );
CKINVDCx5p33_ASAP7_75t_R g934 ( .A(n_51), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_52), .A2(n_332), .B1(n_552), .B2(n_1117), .Y(n_1116) );
AOI221xp5_ASAP7_75t_L g1134 ( .A1(n_52), .A2(n_298), .B1(n_598), .B2(n_610), .C(n_1135), .Y(n_1134) );
AOI221xp5_ASAP7_75t_L g1163 ( .A1(n_53), .A2(n_172), .B1(n_608), .B2(n_609), .C(n_610), .Y(n_1163) );
INVxp33_ASAP7_75t_SL g1184 ( .A(n_53), .Y(n_1184) );
CKINVDCx5p33_ASAP7_75t_R g1326 ( .A(n_54), .Y(n_1326) );
INVx1_ASAP7_75t_L g1150 ( .A(n_55), .Y(n_1150) );
INVx1_ASAP7_75t_L g1616 ( .A(n_56), .Y(n_1616) );
OAI221xp5_ASAP7_75t_L g1909 ( .A1(n_58), .A2(n_112), .B1(n_520), .B2(n_531), .C(n_1910), .Y(n_1909) );
OAI221xp5_ASAP7_75t_SL g1932 ( .A1(n_58), .A2(n_112), .B1(n_776), .B2(n_777), .C(n_1933), .Y(n_1932) );
INVx1_ASAP7_75t_L g1622 ( .A(n_59), .Y(n_1622) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_60), .Y(n_750) );
XOR2xp5_ASAP7_75t_L g1144 ( .A(n_61), .B(n_1145), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1506 ( .A1(n_62), .A2(n_217), .B1(n_883), .B2(n_1262), .Y(n_1506) );
OAI22xp5_ASAP7_75t_L g1552 ( .A1(n_62), .A2(n_217), .B1(n_1553), .B2(n_1555), .Y(n_1552) );
INVxp67_ASAP7_75t_L g1423 ( .A(n_63), .Y(n_1423) );
AOI22xp5_ASAP7_75t_L g1727 ( .A1(n_63), .A2(n_334), .B1(n_1669), .B2(n_1691), .Y(n_1727) );
INVx1_ASAP7_75t_L g1356 ( .A(n_65), .Y(n_1356) );
AOI22xp33_ASAP7_75t_L g1390 ( .A1(n_66), .A2(n_221), .B1(n_1380), .B2(n_1391), .Y(n_1390) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_66), .A2(n_221), .B1(n_1286), .B2(n_1409), .Y(n_1408) );
OAI221xp5_ASAP7_75t_L g676 ( .A1(n_67), .A2(n_141), .B1(n_671), .B2(n_677), .C(n_678), .Y(n_676) );
INVx1_ASAP7_75t_L g726 ( .A(n_67), .Y(n_726) );
INVxp67_ASAP7_75t_L g1441 ( .A(n_68), .Y(n_1441) );
AOI22xp33_ASAP7_75t_L g1464 ( .A1(n_68), .A2(n_102), .B1(n_700), .B2(n_1022), .Y(n_1464) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_69), .A2(n_222), .B1(n_636), .B2(n_638), .C(n_640), .Y(n_635) );
INVx1_ASAP7_75t_L g1598 ( .A(n_71), .Y(n_1598) );
CKINVDCx5p33_ASAP7_75t_R g747 ( .A(n_72), .Y(n_747) );
AOI21xp33_ASAP7_75t_L g443 ( .A1(n_73), .A2(n_444), .B(n_446), .Y(n_443) );
INVxp33_ASAP7_75t_L g507 ( .A(n_73), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_74), .A2(n_216), .B1(n_837), .B2(n_839), .Y(n_836) );
INVxp67_ASAP7_75t_SL g860 ( .A(n_74), .Y(n_860) );
XOR2x2_ASAP7_75t_L g1469 ( .A(n_75), .B(n_1470), .Y(n_1469) );
INVxp33_ASAP7_75t_L g1606 ( .A(n_76), .Y(n_1606) );
AOI21xp33_ASAP7_75t_L g1634 ( .A1(n_76), .A2(n_700), .B(n_701), .Y(n_1634) );
INVxp33_ASAP7_75t_L g1484 ( .A(n_77), .Y(n_1484) );
INVx1_ASAP7_75t_L g1446 ( .A(n_78), .Y(n_1446) );
INVx1_ASAP7_75t_L g842 ( .A(n_79), .Y(n_842) );
AOI22x1_ASAP7_75t_L g1256 ( .A1(n_80), .A2(n_1257), .B1(n_1305), .B2(n_1306), .Y(n_1256) );
INVxp67_ASAP7_75t_L g1305 ( .A(n_80), .Y(n_1305) );
INVxp33_ASAP7_75t_L g1607 ( .A(n_81), .Y(n_1607) );
XNOR2x2_ASAP7_75t_L g1307 ( .A(n_82), .B(n_1308), .Y(n_1307) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_83), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g954 ( .A(n_84), .Y(n_954) );
AOI221xp5_ASAP7_75t_L g1563 ( .A1(n_85), .A2(n_352), .B1(n_446), .B2(n_765), .C(n_834), .Y(n_1563) );
INVxp33_ASAP7_75t_L g1582 ( .A(n_85), .Y(n_1582) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_86), .A2(n_182), .B1(n_553), .B2(n_945), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_86), .A2(n_182), .B1(n_818), .B2(n_975), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_87), .A2(n_245), .B1(n_588), .B2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_88), .A2(n_181), .B1(n_613), .B2(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g651 ( .A(n_88), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g1065 ( .A1(n_89), .A2(n_100), .B1(n_552), .B2(n_1062), .Y(n_1065) );
INVx1_ASAP7_75t_L g1097 ( .A(n_89), .Y(n_1097) );
INVxp33_ASAP7_75t_SL g1395 ( .A(n_90), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g1413 ( .A1(n_90), .A2(n_348), .B1(n_1286), .B2(n_1411), .Y(n_1413) );
AOI22xp33_ASAP7_75t_L g1571 ( .A1(n_91), .A2(n_303), .B1(n_604), .B2(n_1572), .Y(n_1571) );
INVxp67_ASAP7_75t_SL g1593 ( .A(n_91), .Y(n_1593) );
CKINVDCx5p33_ASAP7_75t_R g1010 ( .A(n_92), .Y(n_1010) );
XNOR2xp5_ASAP7_75t_L g1956 ( .A(n_93), .B(n_1901), .Y(n_1956) );
AOI22xp33_ASAP7_75t_SL g1564 ( .A1(n_94), .A2(n_235), .B1(n_603), .B2(n_784), .Y(n_1564) );
INVxp33_ASAP7_75t_SL g1585 ( .A(n_94), .Y(n_1585) );
OR2x2_ASAP7_75t_L g395 ( .A(n_95), .B(n_396), .Y(n_395) );
BUFx2_ASAP7_75t_L g399 ( .A(n_95), .Y(n_399) );
BUFx2_ASAP7_75t_L g487 ( .A(n_95), .Y(n_487) );
INVx1_ASAP7_75t_L g499 ( .A(n_95), .Y(n_499) );
AOI22xp33_ASAP7_75t_SL g946 ( .A1(n_96), .A2(n_110), .B1(n_937), .B2(n_939), .Y(n_946) );
INVx1_ASAP7_75t_L g973 ( .A(n_96), .Y(n_973) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_97), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_98), .A2(n_237), .B1(n_456), .B2(n_459), .C(n_463), .Y(n_455) );
INVxp67_ASAP7_75t_SL g550 ( .A(n_98), .Y(n_550) );
INVx1_ASAP7_75t_L g998 ( .A(n_99), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_99), .A2(n_283), .B1(n_1020), .B2(n_1021), .Y(n_1019) );
INVx1_ASAP7_75t_L g1072 ( .A(n_100), .Y(n_1072) );
AOI221xp5_ASAP7_75t_SL g597 ( .A1(n_101), .A2(n_107), .B1(n_446), .B2(n_598), .C(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g630 ( .A(n_101), .Y(n_630) );
INVxp33_ASAP7_75t_L g1436 ( .A(n_102), .Y(n_1436) );
INVx1_ASAP7_75t_L g592 ( .A(n_103), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g816 ( .A1(n_104), .A2(n_128), .B1(n_817), .B2(n_819), .C(n_820), .Y(n_816) );
INVxp33_ASAP7_75t_L g848 ( .A(n_104), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g1287 ( .A1(n_105), .A2(n_119), .B1(n_1115), .B2(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1920 ( .A(n_106), .Y(n_1920) );
INVx1_ASAP7_75t_L g627 ( .A(n_107), .Y(n_627) );
XOR2x2_ASAP7_75t_L g662 ( .A(n_108), .B(n_663), .Y(n_662) );
INVxp67_ASAP7_75t_SL g1619 ( .A(n_109), .Y(n_1619) );
AOI221xp5_ASAP7_75t_L g1638 ( .A1(n_109), .A2(n_311), .B1(n_690), .B2(n_833), .C(n_1639), .Y(n_1638) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_110), .B(n_478), .Y(n_959) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_111), .A2(n_236), .B1(n_394), .B2(n_734), .Y(n_733) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_111), .Y(n_794) );
OA22x2_ASAP7_75t_L g806 ( .A1(n_113), .A2(n_807), .B1(n_808), .B2(n_873), .Y(n_806) );
CKINVDCx16_ASAP7_75t_R g873 ( .A(n_113), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_114), .Y(n_1006) );
INVx1_ASAP7_75t_L g1453 ( .A(n_115), .Y(n_1453) );
CKINVDCx5p33_ASAP7_75t_R g1929 ( .A(n_116), .Y(n_1929) );
INVxp67_ASAP7_75t_L g1432 ( .A(n_117), .Y(n_1432) );
AOI22xp33_ASAP7_75t_L g1459 ( .A1(n_117), .A2(n_147), .B1(n_614), .B2(n_898), .Y(n_1459) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_118), .A2(n_265), .B1(n_441), .B2(n_698), .Y(n_697) );
OAI211xp5_ASAP7_75t_L g702 ( .A1(n_118), .A2(n_703), .B(n_705), .C(n_707), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g1264 ( .A1(n_119), .A2(n_180), .B1(n_608), .B2(n_1265), .C(n_1267), .Y(n_1264) );
OAI22xp5_ASAP7_75t_L g1151 ( .A1(n_120), .A2(n_187), .B1(n_427), .B2(n_1152), .Y(n_1151) );
OAI221xp5_ASAP7_75t_L g1193 ( .A1(n_120), .A2(n_187), .B1(n_737), .B2(n_738), .C(n_989), .Y(n_1193) );
INVx1_ASAP7_75t_L g1467 ( .A(n_121), .Y(n_1467) );
OAI22xp33_ASAP7_75t_SL g1332 ( .A1(n_122), .A2(n_158), .B1(n_668), .B2(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1357 ( .A(n_122), .Y(n_1357) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_123), .A2(n_192), .B1(n_608), .B2(n_609), .C(n_610), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_123), .A2(n_181), .B1(n_646), .B2(n_648), .C(n_650), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g1711 ( .A1(n_124), .A2(n_328), .B1(n_1669), .B2(n_1691), .Y(n_1711) );
CKINVDCx5p33_ASAP7_75t_R g1323 ( .A(n_125), .Y(n_1323) );
AOI22xp33_ASAP7_75t_SL g1118 ( .A1(n_126), .A2(n_345), .B1(n_1000), .B2(n_1117), .Y(n_1118) );
INVxp33_ASAP7_75t_L g1140 ( .A(n_126), .Y(n_1140) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_127), .Y(n_1013) );
INVxp33_ASAP7_75t_L g851 ( .A(n_128), .Y(n_851) );
OAI222xp33_ASAP7_75t_L g900 ( .A1(n_129), .A2(n_209), .B1(n_344), .B2(n_616), .C1(n_901), .C2(n_902), .Y(n_900) );
INVx1_ASAP7_75t_L g915 ( .A(n_129), .Y(n_915) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_130), .A2(n_320), .B1(n_670), .B2(n_671), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_130), .A2(n_191), .B1(n_628), .B2(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g1431 ( .A(n_131), .Y(n_1431) );
AOI221xp5_ASAP7_75t_L g1458 ( .A1(n_131), .A2(n_201), .B1(n_444), .B2(n_446), .C(n_834), .Y(n_1458) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_132), .A2(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g708 ( .A(n_132), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_133), .A2(n_191), .B1(n_667), .B2(n_668), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_133), .A2(n_320), .B1(n_494), .B2(n_716), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g1700 ( .A1(n_134), .A2(n_137), .B1(n_1701), .B2(n_1704), .Y(n_1700) );
INVx1_ASAP7_75t_L g997 ( .A(n_135), .Y(n_997) );
AOI221xp5_ASAP7_75t_L g1388 ( .A1(n_136), .A2(n_312), .B1(n_609), .B2(n_1267), .C(n_1389), .Y(n_1388) );
AOI22xp33_ASAP7_75t_L g1410 ( .A1(n_136), .A2(n_312), .B1(n_1411), .B2(n_1412), .Y(n_1410) );
AOI22xp5_ASAP7_75t_L g1706 ( .A1(n_138), .A2(n_343), .B1(n_1661), .B2(n_1707), .Y(n_1706) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_139), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g1433 ( .A1(n_140), .A2(n_184), .B1(n_520), .B2(n_737), .C(n_738), .Y(n_1433) );
OAI22xp5_ASAP7_75t_L g1460 ( .A1(n_140), .A2(n_184), .B1(n_1128), .B2(n_1336), .Y(n_1460) );
INVx1_ASAP7_75t_L g706 ( .A(n_141), .Y(n_706) );
INVx1_ASAP7_75t_L g595 ( .A(n_142), .Y(n_595) );
INVx1_ASAP7_75t_L g1159 ( .A(n_143), .Y(n_1159) );
CKINVDCx5p33_ASAP7_75t_R g757 ( .A(n_144), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g885 ( .A1(n_145), .A2(n_310), .B1(n_465), .B2(n_886), .C(n_887), .Y(n_885) );
INVx1_ASAP7_75t_L g923 ( .A(n_145), .Y(n_923) );
AO221x2_ASAP7_75t_L g1735 ( .A1(n_146), .A2(n_226), .B1(n_1661), .B2(n_1669), .C(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1900 ( .A(n_146), .Y(n_1900) );
AOI22xp33_ASAP7_75t_L g1951 ( .A1(n_146), .A2(n_1952), .B1(n_1955), .B2(n_1957), .Y(n_1951) );
INVxp67_ASAP7_75t_L g1428 ( .A(n_147), .Y(n_1428) );
INVxp33_ASAP7_75t_SL g1394 ( .A(n_148), .Y(n_1394) );
AOI22xp33_ASAP7_75t_L g1414 ( .A1(n_148), .A2(n_290), .B1(n_1409), .B2(n_1412), .Y(n_1414) );
INVx1_ASAP7_75t_L g1666 ( .A(n_149), .Y(n_1666) );
INVx1_ASAP7_75t_L g1047 ( .A(n_150), .Y(n_1047) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_150), .A2(n_264), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
XNOR2x1_ASAP7_75t_L g1098 ( .A(n_151), .B(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1667 ( .A(n_151), .Y(n_1667) );
INVx1_ASAP7_75t_L g831 ( .A(n_152), .Y(n_831) );
INVx1_ASAP7_75t_L g1169 ( .A(n_153), .Y(n_1169) );
CKINVDCx5p33_ASAP7_75t_R g1628 ( .A(n_154), .Y(n_1628) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_155), .A2(n_315), .B1(n_939), .B2(n_1060), .Y(n_1059) );
INVxp33_ASAP7_75t_SL g1105 ( .A(n_156), .Y(n_1105) );
AOI221xp5_ASAP7_75t_L g832 ( .A1(n_157), .A2(n_231), .B1(n_688), .B2(n_833), .C(n_835), .Y(n_832) );
INVxp67_ASAP7_75t_SL g865 ( .A(n_157), .Y(n_865) );
INVx1_ASAP7_75t_L g1351 ( .A(n_158), .Y(n_1351) );
AOI22xp5_ASAP7_75t_L g1726 ( .A1(n_159), .A2(n_353), .B1(n_1701), .B2(n_1704), .Y(n_1726) );
INVx1_ASAP7_75t_L g962 ( .A(n_160), .Y(n_962) );
XOR2x1_ASAP7_75t_L g1040 ( .A(n_161), .B(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1604 ( .A(n_162), .Y(n_1604) );
NAND2xp5_ASAP7_75t_L g1635 ( .A(n_162), .B(n_1384), .Y(n_1635) );
INVx1_ASAP7_75t_L g1923 ( .A(n_163), .Y(n_1923) );
INVx1_ASAP7_75t_L g1495 ( .A(n_164), .Y(n_1495) );
AOI221xp5_ASAP7_75t_L g1153 ( .A1(n_165), .A2(n_210), .B1(n_604), .B2(n_1154), .C(n_1156), .Y(n_1153) );
INVxp33_ASAP7_75t_L g1196 ( .A(n_165), .Y(n_1196) );
INVx1_ASAP7_75t_L g1664 ( .A(n_166), .Y(n_1664) );
NAND2xp5_ASAP7_75t_L g1683 ( .A(n_166), .B(n_1677), .Y(n_1683) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_167), .A2(n_252), .B1(n_603), .B2(n_604), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_167), .A2(n_252), .B1(n_624), .B2(n_625), .C(n_626), .Y(n_623) );
INVxp33_ASAP7_75t_L g1139 ( .A(n_168), .Y(n_1139) );
AOI22xp33_ASAP7_75t_SL g1501 ( .A1(n_169), .A2(n_204), .B1(n_819), .B2(n_1502), .Y(n_1501) );
INVxp67_ASAP7_75t_SL g1540 ( .A(n_169), .Y(n_1540) );
INVx1_ASAP7_75t_L g1220 ( .A(n_170), .Y(n_1220) );
INVx2_ASAP7_75t_L g378 ( .A(n_171), .Y(n_378) );
INVxp67_ASAP7_75t_L g1174 ( .A(n_172), .Y(n_1174) );
AOI221xp5_ASAP7_75t_L g1569 ( .A1(n_173), .A2(n_333), .B1(n_415), .B2(n_610), .C(n_1570), .Y(n_1569) );
INVxp33_ASAP7_75t_SL g1590 ( .A(n_173), .Y(n_1590) );
INVx1_ASAP7_75t_L g1934 ( .A(n_174), .Y(n_1934) );
BUFx3_ASAP7_75t_L g408 ( .A(n_175), .Y(n_408) );
INVx1_ASAP7_75t_L g437 ( .A(n_175), .Y(n_437) );
INVx1_ASAP7_75t_L g1272 ( .A(n_176), .Y(n_1272) );
INVx1_ASAP7_75t_L g1737 ( .A(n_178), .Y(n_1737) );
INVx1_ASAP7_75t_L g1478 ( .A(n_179), .Y(n_1478) );
INVx1_ASAP7_75t_L g1624 ( .A(n_183), .Y(n_1624) );
CKINVDCx5p33_ASAP7_75t_R g986 ( .A(n_185), .Y(n_986) );
INVxp33_ASAP7_75t_L g1229 ( .A(n_186), .Y(n_1229) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_186), .A2(n_300), .B1(n_1239), .B2(n_1240), .Y(n_1238) );
INVx1_ASAP7_75t_L g1107 ( .A(n_188), .Y(n_1107) );
CKINVDCx5p33_ASAP7_75t_R g1322 ( .A(n_189), .Y(n_1322) );
INVx1_ASAP7_75t_L g1168 ( .A(n_190), .Y(n_1168) );
INVx1_ASAP7_75t_L g652 ( .A(n_192), .Y(n_652) );
INVxp67_ASAP7_75t_L g1913 ( .A(n_193), .Y(n_1913) );
AOI22xp33_ASAP7_75t_L g1943 ( .A1(n_193), .A2(n_331), .B1(n_1240), .B2(n_1391), .Y(n_1943) );
OAI22xp33_ASAP7_75t_R g827 ( .A1(n_194), .A2(n_357), .B1(n_427), .B2(n_776), .Y(n_827) );
OAI221xp5_ASAP7_75t_L g853 ( .A1(n_194), .A2(n_357), .B1(n_520), .B2(n_854), .C(n_855), .Y(n_853) );
OAI221xp5_ASAP7_75t_SL g421 ( .A1(n_195), .A2(n_350), .B1(n_422), .B2(n_427), .C(n_431), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g519 ( .A1(n_195), .A2(n_350), .B1(n_520), .B2(n_527), .C(n_530), .Y(n_519) );
INVx1_ASAP7_75t_L g1659 ( .A(n_196), .Y(n_1659) );
CKINVDCx5p33_ASAP7_75t_R g984 ( .A(n_197), .Y(n_984) );
INVx1_ASAP7_75t_L g841 ( .A(n_198), .Y(n_841) );
INVx1_ASAP7_75t_L g1907 ( .A(n_199), .Y(n_1907) );
INVxp67_ASAP7_75t_SL g1273 ( .A(n_200), .Y(n_1273) );
INVxp67_ASAP7_75t_L g1429 ( .A(n_201), .Y(n_1429) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_202), .A2(n_337), .B1(n_884), .B2(n_1165), .Y(n_1164) );
INVxp67_ASAP7_75t_SL g1178 ( .A(n_202), .Y(n_1178) );
INVx1_ASAP7_75t_L g594 ( .A(n_203), .Y(n_594) );
INVxp67_ASAP7_75t_SL g1545 ( .A(n_204), .Y(n_1545) );
INVx1_ASAP7_75t_L g1162 ( .A(n_205), .Y(n_1162) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_207), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g1513 ( .A(n_208), .Y(n_1513) );
INVx1_ASAP7_75t_L g907 ( .A(n_209), .Y(n_907) );
INVxp33_ASAP7_75t_L g1199 ( .A(n_210), .Y(n_1199) );
INVx1_ASAP7_75t_L g1147 ( .A(n_211), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_212), .A2(n_297), .B1(n_883), .B2(n_884), .Y(n_882) );
INVx1_ASAP7_75t_L g913 ( .A(n_212), .Y(n_913) );
INVx1_ASAP7_75t_L g1250 ( .A(n_213), .Y(n_1250) );
INVx1_ASAP7_75t_L g1055 ( .A(n_214), .Y(n_1055) );
AOI221xp5_ASAP7_75t_L g1077 ( .A1(n_214), .A2(n_301), .B1(n_603), .B2(n_1022), .C(n_1078), .Y(n_1077) );
INVxp33_ASAP7_75t_SL g1295 ( .A(n_215), .Y(n_1295) );
INVxp67_ASAP7_75t_SL g867 ( .A(n_216), .Y(n_867) );
INVx1_ASAP7_75t_L g1738 ( .A(n_218), .Y(n_1738) );
INVx1_ASAP7_75t_L g480 ( .A(n_219), .Y(n_480) );
INVx1_ASAP7_75t_L g403 ( .A(n_220), .Y(n_403) );
INVx1_ASAP7_75t_L g448 ( .A(n_220), .Y(n_448) );
INVx1_ASAP7_75t_L g591 ( .A(n_222), .Y(n_591) );
INVxp33_ASAP7_75t_SL g1109 ( .A(n_223), .Y(n_1109) );
AOI21xp33_ASAP7_75t_L g1131 ( .A1(n_223), .A2(n_826), .B(n_964), .Y(n_1131) );
INVx1_ASAP7_75t_L g1621 ( .A(n_224), .Y(n_1621) );
INVx1_ASAP7_75t_L g1695 ( .A(n_225), .Y(n_1695) );
INVx1_ASAP7_75t_L g1565 ( .A(n_227), .Y(n_1565) );
CKINVDCx5p33_ASAP7_75t_R g694 ( .A(n_228), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g1319 ( .A1(n_229), .A2(n_321), .B1(n_688), .B2(n_1320), .C(n_1321), .Y(n_1319) );
INVx1_ASAP7_75t_L g1361 ( .A(n_229), .Y(n_1361) );
AOI22xp33_ASAP7_75t_SL g1505 ( .A1(n_230), .A2(n_285), .B1(n_837), .B2(n_1502), .Y(n_1505) );
OAI211xp5_ASAP7_75t_SL g1521 ( .A1(n_230), .A2(n_1522), .B(n_1527), .C(n_1531), .Y(n_1521) );
INVxp67_ASAP7_75t_SL g861 ( .A(n_231), .Y(n_861) );
XNOR2x1_ASAP7_75t_L g977 ( .A(n_232), .B(n_978), .Y(n_977) );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_233), .A2(n_318), .B1(n_446), .B2(n_598), .C(n_600), .Y(n_881) );
INVx1_ASAP7_75t_L g911 ( .A(n_233), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g1710 ( .A1(n_234), .A2(n_293), .B1(n_1701), .B2(n_1704), .Y(n_1710) );
INVxp33_ASAP7_75t_L g1581 ( .A(n_235), .Y(n_1581) );
INVx1_ASAP7_75t_L g545 ( .A(n_237), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g933 ( .A(n_238), .Y(n_933) );
INVx1_ASAP7_75t_L g982 ( .A(n_239), .Y(n_982) );
INVxp67_ASAP7_75t_L g1440 ( .A(n_240), .Y(n_1440) );
AOI221xp5_ASAP7_75t_L g1462 ( .A1(n_240), .A2(n_253), .B1(n_440), .B2(n_1318), .C(n_1463), .Y(n_1462) );
INVxp33_ASAP7_75t_L g1211 ( .A(n_241), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g1233 ( .A1(n_241), .A2(n_270), .B1(n_458), .B2(n_610), .C(n_887), .Y(n_1233) );
INVx1_ASAP7_75t_L g824 ( .A(n_242), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_243), .A2(n_305), .B1(n_468), .B2(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g539 ( .A(n_243), .Y(n_539) );
INVx1_ASAP7_75t_L g814 ( .A(n_244), .Y(n_814) );
INVx1_ASAP7_75t_L g721 ( .A(n_245), .Y(n_721) );
CKINVDCx16_ASAP7_75t_R g1692 ( .A(n_246), .Y(n_1692) );
OAI211xp5_ASAP7_75t_SL g1274 ( .A1(n_247), .A2(n_1275), .B(n_1276), .C(n_1280), .Y(n_1274) );
INVx1_ASAP7_75t_L g1302 ( .A(n_247), .Y(n_1302) );
INVx1_ASAP7_75t_L g957 ( .A(n_248), .Y(n_957) );
OAI211xp5_ASAP7_75t_L g971 ( .A1(n_248), .A2(n_616), .B(n_972), .C(n_976), .Y(n_971) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_249), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_250), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_251), .A2(n_288), .B1(n_1060), .B2(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1096 ( .A(n_251), .Y(n_1096) );
INVxp33_ASAP7_75t_L g1437 ( .A(n_253), .Y(n_1437) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_254), .A2(n_260), .B1(n_440), .B2(n_441), .Y(n_439) );
INVxp33_ASAP7_75t_L g512 ( .A(n_254), .Y(n_512) );
XNOR2x1_ASAP7_75t_L g877 ( .A(n_255), .B(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g1921 ( .A(n_256), .Y(n_1921) );
BUFx3_ASAP7_75t_L g410 ( .A(n_257), .Y(n_410) );
INVx1_ASAP7_75t_L g417 ( .A(n_257), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g745 ( .A(n_258), .Y(n_745) );
CKINVDCx5p33_ASAP7_75t_R g1316 ( .A(n_259), .Y(n_1316) );
INVxp33_ASAP7_75t_L g491 ( .A(n_260), .Y(n_491) );
INVx1_ASAP7_75t_L g575 ( .A(n_261), .Y(n_575) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_262), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_262), .B(n_341), .Y(n_396) );
AND2x2_ASAP7_75t_L g500 ( .A(n_262), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g574 ( .A(n_262), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g1003 ( .A(n_263), .Y(n_1003) );
INVx1_ASAP7_75t_L g1046 ( .A(n_264), .Y(n_1046) );
INVx1_ASAP7_75t_L g711 ( .A(n_265), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g1383 ( .A1(n_266), .A2(n_1245), .B(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1403 ( .A(n_266), .Y(n_1403) );
OAI332xp33_ASAP7_75t_L g739 ( .A1(n_267), .A2(n_533), .A3(n_570), .B1(n_740), .B2(n_744), .B3(n_749), .C1(n_756), .C2(n_761), .Y(n_739) );
INVx1_ASAP7_75t_L g798 ( .A(n_267), .Y(n_798) );
INVx1_ASAP7_75t_L g1678 ( .A(n_268), .Y(n_1678) );
INVx1_ASAP7_75t_L g1158 ( .A(n_269), .Y(n_1158) );
INVxp67_ASAP7_75t_L g1206 ( .A(n_270), .Y(n_1206) );
INVx1_ASAP7_75t_L g1575 ( .A(n_271), .Y(n_1575) );
INVx1_ASAP7_75t_L g1696 ( .A(n_273), .Y(n_1696) );
INVx2_ASAP7_75t_L g405 ( .A(n_274), .Y(n_405) );
OR2x2_ASAP7_75t_L g419 ( .A(n_274), .B(n_403), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_275), .Y(n_742) );
INVx1_ASAP7_75t_L g1671 ( .A(n_276), .Y(n_1671) );
INVx1_ASAP7_75t_L g1444 ( .A(n_277), .Y(n_1444) );
INVxp67_ASAP7_75t_L g1917 ( .A(n_278), .Y(n_1917) );
AOI221xp5_ASAP7_75t_L g1940 ( .A1(n_278), .A2(n_329), .B1(n_835), .B2(n_1941), .C(n_1942), .Y(n_1940) );
INVx1_ASAP7_75t_L g928 ( .A(n_279), .Y(n_928) );
CKINVDCx16_ASAP7_75t_R g580 ( .A(n_280), .Y(n_580) );
INVx1_ASAP7_75t_L g1576 ( .A(n_281), .Y(n_1576) );
INVxp67_ASAP7_75t_SL g1277 ( .A(n_282), .Y(n_1277) );
OAI211xp5_ASAP7_75t_SL g1289 ( .A1(n_282), .A2(n_759), .B(n_1290), .C(n_1292), .Y(n_1289) );
INVx1_ASAP7_75t_L g992 ( .A(n_283), .Y(n_992) );
INVx1_ASAP7_75t_L g454 ( .A(n_284), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g1536 ( .A1(n_285), .A2(n_1537), .B1(n_1539), .B2(n_1544), .C(n_1551), .Y(n_1536) );
INVx1_ASAP7_75t_L g1720 ( .A(n_286), .Y(n_1720) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_287), .A2(n_316), .B1(n_784), .B2(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g921 ( .A(n_287), .Y(n_921) );
INVx1_ASAP7_75t_L g1085 ( .A(n_288), .Y(n_1085) );
CKINVDCx5p33_ASAP7_75t_R g1054 ( .A(n_289), .Y(n_1054) );
INVxp67_ASAP7_75t_SL g1387 ( .A(n_290), .Y(n_1387) );
INVx1_ASAP7_75t_L g1924 ( .A(n_291), .Y(n_1924) );
AOI221xp5_ASAP7_75t_L g1379 ( .A1(n_292), .A2(n_302), .B1(n_609), .B2(n_1380), .C(n_1381), .Y(n_1379) );
INVxp33_ASAP7_75t_L g1402 ( .A(n_292), .Y(n_1402) );
INVx1_ASAP7_75t_L g1596 ( .A(n_294), .Y(n_1596) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_295), .Y(n_811) );
INVx1_ASAP7_75t_L g950 ( .A(n_296), .Y(n_950) );
AOI21xp5_ASAP7_75t_L g968 ( .A1(n_296), .A2(n_686), .B(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g909 ( .A(n_297), .Y(n_909) );
INVxp33_ASAP7_75t_L g1296 ( .A(n_299), .Y(n_1296) );
INVxp33_ASAP7_75t_L g1225 ( .A(n_300), .Y(n_1225) );
INVx1_ASAP7_75t_L g1050 ( .A(n_301), .Y(n_1050) );
INVxp33_ASAP7_75t_L g1589 ( .A(n_303), .Y(n_1589) );
CKINVDCx5p33_ASAP7_75t_R g1315 ( .A(n_304), .Y(n_1315) );
INVx1_ASAP7_75t_L g554 ( .A(n_305), .Y(n_554) );
INVx1_ASAP7_75t_L g1217 ( .A(n_306), .Y(n_1217) );
INVxp67_ASAP7_75t_SL g1102 ( .A(n_307), .Y(n_1102) );
OAI221xp5_ASAP7_75t_L g1127 ( .A1(n_307), .A2(n_335), .B1(n_422), .B2(n_1128), .C(n_1129), .Y(n_1127) );
INVx1_ASAP7_75t_L g1626 ( .A(n_308), .Y(n_1626) );
INVx1_ASAP7_75t_L g953 ( .A(n_309), .Y(n_953) );
AOI221xp5_ASAP7_75t_L g918 ( .A1(n_310), .A2(n_316), .B1(n_636), .B2(n_919), .C(n_920), .Y(n_918) );
INVxp33_ASAP7_75t_L g1614 ( .A(n_311), .Y(n_1614) );
INVx1_ASAP7_75t_L g1715 ( .A(n_313), .Y(n_1715) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_315), .A2(n_317), .B1(n_817), .B2(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g917 ( .A(n_318), .Y(n_917) );
CKINVDCx5p33_ASAP7_75t_R g893 ( .A(n_319), .Y(n_893) );
INVx1_ASAP7_75t_L g1363 ( .A(n_321), .Y(n_1363) );
INVx1_ASAP7_75t_L g1452 ( .A(n_322), .Y(n_1452) );
INVx1_ASAP7_75t_L g1577 ( .A(n_323), .Y(n_1577) );
INVx1_ASAP7_75t_L g432 ( .A(n_324), .Y(n_432) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_325), .Y(n_368) );
AND3x2_ASAP7_75t_L g1665 ( .A(n_325), .B(n_366), .C(n_1666), .Y(n_1665) );
NAND2xp5_ASAP7_75t_L g1675 ( .A(n_325), .B(n_366), .Y(n_1675) );
INVx1_ASAP7_75t_L g1247 ( .A(n_326), .Y(n_1247) );
INVx2_ASAP7_75t_L g379 ( .A(n_327), .Y(n_379) );
INVxp67_ASAP7_75t_SL g1918 ( .A(n_329), .Y(n_1918) );
CKINVDCx5p33_ASAP7_75t_R g1052 ( .A(n_330), .Y(n_1052) );
INVxp33_ASAP7_75t_SL g1915 ( .A(n_331), .Y(n_1915) );
INVxp67_ASAP7_75t_SL g1592 ( .A(n_333), .Y(n_1592) );
INVxp67_ASAP7_75t_SL g1103 ( .A(n_335), .Y(n_1103) );
AOI22x1_ASAP7_75t_L g1200 ( .A1(n_336), .A2(n_1201), .B1(n_1202), .B2(n_1251), .Y(n_1200) );
INVx1_ASAP7_75t_L g1251 ( .A(n_336), .Y(n_1251) );
INVxp33_ASAP7_75t_L g1182 ( .A(n_337), .Y(n_1182) );
CKINVDCx5p33_ASAP7_75t_R g741 ( .A(n_338), .Y(n_741) );
INVx1_ASAP7_75t_L g822 ( .A(n_339), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g1338 ( .A(n_340), .Y(n_1338) );
INVx1_ASAP7_75t_L g381 ( .A(n_341), .Y(n_381) );
INVx2_ASAP7_75t_L g501 ( .A(n_341), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g1337 ( .A(n_342), .Y(n_1337) );
INVx1_ASAP7_75t_L g906 ( .A(n_344), .Y(n_906) );
INVxp67_ASAP7_75t_L g1126 ( .A(n_345), .Y(n_1126) );
INVxp67_ASAP7_75t_SL g1550 ( .A(n_346), .Y(n_1550) );
INVxp33_ASAP7_75t_L g1210 ( .A(n_347), .Y(n_1210) );
INVxp67_ASAP7_75t_SL g1375 ( .A(n_348), .Y(n_1375) );
INVxp67_ASAP7_75t_SL g1417 ( .A(n_349), .Y(n_1417) );
INVx1_ASAP7_75t_L g1721 ( .A(n_351), .Y(n_1721) );
INVxp33_ASAP7_75t_L g1584 ( .A(n_352), .Y(n_1584) );
INVx1_ASAP7_75t_L g1279 ( .A(n_354), .Y(n_1279) );
INVx1_ASAP7_75t_L g1349 ( .A(n_355), .Y(n_1349) );
CKINVDCx5p33_ASAP7_75t_R g1372 ( .A(n_356), .Y(n_1372) );
INVx1_ASAP7_75t_L g476 ( .A(n_358), .Y(n_476) );
INVxp33_ASAP7_75t_SL g1906 ( .A(n_359), .Y(n_1906) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_382), .B(n_1653), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_364), .B(n_369), .Y(n_363) );
AND2x4_ASAP7_75t_L g1950 ( .A(n_364), .B(n_370), .Y(n_1950) );
NOR2xp33_ASAP7_75t_SL g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_SL g1954 ( .A(n_365), .Y(n_1954) );
NAND2xp5_ASAP7_75t_L g1964 ( .A(n_365), .B(n_367), .Y(n_1964) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g1953 ( .A(n_367), .B(n_1954), .Y(n_1953) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_375), .Y(n_370) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g644 ( .A(n_373), .B(n_381), .Y(n_644) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g534 ( .A(n_374), .B(n_535), .Y(n_534) );
OR2x6_ASAP7_75t_L g375 ( .A(n_376), .B(n_380), .Y(n_375) );
OR2x2_ASAP7_75t_L g394 ( .A(n_376), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g538 ( .A(n_376), .Y(n_538) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_376), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_376), .A2(n_682), .B1(n_721), .B2(n_722), .Y(n_720) );
INVx2_ASAP7_75t_SL g859 ( .A(n_376), .Y(n_859) );
BUFx2_ASAP7_75t_L g922 ( .A(n_376), .Y(n_922) );
OAI22xp33_ASAP7_75t_L g927 ( .A1(n_376), .A2(n_722), .B1(n_893), .B2(n_928), .Y(n_927) );
INVx2_ASAP7_75t_SL g1192 ( .A(n_376), .Y(n_1192) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
AND2x4_ASAP7_75t_L g496 ( .A(n_378), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g505 ( .A(n_378), .Y(n_505) );
AND2x2_ASAP7_75t_L g511 ( .A(n_378), .B(n_379), .Y(n_511) );
INVx2_ASAP7_75t_L g516 ( .A(n_378), .Y(n_516) );
INVx1_ASAP7_75t_L g544 ( .A(n_378), .Y(n_544) );
INVx2_ASAP7_75t_L g497 ( .A(n_379), .Y(n_497) );
INVx1_ASAP7_75t_L g518 ( .A(n_379), .Y(n_518) );
INVx1_ASAP7_75t_L g525 ( .A(n_379), .Y(n_525) );
INVx1_ASAP7_75t_L g543 ( .A(n_379), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_379), .B(n_516), .Y(n_549) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_1034), .B1(n_1650), .B2(n_1651), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g1652 ( .A(n_385), .Y(n_1652) );
AO22x2_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_805), .B2(n_1033), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
XNOR2x1_ASAP7_75t_L g387 ( .A(n_388), .B(n_576), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
XNOR2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_575), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_488), .Y(n_390) );
AOI21xp33_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_411), .B(n_412), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g1122 ( .A1(n_392), .A2(n_1123), .B1(n_1124), .B2(n_1141), .Y(n_1122) );
AOI21xp33_ASAP7_75t_L g1146 ( .A1(n_392), .A2(n_1147), .B(n_1148), .Y(n_1146) );
AOI22xp5_ASAP7_75t_L g1230 ( .A1(n_392), .A2(n_1123), .B1(n_1231), .B2(n_1250), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1560 ( .A1(n_392), .A2(n_1123), .B1(n_1561), .B2(n_1577), .Y(n_1560) );
INVx1_ASAP7_75t_L g1928 ( .A(n_392), .Y(n_1928) );
INVx5_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g810 ( .A(n_393), .Y(n_810) );
INVx1_ASAP7_75t_L g1012 ( .A(n_393), .Y(n_1012) );
INVx1_ASAP7_75t_L g1371 ( .A(n_393), .Y(n_1371) );
INVx2_ASAP7_75t_SL g1466 ( .A(n_393), .Y(n_1466) );
AND2x4_ASAP7_75t_L g393 ( .A(n_394), .B(n_397), .Y(n_393) );
INVx2_ASAP7_75t_L g653 ( .A(n_394), .Y(n_653) );
INVx3_ASAP7_75t_L g526 ( .A(n_395), .Y(n_526) );
INVx1_ASAP7_75t_L g1519 ( .A(n_396), .Y(n_1519) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x6_ASAP7_75t_L g1514 ( .A(n_398), .B(n_1515), .Y(n_1514) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
AND2x4_ASAP7_75t_L g1507 ( .A(n_399), .B(n_447), .Y(n_1507) );
INVx2_ASAP7_75t_L g616 ( .A(n_400), .Y(n_616) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_406), .Y(n_400) );
AND2x4_ASAP7_75t_L g423 ( .A(n_401), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g428 ( .A(n_401), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g473 ( .A(n_401), .Y(n_473) );
AND2x4_ASAP7_75t_L g593 ( .A(n_401), .B(n_424), .Y(n_593) );
BUFx2_ASAP7_75t_L g680 ( .A(n_401), .Y(n_680) );
AND2x4_ASAP7_75t_L g903 ( .A(n_401), .B(n_429), .Y(n_903) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_401), .B(n_429), .Y(n_1076) );
NAND2x1p5_ASAP7_75t_L g1494 ( .A(n_401), .B(n_571), .Y(n_1494) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_404), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g447 ( .A(n_404), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g466 ( .A(n_405), .B(n_448), .Y(n_466) );
INVx6_ASAP7_75t_L g445 ( .A(n_406), .Y(n_445) );
BUFx2_ASAP7_75t_L g700 ( .A(n_406), .Y(n_700) );
INVx2_ASAP7_75t_L g1094 ( .A(n_406), .Y(n_1094) );
AND2x4_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g430 ( .A(n_407), .Y(n_430) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g416 ( .A(n_408), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g453 ( .A(n_408), .B(n_410), .Y(n_453) );
INVx1_ASAP7_75t_L g426 ( .A(n_409), .Y(n_426) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g442 ( .A(n_410), .B(n_437), .Y(n_442) );
AOI31xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_449), .A3(n_475), .B(n_484), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_420), .B(n_421), .Y(n_413) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_414), .Y(n_815) );
AOI211xp5_ASAP7_75t_L g1023 ( .A1(n_414), .A2(n_1003), .B(n_1024), .C(n_1025), .Y(n_1023) );
AOI211xp5_ASAP7_75t_L g1071 ( .A1(n_414), .A2(n_1072), .B(n_1073), .C(n_1077), .Y(n_1071) );
AOI21xp33_ASAP7_75t_L g1125 ( .A1(n_414), .A2(n_1126), .B(n_1127), .Y(n_1125) );
AOI211xp5_ASAP7_75t_L g1149 ( .A1(n_414), .A2(n_1150), .B(n_1151), .C(n_1153), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_414), .A2(n_477), .B1(n_1216), .B2(n_1219), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1271 ( .A1(n_414), .A2(n_477), .B1(n_1272), .B2(n_1273), .Y(n_1271) );
INVx1_ASAP7_75t_L g1377 ( .A(n_414), .Y(n_1377) );
AOI221xp5_ASAP7_75t_L g1562 ( .A1(n_414), .A2(n_1563), .B1(n_1564), .B2(n_1565), .C(n_1566), .Y(n_1562) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .Y(n_414) );
BUFx3_ASAP7_75t_L g603 ( .A(n_415), .Y(n_603) );
INVx2_ASAP7_75t_SL g1640 ( .A(n_415), .Y(n_1640) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_416), .Y(n_440) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_416), .Y(n_458) );
BUFx2_ASAP7_75t_L g609 ( .A(n_416), .Y(n_609) );
INVx2_ASAP7_75t_SL g689 ( .A(n_416), .Y(n_689) );
BUFx3_ASAP7_75t_L g698 ( .A(n_416), .Y(n_698) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_416), .Y(n_790) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_416), .Y(n_886) );
BUFx2_ASAP7_75t_L g898 ( .A(n_416), .Y(n_898) );
INVx1_ASAP7_75t_L g438 ( .A(n_417), .Y(n_438) );
AND2x4_ASAP7_75t_L g451 ( .A(n_418), .B(n_452), .Y(n_451) );
AOI222xp33_ASAP7_75t_L g583 ( .A1(n_418), .A2(n_428), .B1(n_584), .B2(n_593), .C1(n_594), .C2(n_595), .Y(n_583) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_418), .A2(n_666), .B(n_669), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g892 ( .A1(n_418), .A2(n_477), .B1(n_893), .B2(n_894), .C(n_900), .Y(n_892) );
A2O1A1Ixp33_ASAP7_75t_L g972 ( .A1(n_418), .A2(n_834), .B(n_973), .C(n_974), .Y(n_972) );
OAI21xp33_ASAP7_75t_L g1329 ( .A1(n_418), .A2(n_1330), .B(n_1332), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_418), .B(n_458), .Y(n_1457) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g478 ( .A(n_419), .B(n_479), .Y(n_478) );
OR2x2_ASAP7_75t_L g482 ( .A(n_419), .B(n_483), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_SL g763 ( .A1(n_419), .A2(n_764), .B(n_769), .C(n_774), .Y(n_763) );
OR2x2_ASAP7_75t_L g1477 ( .A(n_419), .B(n_499), .Y(n_1477) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_420), .A2(n_480), .B1(n_556), .B2(n_559), .Y(n_555) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g901 ( .A(n_423), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_423), .A2(n_903), .B1(n_933), .B2(n_934), .Y(n_976) );
INVx4_ASAP7_75t_L g1336 ( .A(n_423), .Y(n_1336) );
INVxp67_ASAP7_75t_L g677 ( .A(n_424), .Y(n_677) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g1492 ( .A(n_425), .Y(n_1492) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g678 ( .A(n_429), .Y(n_678) );
INVx2_ASAP7_75t_L g778 ( .A(n_429), .Y(n_778) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI211xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B(n_439), .C(n_443), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_432), .A2(n_491), .B1(n_492), .B2(n_502), .Y(n_490) );
OAI211xp5_ASAP7_75t_L g1129 ( .A1(n_433), .A2(n_1107), .B(n_1130), .C(n_1131), .Y(n_1129) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_SL g671 ( .A(n_434), .Y(n_671) );
INVx1_ASAP7_75t_L g821 ( .A(n_434), .Y(n_821) );
INVx1_ASAP7_75t_L g1079 ( .A(n_434), .Y(n_1079) );
BUFx4f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g684 ( .A(n_435), .Y(n_684) );
INVx1_ASAP7_75t_L g787 ( .A(n_435), .Y(n_787) );
INVx1_ASAP7_75t_L g896 ( .A(n_435), .Y(n_896) );
BUFx2_ASAP7_75t_L g1029 ( .A(n_435), .Y(n_1029) );
INVx1_ASAP7_75t_L g1157 ( .A(n_435), .Y(n_1157) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
OR2x2_ASAP7_75t_L g479 ( .A(n_436), .B(n_438), .Y(n_479) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g883 ( .A(n_440), .Y(n_883) );
INVx1_ASAP7_75t_L g975 ( .A(n_440), .Y(n_975) );
INVx2_ASAP7_75t_L g1136 ( .A(n_440), .Y(n_1136) );
BUFx2_ASAP7_75t_L g1941 ( .A(n_440), .Y(n_1941) );
BUFx6f_ASAP7_75t_L g784 ( .A(n_441), .Y(n_784) );
INVx1_ASAP7_75t_L g1263 ( .A(n_441), .Y(n_1263) );
BUFx3_ASAP7_75t_L g1320 ( .A(n_441), .Y(n_1320) );
INVx1_ASAP7_75t_L g1331 ( .A(n_441), .Y(n_1331) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_442), .Y(n_470) );
INVx2_ASAP7_75t_L g483 ( .A(n_442), .Y(n_483) );
INVx1_ASAP7_75t_L g605 ( .A(n_442), .Y(n_605) );
INVx1_ASAP7_75t_L g768 ( .A(n_442), .Y(n_768) );
BUFx3_ASAP7_75t_L g468 ( .A(n_444), .Y(n_468) );
HB1xp67_ASAP7_75t_L g1020 ( .A(n_444), .Y(n_1020) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g601 ( .A(n_445), .Y(n_601) );
INVx1_ASAP7_75t_L g613 ( .A(n_445), .Y(n_613) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_445), .Y(n_675) );
INVx1_ASAP7_75t_L g686 ( .A(n_445), .Y(n_686) );
HB1xp67_ASAP7_75t_L g890 ( .A(n_445), .Y(n_890) );
INVx2_ASAP7_75t_SL g964 ( .A(n_445), .Y(n_964) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g701 ( .A(n_447), .Y(n_701) );
INVx2_ASAP7_75t_L g826 ( .A(n_447), .Y(n_826) );
INVx2_ASAP7_75t_SL g969 ( .A(n_447), .Y(n_969) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_454), .B1(n_455), .B2(n_467), .C(n_471), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g1015 ( .A1(n_450), .A2(n_471), .B1(n_1010), .B2(n_1016), .C(n_1019), .Y(n_1015) );
INVx1_ASAP7_75t_L g1939 ( .A(n_450), .Y(n_1939) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g830 ( .A(n_451), .Y(n_830) );
INVx1_ASAP7_75t_L g1084 ( .A(n_451), .Y(n_1084) );
INVx1_ASAP7_75t_L g1275 ( .A(n_451), .Y(n_1275) );
AOI221xp5_ASAP7_75t_L g1461 ( .A1(n_451), .A2(n_891), .B1(n_1453), .B2(n_1462), .C(n_1464), .Y(n_1461) );
AOI221xp5_ASAP7_75t_L g1568 ( .A1(n_451), .A2(n_471), .B1(n_1569), .B2(n_1571), .C(n_1573), .Y(n_1568) );
INVx2_ASAP7_75t_SL g599 ( .A(n_452), .Y(n_599) );
BUFx3_ASAP7_75t_L g608 ( .A(n_452), .Y(n_608) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_452), .Y(n_773) );
BUFx4f_ASAP7_75t_L g834 ( .A(n_452), .Y(n_834) );
AND2x4_ASAP7_75t_L g891 ( .A(n_452), .B(n_680), .Y(n_891) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_453), .Y(n_462) );
OAI22xp33_ASAP7_75t_L g562 ( .A1(n_454), .A2(n_476), .B1(n_563), .B2(n_566), .Y(n_562) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_458), .A2(n_474), .B1(n_591), .B2(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g668 ( .A(n_458), .Y(n_668) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_462), .Y(n_474) );
INVx2_ASAP7_75t_L g1090 ( .A(n_462), .Y(n_1090) );
BUFx6f_ASAP7_75t_L g1463 ( .A(n_462), .Y(n_1463) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g835 ( .A(n_465), .Y(n_835) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
BUFx3_ASAP7_75t_L g611 ( .A(n_466), .Y(n_611) );
INVx2_ASAP7_75t_L g692 ( .A(n_466), .Y(n_692) );
INVx1_ASAP7_75t_L g1318 ( .A(n_466), .Y(n_1318) );
INVx2_ASAP7_75t_SL g899 ( .A(n_469), .Y(n_899) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g670 ( .A(n_470), .Y(n_670) );
BUFx6f_ASAP7_75t_L g1022 ( .A(n_470), .Y(n_1022) );
INVx1_ASAP7_75t_L g1241 ( .A(n_470), .Y(n_1241) );
INVx1_ASAP7_75t_L g1644 ( .A(n_470), .Y(n_1644) );
AOI21xp33_ASAP7_75t_L g596 ( .A1(n_471), .A2(n_597), .B(n_602), .Y(n_596) );
INVx1_ASAP7_75t_L g774 ( .A(n_471), .Y(n_774) );
AOI221xp5_ASAP7_75t_L g828 ( .A1(n_471), .A2(n_829), .B1(n_831), .B2(n_832), .C(n_836), .Y(n_828) );
AOI221xp5_ASAP7_75t_L g1082 ( .A1(n_471), .A2(n_1083), .B1(n_1085), .B2(n_1086), .C(n_1091), .Y(n_1082) );
AOI221xp5_ASAP7_75t_L g1161 ( .A1(n_471), .A2(n_829), .B1(n_1162), .B2(n_1163), .C(n_1164), .Y(n_1161) );
AOI221xp5_ASAP7_75t_L g1232 ( .A1(n_471), .A2(n_829), .B1(n_1217), .B2(n_1233), .C(n_1234), .Y(n_1232) );
INVx1_ASAP7_75t_L g1280 ( .A(n_471), .Y(n_1280) );
HB1xp67_ASAP7_75t_L g1392 ( .A(n_471), .Y(n_1392) );
AOI221xp5_ASAP7_75t_L g1637 ( .A1(n_471), .A2(n_1083), .B1(n_1626), .B2(n_1638), .C(n_1641), .Y(n_1637) );
INVx1_ASAP7_75t_L g1945 ( .A(n_471), .Y(n_1945) );
AND2x4_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g777 ( .A(n_473), .B(n_778), .Y(n_777) );
BUFx6f_ASAP7_75t_L g887 ( .A(n_474), .Y(n_887) );
INVx1_ASAP7_75t_L g1018 ( .A(n_474), .Y(n_1018) );
INVx1_ASAP7_75t_L g1328 ( .A(n_474), .Y(n_1328) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B1(n_480), .B2(n_481), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_477), .A2(n_481), .B1(n_841), .B2(n_842), .Y(n_840) );
AOI22xp33_ASAP7_75t_SL g1031 ( .A1(n_477), .A2(n_481), .B1(n_1006), .B2(n_1008), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_477), .A2(n_481), .B1(n_1096), .B2(n_1097), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_477), .A2(n_481), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
AOI22xp33_ASAP7_75t_SL g1167 ( .A1(n_477), .A2(n_481), .B1(n_1168), .B2(n_1169), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g1393 ( .A1(n_477), .A2(n_481), .B1(n_1394), .B2(n_1395), .Y(n_1393) );
AOI22xp5_ASAP7_75t_L g1465 ( .A1(n_477), .A2(n_481), .B1(n_1446), .B2(n_1452), .Y(n_1465) );
AOI22xp33_ASAP7_75t_L g1574 ( .A1(n_477), .A2(n_481), .B1(n_1575), .B2(n_1576), .Y(n_1574) );
AOI22xp33_ASAP7_75t_L g1645 ( .A1(n_477), .A2(n_481), .B1(n_1622), .B2(n_1624), .Y(n_1645) );
AOI22xp33_ASAP7_75t_L g1946 ( .A1(n_477), .A2(n_481), .B1(n_1921), .B2(n_1923), .Y(n_1946) );
INVx6_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g586 ( .A(n_479), .Y(n_586) );
BUFx2_ASAP7_75t_L g823 ( .A(n_479), .Y(n_823) );
INVx1_ASAP7_75t_L g1081 ( .A(n_479), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_481), .B(n_1220), .Y(n_1249) );
INVx4_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g589 ( .A(n_483), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g879 ( .A1(n_484), .A2(n_880), .B(n_892), .Y(n_879) );
AOI31xp33_ASAP7_75t_L g1014 ( .A1(n_484), .A2(n_1015), .A3(n_1023), .B(n_1031), .Y(n_1014) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI31xp33_ASAP7_75t_L g958 ( .A1(n_485), .A2(n_959), .A3(n_960), .B(n_971), .Y(n_958) );
OAI31xp33_ASAP7_75t_SL g1309 ( .A1(n_485), .A2(n_1310), .A3(n_1319), .B(n_1324), .Y(n_1309) );
BUFx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g843 ( .A(n_486), .Y(n_843) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR2x6_ASAP7_75t_L g533 ( .A(n_487), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g620 ( .A(n_487), .Y(n_620) );
NOR3xp33_ASAP7_75t_SL g488 ( .A(n_489), .B(n_519), .C(n_532), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_506), .Y(n_489) );
BUFx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_493), .A2(n_822), .B1(n_851), .B2(n_852), .Y(n_850) );
BUFx2_ASAP7_75t_L g914 ( .A(n_493), .Y(n_914) );
BUFx2_ASAP7_75t_L g983 ( .A(n_493), .Y(n_983) );
BUFx2_ASAP7_75t_L g1051 ( .A(n_493), .Y(n_1051) );
BUFx2_ASAP7_75t_L g1106 ( .A(n_493), .Y(n_1106) );
BUFx2_ASAP7_75t_L g1197 ( .A(n_493), .Y(n_1197) );
BUFx2_ASAP7_75t_L g1304 ( .A(n_493), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_493), .A2(n_502), .B1(n_1322), .B2(n_1361), .Y(n_1360) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_498), .Y(n_493) );
BUFx3_ASAP7_75t_L g1180 ( .A(n_494), .Y(n_1180) );
INVx1_ASAP7_75t_L g1189 ( .A(n_494), .Y(n_1189) );
INVx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx3_ASAP7_75t_L g561 ( .A(n_495), .Y(n_561) );
BUFx6f_ASAP7_75t_L g943 ( .A(n_495), .Y(n_943) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_496), .Y(n_553) );
INVx1_ASAP7_75t_L g1450 ( .A(n_496), .Y(n_1450) );
AND2x4_ASAP7_75t_L g504 ( .A(n_497), .B(n_505), .Y(n_504) );
AND2x6_ASAP7_75t_L g502 ( .A(n_498), .B(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g508 ( .A(n_498), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g513 ( .A(n_498), .B(n_514), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_498), .A2(n_623), .B1(n_634), .B2(n_635), .Y(n_622) );
AND2x2_ASAP7_75t_L g704 ( .A(n_498), .B(n_514), .Y(n_704) );
AND2x2_ASAP7_75t_L g709 ( .A(n_498), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g712 ( .A(n_498), .B(n_561), .Y(n_712) );
AND2x2_ASAP7_75t_L g724 ( .A(n_498), .B(n_718), .Y(n_724) );
AND2x2_ASAP7_75t_L g849 ( .A(n_498), .B(n_514), .Y(n_849) );
AND2x2_ASAP7_75t_L g910 ( .A(n_498), .B(n_514), .Y(n_910) );
AND2x2_ASAP7_75t_L g1608 ( .A(n_498), .B(n_514), .Y(n_1608) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g571 ( .A(n_499), .Y(n_571) );
INVx2_ASAP7_75t_L g1525 ( .A(n_500), .Y(n_1525) );
AND2x4_ASAP7_75t_L g1538 ( .A(n_500), .B(n_629), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_500), .B(n_515), .Y(n_1554) );
INVx1_ASAP7_75t_L g535 ( .A(n_501), .Y(n_535) );
INVx1_ASAP7_75t_L g573 ( .A(n_501), .Y(n_573) );
INVx1_ASAP7_75t_SL g732 ( .A(n_502), .Y(n_732) );
BUFx2_ASAP7_75t_L g852 ( .A(n_502), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g908 ( .A1(n_502), .A2(n_909), .B1(n_910), .B2(n_911), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_502), .A2(n_704), .B1(n_953), .B2(n_954), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_502), .A2(n_982), .B1(n_983), .B2(n_984), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_502), .A2(n_1050), .B1(n_1051), .B2(n_1052), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_502), .A2(n_1105), .B1(n_1106), .B2(n_1107), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_502), .A2(n_1158), .B1(n_1196), .B2(n_1197), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_502), .A2(n_1106), .B1(n_1225), .B2(n_1226), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1580 ( .A1(n_502), .A2(n_1304), .B1(n_1581), .B2(n_1582), .Y(n_1580) );
AOI22xp33_ASAP7_75t_L g1602 ( .A1(n_502), .A2(n_1051), .B1(n_1603), .B2(n_1604), .Y(n_1602) );
NAND2x1p5_ASAP7_75t_L g531 ( .A(n_503), .B(n_526), .Y(n_531) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_503), .Y(n_1115) );
BUFx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_504), .Y(n_633) );
BUFx2_ASAP7_75t_L g661 ( .A(n_504), .Y(n_661) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_504), .Y(n_718) );
INVx1_ASAP7_75t_L g940 ( .A(n_504), .Y(n_940) );
BUFx3_ASAP7_75t_L g1526 ( .A(n_504), .Y(n_1526) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_512), .B2(n_513), .Y(n_506) );
BUFx2_ASAP7_75t_L g847 ( .A(n_508), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_508), .B(n_950), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_508), .A2(n_849), .B1(n_986), .B2(n_987), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_508), .A2(n_513), .B1(n_1054), .B2(n_1055), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_508), .A2(n_513), .B1(n_1109), .B2(n_1110), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_508), .A2(n_910), .B1(n_1159), .B2(n_1199), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_508), .A2(n_910), .B1(n_1228), .B2(n_1229), .Y(n_1227) );
AOI22xp33_ASAP7_75t_L g1294 ( .A1(n_508), .A2(n_513), .B1(n_1295), .B2(n_1296), .Y(n_1294) );
AOI22xp33_ASAP7_75t_L g1583 ( .A1(n_508), .A2(n_513), .B1(n_1584), .B2(n_1585), .Y(n_1583) );
AOI22xp33_ASAP7_75t_L g1605 ( .A1(n_508), .A2(n_1606), .B1(n_1607), .B2(n_1608), .Y(n_1605) );
INVx2_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_SL g710 ( .A(n_510), .Y(n_710) );
INVx2_ASAP7_75t_L g1288 ( .A(n_510), .Y(n_1288) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_511), .Y(n_629) );
AOI22xp33_ASAP7_75t_SL g1362 ( .A1(n_513), .A2(n_653), .B1(n_1326), .B2(n_1363), .Y(n_1362) );
INVx2_ASAP7_75t_SL g1300 ( .A(n_514), .Y(n_1300) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g637 ( .A(n_515), .Y(n_637) );
INVx1_ASAP7_75t_L g647 ( .A(n_515), .Y(n_647) );
BUFx6f_ASAP7_75t_L g716 ( .A(n_515), .Y(n_716) );
BUFx6f_ASAP7_75t_L g945 ( .A(n_515), .Y(n_945) );
BUFx2_ASAP7_75t_L g1117 ( .A(n_515), .Y(n_1117) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g529 ( .A(n_516), .Y(n_529) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_SL g989 ( .A(n_521), .Y(n_989) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2x1_ASAP7_75t_SL g522 ( .A(n_523), .B(n_526), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g1292 ( .A1(n_523), .A2(n_528), .B1(n_1278), .B2(n_1279), .Y(n_1292) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_525), .Y(n_656) );
NAND2x1p5_ASAP7_75t_L g527 ( .A(n_526), .B(n_528), .Y(n_527) );
AND2x4_ASAP7_75t_L g655 ( .A(n_526), .B(n_656), .Y(n_655) );
AND2x4_ASAP7_75t_L g657 ( .A(n_526), .B(n_658), .Y(n_657) );
AND2x4_ASAP7_75t_L g660 ( .A(n_526), .B(n_661), .Y(n_660) );
AOI32xp33_ASAP7_75t_L g1284 ( .A1(n_526), .A2(n_1058), .A3(n_1285), .B1(n_1287), .B2(n_1289), .Y(n_1284) );
BUFx4f_ASAP7_75t_L g737 ( .A(n_527), .Y(n_737) );
BUFx4f_ASAP7_75t_L g1222 ( .A(n_527), .Y(n_1222) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OR2x6_ASAP7_75t_L g1535 ( .A(n_529), .B(n_1518), .Y(n_1535) );
BUFx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx3_ASAP7_75t_L g738 ( .A(n_531), .Y(n_738) );
BUFx2_ASAP7_75t_L g855 ( .A(n_531), .Y(n_855) );
OAI33xp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_536), .A3(n_546), .B1(n_555), .B2(n_562), .B3(n_568), .Y(n_532) );
OAI33xp33_ASAP7_75t_L g856 ( .A1(n_533), .A2(n_857), .A3(n_862), .B1(n_868), .B2(n_871), .B3(n_872), .Y(n_856) );
OAI33xp33_ASAP7_75t_L g990 ( .A1(n_533), .A2(n_568), .A3(n_991), .B1(n_996), .B2(n_1001), .B3(n_1007), .Y(n_990) );
OAI33xp33_ASAP7_75t_L g1172 ( .A1(n_533), .A2(n_568), .A3(n_1173), .B1(n_1181), .B2(n_1187), .B3(n_1190), .Y(n_1172) );
OAI33xp33_ASAP7_75t_L g1204 ( .A1(n_533), .A2(n_568), .A3(n_1205), .B1(n_1209), .B2(n_1213), .B3(n_1218), .Y(n_1204) );
OAI33xp33_ASAP7_75t_L g1340 ( .A1(n_533), .A2(n_1341), .A3(n_1346), .B1(n_1350), .B2(n_1355), .B3(n_1358), .Y(n_1340) );
OAI33xp33_ASAP7_75t_L g1434 ( .A1(n_533), .A2(n_872), .A3(n_1435), .B1(n_1439), .B2(n_1443), .B3(n_1451), .Y(n_1434) );
OAI33xp33_ASAP7_75t_L g1587 ( .A1(n_533), .A2(n_568), .A3(n_1588), .B1(n_1591), .B2(n_1594), .B3(n_1595), .Y(n_1587) );
HB1xp67_ASAP7_75t_L g1611 ( .A(n_533), .Y(n_1611) );
OAI22xp33_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_539), .B1(n_540), .B2(n_545), .Y(n_536) );
OAI22xp33_ASAP7_75t_L g1301 ( .A1(n_537), .A2(n_1009), .B1(n_1272), .B2(n_1302), .Y(n_1301) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g746 ( .A(n_538), .Y(n_746) );
INVx1_ASAP7_75t_L g1914 ( .A(n_538), .Y(n_1914) );
OAI22xp33_ASAP7_75t_L g1213 ( .A1(n_540), .A2(n_1214), .B1(n_1216), .B2(n_1217), .Y(n_1213) );
OAI22xp33_ASAP7_75t_L g1595 ( .A1(n_540), .A2(n_1183), .B1(n_1573), .B2(n_1575), .Y(n_1595) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx3_ASAP7_75t_L g567 ( .A(n_542), .Y(n_567) );
INVx2_ASAP7_75t_L g1345 ( .A(n_542), .Y(n_1345) );
INVx2_ASAP7_75t_L g1438 ( .A(n_542), .Y(n_1438) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_543), .B(n_544), .Y(n_723) );
INVx1_ASAP7_75t_L g659 ( .A(n_544), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_550), .B1(n_551), .B2(n_554), .Y(n_546) );
BUFx2_ASAP7_75t_L g1207 ( .A(n_547), .Y(n_1207) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_548), .Y(n_864) );
INVx1_ASAP7_75t_L g1348 ( .A(n_548), .Y(n_1348) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g558 ( .A(n_549), .Y(n_558) );
BUFx2_ASAP7_75t_L g753 ( .A(n_549), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g1218 ( .A1(n_551), .A2(n_556), .B1(n_1219), .B2(n_1220), .Y(n_1218) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_SL g625 ( .A(n_553), .Y(n_625) );
INVx2_ASAP7_75t_SL g649 ( .A(n_553), .Y(n_649) );
INVx4_ASAP7_75t_L g743 ( .A(n_553), .Y(n_743) );
INVx2_ASAP7_75t_SL g866 ( .A(n_553), .Y(n_866) );
INVx2_ASAP7_75t_SL g1064 ( .A(n_553), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_556), .A2(n_741), .B1(n_742), .B2(n_743), .Y(n_740) );
INVx2_ASAP7_75t_L g1618 ( .A(n_556), .Y(n_1618) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g624 ( .A(n_557), .Y(n_624) );
INVx2_ASAP7_75t_SL g870 ( .A(n_557), .Y(n_870) );
INVx2_ASAP7_75t_L g1445 ( .A(n_557), .Y(n_1445) );
BUFx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g1177 ( .A(n_558), .Y(n_1177) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g919 ( .A(n_560), .Y(n_919) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g639 ( .A(n_561), .Y(n_639) );
INVx2_ASAP7_75t_L g754 ( .A(n_561), .Y(n_754) );
OAI22xp33_ASAP7_75t_L g1209 ( .A1(n_563), .A2(n_1210), .B1(n_1211), .B2(n_1212), .Y(n_1209) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OAI22xp33_ASAP7_75t_L g640 ( .A1(n_565), .A2(n_567), .B1(n_592), .B2(n_641), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_565), .A2(n_567), .B1(n_651), .B2(n_652), .Y(n_650) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_565), .A2(n_757), .B1(n_758), .B2(n_759), .Y(n_756) );
BUFx2_ASAP7_75t_L g1183 ( .A(n_565), .Y(n_1183) );
INVx1_ASAP7_75t_L g1215 ( .A(n_565), .Y(n_1215) );
OAI22xp33_ASAP7_75t_L g1623 ( .A1(n_565), .A2(n_1624), .B1(n_1625), .B2(n_1626), .Y(n_1623) );
OAI22xp33_ASAP7_75t_L g1190 ( .A1(n_566), .A2(n_1162), .B1(n_1168), .B2(n_1191), .Y(n_1190) );
BUFx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g1186 ( .A(n_567), .Y(n_1186) );
INVx1_ASAP7_75t_L g1415 ( .A(n_568), .Y(n_1415) );
CKINVDCx8_ASAP7_75t_R g568 ( .A(n_569), .Y(n_568) );
INVx5_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx6_ASAP7_75t_L g634 ( .A(n_570), .Y(n_634) );
OR2x6_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx2_ASAP7_75t_L g948 ( .A(n_572), .Y(n_948) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
OAI22x1_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_727), .B2(n_804), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
XNOR2x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_662), .Y(n_578) );
XNOR2x1_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g1689 ( .A1(n_580), .A2(n_1690), .B1(n_1692), .B2(n_1693), .Y(n_1689) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_621), .Y(n_581) );
AOI31xp33_ASAP7_75t_SL g582 ( .A1(n_583), .A2(n_596), .A3(n_606), .B(n_618), .Y(n_582) );
OAI221xp5_ASAP7_75t_L g1027 ( .A1(n_585), .A2(n_984), .B1(n_986), .B2(n_1028), .C(n_1030), .Y(n_1027) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g667 ( .A(n_586), .Y(n_667) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_586), .Y(n_782) );
INVx2_ASAP7_75t_L g797 ( .A(n_586), .Y(n_797) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g818 ( .A(n_589), .Y(n_818) );
INVx2_ASAP7_75t_SL g776 ( .A(n_593), .Y(n_776) );
INVx1_ASAP7_75t_L g1074 ( .A(n_593), .Y(n_1074) );
INVx1_ASAP7_75t_L g1152 ( .A(n_593), .Y(n_1152) );
AOI322xp5_ASAP7_75t_L g1237 ( .A1(n_593), .A2(n_1076), .A3(n_1238), .B1(n_1242), .B2(n_1244), .C1(n_1246), .C2(n_1247), .Y(n_1237) );
AOI222xp33_ASAP7_75t_L g1276 ( .A1(n_593), .A2(n_615), .B1(n_1076), .B2(n_1277), .C1(n_1278), .C2(n_1279), .Y(n_1276) );
INVx2_ASAP7_75t_SL g1567 ( .A(n_593), .Y(n_1567) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_594), .A2(n_595), .B1(n_655), .B2(n_657), .C(n_660), .Y(n_654) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g1243 ( .A(n_599), .Y(n_1243) );
INVx1_ASAP7_75t_L g1270 ( .A(n_599), .Y(n_1270) );
HB1xp67_ASAP7_75t_L g1391 ( .A(n_600), .Y(n_1391) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g1166 ( .A(n_601), .Y(n_1166) );
INVxp67_ASAP7_75t_L g793 ( .A(n_603), .Y(n_793) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g614 ( .A(n_605), .Y(n_614) );
INVx1_ASAP7_75t_L g839 ( .A(n_605), .Y(n_839) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_612), .B1(n_615), .B2(n_617), .Y(n_606) );
INVx3_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI221xp5_ASAP7_75t_L g785 ( .A1(n_611), .A2(n_741), .B1(n_747), .B2(n_786), .C(n_788), .Y(n_785) );
INVx1_ASAP7_75t_L g1267 ( .A(n_611), .Y(n_1267) );
BUFx2_ASAP7_75t_L g1504 ( .A(n_613), .Y(n_1504) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_617), .A2(n_643), .B1(n_645), .B2(n_653), .Y(n_642) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AOI211xp5_ASAP7_75t_L g663 ( .A1(n_619), .A2(n_664), .B(n_702), .C(n_713), .Y(n_663) );
NOR2xp67_ASAP7_75t_L g1515 ( .A(n_619), .B(n_1516), .Y(n_1515) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x4_ASAP7_75t_L g643 ( .A(n_620), .B(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g801 ( .A(n_620), .Y(n_801) );
AND2x2_ASAP7_75t_L g947 ( .A(n_620), .B(n_948), .Y(n_947) );
AND2x4_ASAP7_75t_L g1058 ( .A(n_620), .B(n_644), .Y(n_1058) );
OR2x6_ASAP7_75t_L g1500 ( .A(n_620), .B(n_692), .Y(n_1500) );
AOI31xp33_ASAP7_75t_L g1629 ( .A1(n_620), .A2(n_1630), .A3(n_1637), .B(n_1645), .Y(n_1629) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_642), .C(n_654), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_624), .A2(n_997), .B1(n_998), .B2(n_999), .Y(n_996) );
OAI221xp5_ASAP7_75t_L g1527 ( .A1(n_624), .A2(n_649), .B1(n_1474), .B2(n_1478), .C(n_1528), .Y(n_1527) );
OAI22xp5_ASAP7_75t_L g1912 ( .A1(n_625), .A2(n_1913), .B1(n_1914), .B2(n_1915), .Y(n_1912) );
OAI22xp5_ASAP7_75t_L g1919 ( .A1(n_625), .A2(n_1617), .B1(n_1920), .B2(n_1921), .Y(n_1919) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_630), .B2(n_631), .Y(n_626) );
HB1xp67_ASAP7_75t_L g1114 ( .A(n_628), .Y(n_1114) );
INVx1_ASAP7_75t_L g1121 ( .A(n_628), .Y(n_1121) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx3_ASAP7_75t_L g938 ( .A(n_629), .Y(n_938) );
BUFx2_ASAP7_75t_L g1060 ( .A(n_629), .Y(n_1060) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
AOI322xp5_ASAP7_75t_L g714 ( .A1(n_634), .A2(n_643), .A3(n_694), .B1(n_715), .B2(n_717), .C1(n_719), .C2(n_724), .Y(n_714) );
INVx1_ASAP7_75t_L g872 ( .A(n_634), .Y(n_872) );
AOI222xp33_ASAP7_75t_L g916 ( .A1(n_634), .A2(n_643), .B1(n_709), .B2(n_917), .C1(n_918), .C2(n_924), .Y(n_916) );
AOI33xp33_ASAP7_75t_L g1056 ( .A1(n_634), .A2(n_1057), .A3(n_1059), .B1(n_1061), .B2(n_1065), .B3(n_1066), .Y(n_1056) );
AOI33xp33_ASAP7_75t_L g1111 ( .A1(n_634), .A2(n_1112), .A3(n_1113), .B1(n_1116), .B2(n_1118), .B3(n_1119), .Y(n_1111) );
AOI22xp5_ASAP7_75t_L g1297 ( .A1(n_634), .A2(n_1298), .B1(n_1303), .B2(n_1304), .Y(n_1297) );
INVx2_ASAP7_75t_L g1358 ( .A(n_634), .Y(n_1358) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g1000 ( .A(n_639), .Y(n_1000) );
AOI33xp33_ASAP7_75t_L g935 ( .A1(n_643), .A2(n_936), .A3(n_941), .B1(n_944), .B2(n_946), .B3(n_947), .Y(n_935) );
BUFx2_ASAP7_75t_L g1112 ( .A(n_643), .Y(n_1112) );
INVx1_ASAP7_75t_L g1543 ( .A(n_644), .Y(n_1543) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g925 ( .A(n_647), .Y(n_925) );
INVxp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI22xp33_ASAP7_75t_L g1612 ( .A1(n_649), .A2(n_759), .B1(n_1613), .B2(n_1614), .Y(n_1612) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_653), .A2(n_657), .B1(n_673), .B2(n_706), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g912 ( .A1(n_653), .A2(n_913), .B1(n_914), .B2(n_915), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_653), .A2(n_712), .B1(n_956), .B2(n_957), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_655), .A2(n_660), .B(n_726), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g905 ( .A1(n_655), .A2(n_657), .B1(n_660), .B2(n_906), .C(n_907), .Y(n_905) );
AOI221xp5_ASAP7_75t_L g932 ( .A1(n_655), .A2(n_657), .B1(n_660), .B2(n_933), .C(n_934), .Y(n_932) );
AOI221xp5_ASAP7_75t_L g1043 ( .A1(n_655), .A2(n_1044), .B1(n_1046), .B2(n_1047), .C(n_1048), .Y(n_1043) );
AOI221xp5_ASAP7_75t_L g1101 ( .A1(n_655), .A2(n_657), .B1(n_660), .B2(n_1102), .C(n_1103), .Y(n_1101) );
INVx1_ASAP7_75t_L g1366 ( .A(n_655), .Y(n_1366) );
AOI221xp5_ASAP7_75t_L g1416 ( .A1(n_655), .A2(n_657), .B1(n_660), .B2(n_1417), .C(n_1418), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_656), .B(n_1517), .Y(n_1533) );
INVx1_ASAP7_75t_L g1045 ( .A(n_657), .Y(n_1045) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
HB1xp67_ASAP7_75t_L g1048 ( .A(n_660), .Y(n_1048) );
AOI221xp5_ASAP7_75t_L g1364 ( .A1(n_660), .A2(n_1044), .B1(n_1337), .B2(n_1338), .C(n_1365), .Y(n_1364) );
HB1xp67_ASAP7_75t_L g1412 ( .A(n_661), .Y(n_1412) );
NAND4xp25_ASAP7_75t_L g664 ( .A(n_665), .B(n_672), .C(n_681), .D(n_693), .Y(n_664) );
INVx1_ASAP7_75t_L g1026 ( .A(n_668), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_670), .A2(n_792), .B1(n_793), .B2(n_794), .Y(n_791) );
INVx1_ASAP7_75t_L g884 ( .A(n_670), .Y(n_884) );
INVx1_ASAP7_75t_L g1380 ( .A(n_670), .Y(n_1380) );
OAI221xp5_ASAP7_75t_L g1933 ( .A1(n_670), .A2(n_1640), .B1(n_1907), .B2(n_1934), .C(n_1935), .Y(n_1933) );
OAI221xp5_ASAP7_75t_L g1321 ( .A1(n_671), .A2(n_1030), .B1(n_1080), .B2(n_1322), .C(n_1323), .Y(n_1321) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B(n_676), .C(n_679), .Y(n_672) );
A2O1A1Ixp33_ASAP7_75t_SL g1325 ( .A1(n_674), .A2(n_679), .B(n_1326), .C(n_1327), .Y(n_1325) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx4_ASAP7_75t_L g765 ( .A(n_675), .Y(n_765) );
INVx2_ASAP7_75t_L g838 ( .A(n_675), .Y(n_838) );
BUFx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI211xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B(n_685), .C(n_687), .Y(n_681) );
OAI211xp5_ASAP7_75t_L g966 ( .A1(n_683), .A2(n_954), .B(n_967), .C(n_968), .Y(n_966) );
BUFx3_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g696 ( .A(n_684), .Y(n_696) );
OR2x6_ASAP7_75t_L g1486 ( .A(n_684), .B(n_1477), .Y(n_1486) );
INVx1_ASAP7_75t_L g1312 ( .A(n_686), .Y(n_1312) );
HB1xp67_ASAP7_75t_L g1642 ( .A(n_686), .Y(n_1642) );
INVx2_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g1239 ( .A(n_689), .Y(n_1239) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI211xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B(n_697), .C(n_699), .Y(n_693) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_SL g771 ( .A(n_698), .Y(n_771) );
BUFx3_ASAP7_75t_L g819 ( .A(n_698), .Y(n_819) );
INVx1_ASAP7_75t_L g799 ( .A(n_701), .Y(n_799) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g731 ( .A(n_704), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g1430 ( .A1(n_704), .A2(n_709), .B1(n_1431), .B2(n_1432), .Y(n_1430) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_709), .B1(n_711), .B2(n_712), .Y(n_707) );
INVx1_ASAP7_75t_L g761 ( .A(n_709), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g1516 ( .A(n_710), .B(n_1517), .Y(n_1516) );
INVx2_ASAP7_75t_L g734 ( .A(n_712), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g1427 ( .A1(n_712), .A2(n_724), .B1(n_1428), .B2(n_1429), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_725), .Y(n_713) );
BUFx6f_ASAP7_75t_L g1067 ( .A(n_718), .Y(n_1067) );
BUFx3_ASAP7_75t_L g748 ( .A(n_722), .Y(n_748) );
INVx2_ASAP7_75t_L g760 ( .A(n_722), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_722), .A2(n_921), .B1(n_922), .B2(n_923), .Y(n_920) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g804 ( .A(n_727), .Y(n_804) );
INVx1_ASAP7_75t_L g802 ( .A(n_728), .Y(n_802) );
NAND3xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_735), .C(n_762), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_733), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_739), .Y(n_735) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_737), .Y(n_854) );
HB1xp67_ASAP7_75t_L g1910 ( .A(n_737), .Y(n_1910) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_742), .A2(n_745), .B1(n_781), .B2(n_783), .Y(n_780) );
INVx2_ASAP7_75t_L g1286 ( .A(n_743), .Y(n_1286) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_744) );
OAI22xp33_ASAP7_75t_L g1341 ( .A1(n_746), .A2(n_1315), .B1(n_1342), .B2(n_1343), .Y(n_1341) );
OAI22xp33_ASAP7_75t_L g1355 ( .A1(n_746), .A2(n_1009), .B1(n_1356), .B2(n_1357), .Y(n_1355) );
BUFx3_ASAP7_75t_L g995 ( .A(n_748), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_751), .B1(n_754), .B2(n_755), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_750), .A2(n_758), .B1(n_770), .B2(n_772), .Y(n_769) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
BUFx2_ASAP7_75t_L g1002 ( .A(n_753), .Y(n_1002) );
INVx2_ASAP7_75t_L g926 ( .A(n_754), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_754), .A2(n_1206), .B1(n_1207), .B2(n_1208), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_755), .A2(n_757), .B1(n_765), .B2(n_766), .Y(n_764) );
OAI22xp33_ASAP7_75t_L g857 ( .A1(n_759), .A2(n_858), .B1(n_860), .B2(n_861), .Y(n_857) );
OAI22xp33_ASAP7_75t_L g871 ( .A1(n_759), .A2(n_831), .B1(n_842), .B2(n_866), .Y(n_871) );
OAI22xp5_ASAP7_75t_SL g1451 ( .A1(n_759), .A2(n_858), .B1(n_1452), .B2(n_1453), .Y(n_1451) );
OAI22xp5_ASAP7_75t_L g1916 ( .A1(n_759), .A2(n_1617), .B1(n_1917), .B2(n_1918), .Y(n_1916) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g1009 ( .A(n_760), .Y(n_1009) );
INVx1_ASAP7_75t_L g1212 ( .A(n_760), .Y(n_1212) );
OAI31xp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_775), .A3(n_779), .B(n_800), .Y(n_762) );
BUFx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OR2x6_ASAP7_75t_L g1480 ( .A(n_768), .B(n_1477), .Y(n_1480) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
BUFx2_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
HB1xp67_ASAP7_75t_L g1502 ( .A(n_773), .Y(n_1502) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_773), .B(n_1511), .Y(n_1510) );
OR2x6_ASAP7_75t_L g1497 ( .A(n_778), .B(n_1494), .Y(n_1497) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_785), .B1(n_791), .B2(n_795), .Y(n_779) );
OAI21xp5_ASAP7_75t_SL g1381 ( .A1(n_781), .A2(n_1382), .B(n_1383), .Y(n_1381) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
OAI221xp5_ASAP7_75t_L g795 ( .A1(n_786), .A2(n_796), .B1(n_797), .B2(n_798), .C(n_799), .Y(n_795) );
INVx1_ASAP7_75t_L g1384 ( .A(n_786), .Y(n_1384) );
BUFx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
BUFx3_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g1155 ( .A(n_790), .Y(n_1155) );
INVx2_ASAP7_75t_SL g1266 ( .A(n_790), .Y(n_1266) );
AOI22xp5_ASAP7_75t_L g1454 ( .A1(n_800), .A2(n_1455), .B1(n_1466), .B2(n_1467), .Y(n_1454) );
CKINVDCx8_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
AOI31xp33_ASAP7_75t_L g1070 ( .A1(n_801), .A2(n_1071), .A3(n_1082), .B(n_1095), .Y(n_1070) );
INVx1_ASAP7_75t_SL g1033 ( .A(n_805), .Y(n_1033) );
XNOR2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_874), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_844), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B(n_812), .Y(n_809) );
AOI31xp33_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_828), .A3(n_840), .B(n_843), .Y(n_812) );
AOI211xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B(n_816), .C(n_827), .Y(n_813) );
OAI22xp33_ASAP7_75t_L g868 ( .A1(n_814), .A2(n_841), .B1(n_858), .B2(n_869), .Y(n_868) );
AOI21xp5_ASAP7_75t_L g1931 ( .A1(n_815), .A2(n_1920), .B(n_1932), .Y(n_1931) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_822), .B1(n_823), .B2(n_824), .C(n_825), .Y(n_820) );
OAI211xp5_ASAP7_75t_L g961 ( .A1(n_821), .A2(n_962), .B(n_963), .C(n_965), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_824), .A2(n_847), .B1(n_848), .B2(n_849), .Y(n_846) );
OAI221xp5_ASAP7_75t_L g1078 ( .A1(n_825), .A2(n_1052), .B1(n_1054), .B2(n_1079), .C(n_1080), .Y(n_1078) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
BUFx2_ASAP7_75t_L g1245 ( .A(n_826), .Y(n_1245) );
AOI221xp5_ASAP7_75t_L g1132 ( .A1(n_829), .A2(n_891), .B1(n_1133), .B2(n_1134), .C(n_1137), .Y(n_1132) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
BUFx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g1123 ( .A(n_843), .Y(n_1123) );
BUFx8_ASAP7_75t_SL g1170 ( .A(n_843), .Y(n_1170) );
NOR3xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_853), .C(n_856), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_850), .Y(n_845) );
AOI21xp5_ASAP7_75t_L g1339 ( .A1(n_847), .A2(n_1323), .B(n_1340), .Y(n_1339) );
INVx1_ASAP7_75t_L g1399 ( .A(n_847), .Y(n_1399) );
AOI22xp33_ASAP7_75t_L g1905 ( .A1(n_847), .A2(n_1906), .B1(n_1907), .B2(n_1908), .Y(n_1905) );
INVx1_ASAP7_75t_L g1400 ( .A(n_849), .Y(n_1400) );
AOI22xp33_ASAP7_75t_L g1401 ( .A1(n_852), .A2(n_914), .B1(n_1402), .B2(n_1403), .Y(n_1401) );
INVxp67_ASAP7_75t_SL g1904 ( .A(n_852), .Y(n_1904) );
BUFx2_ASAP7_75t_L g993 ( .A(n_858), .Y(n_993) );
OAI221xp5_ASAP7_75t_L g1539 ( .A1(n_858), .A2(n_995), .B1(n_1540), .B2(n_1541), .C(n_1542), .Y(n_1539) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g1544 ( .A1(n_863), .A2(n_1545), .B1(n_1546), .B2(n_1550), .Y(n_1544) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
OAI22xp5_ASAP7_75t_SL g1591 ( .A1(n_866), .A2(n_1188), .B1(n_1592), .B2(n_1593), .Y(n_1591) );
OAI22xp5_ASAP7_75t_L g1620 ( .A1(n_866), .A2(n_869), .B1(n_1621), .B2(n_1622), .Y(n_1620) );
BUFx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_870), .A2(n_1351), .B1(n_1352), .B2(n_1354), .Y(n_1350) );
OAI33xp33_ASAP7_75t_L g1610 ( .A1(n_872), .A2(n_1611), .A3(n_1612), .B1(n_1615), .B2(n_1620), .B3(n_1623), .Y(n_1610) );
OAI22xp5_ASAP7_75t_L g1722 ( .A1(n_873), .A2(n_1693), .B1(n_1723), .B2(n_1724), .Y(n_1722) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_875), .A2(n_876), .B1(n_977), .B2(n_1032), .Y(n_874) );
INVx1_ASAP7_75t_SL g875 ( .A(n_876), .Y(n_875) );
XNOR2x1_ASAP7_75t_L g876 ( .A(n_877), .B(n_929), .Y(n_876) );
NOR2x1_ASAP7_75t_L g878 ( .A(n_879), .B(n_904), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_882), .B1(n_885), .B2(n_888), .C(n_891), .Y(n_880) );
HB1xp67_ASAP7_75t_L g1389 ( .A(n_887), .Y(n_1389) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g970 ( .A(n_891), .Y(n_970) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx2_ASAP7_75t_SL g1128 ( .A(n_903), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1334 ( .A1(n_903), .A2(n_1335), .B1(n_1337), .B2(n_1338), .Y(n_1334) );
NAND4xp25_ASAP7_75t_L g904 ( .A(n_905), .B(n_908), .C(n_912), .D(n_916), .Y(n_904) );
INVx2_ASAP7_75t_SL g1291 ( .A(n_922), .Y(n_1291) );
INVx1_ASAP7_75t_L g1442 ( .A(n_926), .Y(n_1442) );
NAND3xp33_ASAP7_75t_L g930 ( .A(n_931), .B(n_951), .C(n_958), .Y(n_930) );
AND3x1_ASAP7_75t_L g931 ( .A(n_932), .B(n_935), .C(n_949), .Y(n_931) );
INVx2_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx2_ASAP7_75t_SL g1529 ( .A(n_938), .Y(n_1529) );
INVx2_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx2_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx2_ASAP7_75t_L g1005 ( .A(n_943), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_943), .A2(n_1316), .B1(n_1347), .B2(n_1349), .Y(n_1346) );
INVx3_ASAP7_75t_L g1353 ( .A(n_943), .Y(n_1353) );
BUFx3_ASAP7_75t_L g1062 ( .A(n_945), .Y(n_1062) );
INVx2_ASAP7_75t_SL g1530 ( .A(n_948), .Y(n_1530) );
AND2x2_ASAP7_75t_L g951 ( .A(n_952), .B(n_955), .Y(n_951) );
NAND3xp33_ASAP7_75t_L g960 ( .A(n_961), .B(n_966), .C(n_970), .Y(n_960) );
INVx1_ASAP7_75t_L g1236 ( .A(n_964), .Y(n_1236) );
INVx1_ASAP7_75t_L g1030 ( .A(n_969), .Y(n_1030) );
INVx1_ASAP7_75t_L g1160 ( .A(n_969), .Y(n_1160) );
INVx2_ASAP7_75t_L g1032 ( .A(n_977), .Y(n_1032) );
AND2x2_ASAP7_75t_L g978 ( .A(n_979), .B(n_1011), .Y(n_978) );
NOR3xp33_ASAP7_75t_SL g979 ( .A(n_980), .B(n_988), .C(n_990), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_981), .B(n_985), .Y(n_980) );
OAI22xp33_ASAP7_75t_L g991 ( .A1(n_992), .A2(n_993), .B1(n_994), .B2(n_995), .Y(n_991) );
OAI22xp33_ASAP7_75t_L g1007 ( .A1(n_993), .A2(n_1008), .B1(n_1009), .B2(n_1010), .Y(n_1007) );
OAI22xp33_ASAP7_75t_L g1922 ( .A1(n_995), .A2(n_1914), .B1(n_1923), .B2(n_1924), .Y(n_1922) );
INVx2_ASAP7_75t_SL g999 ( .A(n_1000), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_1002), .A2(n_1003), .B1(n_1004), .B2(n_1006), .Y(n_1001) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
AOI21xp5_ASAP7_75t_L g1011 ( .A1(n_1012), .A2(n_1013), .B(n_1014), .Y(n_1011) );
AOI21xp33_ASAP7_75t_L g1068 ( .A1(n_1012), .A2(n_1069), .B(n_1070), .Y(n_1068) );
AOI21xp5_ASAP7_75t_L g1627 ( .A1(n_1012), .A2(n_1628), .B(n_1629), .Y(n_1627) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1029), .Y(n_1314) );
INVx2_ASAP7_75t_SL g1333 ( .A(n_1029), .Y(n_1333) );
INVx1_ASAP7_75t_L g1936 ( .A(n_1030), .Y(n_1936) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1034), .Y(n_1650) );
XNOR2xp5_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1421), .Y(n_1034) );
AOI22xp5_ASAP7_75t_L g1035 ( .A1(n_1036), .A2(n_1037), .B1(n_1252), .B2(n_1420), .Y(n_1035) );
INVx2_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
AO22x2_ASAP7_75t_L g1037 ( .A1(n_1038), .A2(n_1039), .B1(n_1142), .B2(n_1143), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
XNOR2xp5_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1098), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1068), .Y(n_1041) );
AND4x1_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1049), .C(n_1053), .D(n_1056), .Y(n_1042) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
HB1xp67_ASAP7_75t_L g1908 ( .A(n_1051), .Y(n_1908) );
BUFx3_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx2_ASAP7_75t_L g1407 ( .A(n_1058), .Y(n_1407) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx2_ASAP7_75t_SL g1075 ( .A(n_1076), .Y(n_1075) );
OAI221xp5_ASAP7_75t_L g1156 ( .A1(n_1080), .A2(n_1157), .B1(n_1158), .B2(n_1159), .C(n_1160), .Y(n_1156) );
INVx2_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1942 ( .A(n_1088), .Y(n_1942) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1093), .B(n_1476), .Y(n_1483) );
INVx2_ASAP7_75t_SL g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1094), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1122), .Y(n_1099) );
AND4x1_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1104), .C(n_1108), .D(n_1111), .Y(n_1100) );
HB1xp67_ASAP7_75t_L g1411 ( .A(n_1117), .Y(n_1411) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
NAND3xp33_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1132), .C(n_1138), .Y(n_1124) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
XOR2xp5_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1200), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1171), .Y(n_1145) );
AOI31xp33_ASAP7_75t_L g1148 ( .A1(n_1149), .A2(n_1161), .A3(n_1167), .B(n_1170), .Y(n_1148) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_1150), .A2(n_1169), .B1(n_1188), .B2(n_1189), .Y(n_1187) );
INVx2_ASAP7_75t_SL g1154 ( .A(n_1155), .Y(n_1154) );
INVx2_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
INVx5_ASAP7_75t_L g1281 ( .A(n_1170), .Y(n_1281) );
OAI31xp33_ASAP7_75t_L g1520 ( .A1(n_1170), .A2(n_1521), .A3(n_1536), .B(n_1552), .Y(n_1520) );
AOI31xp33_ASAP7_75t_L g1930 ( .A1(n_1170), .A2(n_1931), .A3(n_1937), .B(n_1946), .Y(n_1930) );
NOR3xp33_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1193), .C(n_1194), .Y(n_1171) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_1174), .A2(n_1175), .B1(n_1178), .B2(n_1179), .Y(n_1173) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
INVx2_ASAP7_75t_L g1188 ( .A(n_1176), .Y(n_1188) );
INVx2_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
OAI22xp5_ASAP7_75t_L g1594 ( .A1(n_1179), .A2(n_1188), .B1(n_1565), .B2(n_1576), .Y(n_1594) );
CKINVDCx5p33_ASAP7_75t_R g1179 ( .A(n_1180), .Y(n_1179) );
OAI22xp33_ASAP7_75t_L g1181 ( .A1(n_1182), .A2(n_1183), .B1(n_1184), .B2(n_1185), .Y(n_1181) );
OAI22xp33_ASAP7_75t_L g1588 ( .A1(n_1183), .A2(n_1438), .B1(n_1589), .B2(n_1590), .Y(n_1588) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
OAI22xp33_ASAP7_75t_SL g1615 ( .A1(n_1191), .A2(n_1616), .B1(n_1617), .B2(n_1619), .Y(n_1615) );
INVx3_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1198), .Y(n_1194) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1230), .Y(n_1202) );
NOR3xp33_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1221), .C(n_1223), .Y(n_1203) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1227), .Y(n_1223) );
NAND4xp25_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1237), .C(n_1248), .D(n_1249), .Y(n_1231) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1239), .B(n_1476), .Y(n_1475) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1252), .Y(n_1420) );
BUFx3_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
AOI22xp5_ASAP7_75t_L g1253 ( .A1(n_1254), .A2(n_1255), .B1(n_1367), .B2(n_1419), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
XNOR2xp5_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1307), .Y(n_1255) );
INVx2_ASAP7_75t_SL g1306 ( .A(n_1257), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1282), .Y(n_1257) );
OAI21xp33_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1274), .B(n_1281), .Y(n_1258) );
AOI22xp5_ASAP7_75t_L g1260 ( .A1(n_1261), .A2(n_1264), .B1(n_1268), .B2(n_1269), .Y(n_1260) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
OAI221xp5_ASAP7_75t_L g1313 ( .A1(n_1266), .A2(n_1314), .B1(n_1315), .B2(n_1316), .C(n_1317), .Y(n_1313) );
CKINVDCx5p33_ASAP7_75t_R g1386 ( .A(n_1275), .Y(n_1386) );
INVx1_ASAP7_75t_SL g1396 ( .A(n_1281), .Y(n_1396) );
NOR2xp33_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1293), .Y(n_1282) );
BUFx3_ASAP7_75t_L g1409 ( .A(n_1288), .Y(n_1409) );
OAI22xp33_ASAP7_75t_L g1435 ( .A1(n_1290), .A2(n_1436), .B1(n_1437), .B2(n_1438), .Y(n_1435) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1297), .Y(n_1293) );
INVx3_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
NAND4xp25_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1339), .C(n_1359), .D(n_1364), .Y(n_1308) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
NAND3xp33_ASAP7_75t_SL g1324 ( .A(n_1325), .B(n_1329), .C(n_1334), .Y(n_1324) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1328), .Y(n_1570) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
OR2x2_ASAP7_75t_L g1551 ( .A(n_1345), .B(n_1518), .Y(n_1551) );
HB1xp67_ASAP7_75t_L g1625 ( .A(n_1345), .Y(n_1625) );
OAI22xp5_ASAP7_75t_L g1439 ( .A1(n_1347), .A2(n_1440), .B1(n_1441), .B2(n_1442), .Y(n_1439) );
BUFx2_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1360), .B(n_1362), .Y(n_1359) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx2_ASAP7_75t_SL g1419 ( .A(n_1367), .Y(n_1419) );
XNOR2x1_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1369), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1397), .Y(n_1369) );
AOI21xp5_ASAP7_75t_L g1370 ( .A1(n_1371), .A2(n_1372), .B(n_1373), .Y(n_1370) );
AOI31xp33_ASAP7_75t_L g1373 ( .A1(n_1374), .A2(n_1385), .A3(n_1393), .B(n_1396), .Y(n_1373) );
AOI211xp5_ASAP7_75t_SL g1374 ( .A1(n_1375), .A2(n_1376), .B(n_1378), .C(n_1379), .Y(n_1374) );
AOI21xp5_ASAP7_75t_L g1630 ( .A1(n_1376), .A2(n_1621), .B(n_1631), .Y(n_1630) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
AOI221xp5_ASAP7_75t_L g1385 ( .A1(n_1386), .A2(n_1387), .B1(n_1388), .B2(n_1390), .C(n_1392), .Y(n_1385) );
NOR2xp33_ASAP7_75t_L g1397 ( .A(n_1398), .B(n_1404), .Y(n_1397) );
NAND2xp5_ASAP7_75t_SL g1404 ( .A(n_1405), .B(n_1416), .Y(n_1404) );
AOI33xp33_ASAP7_75t_L g1405 ( .A1(n_1406), .A2(n_1408), .A3(n_1410), .B1(n_1413), .B2(n_1414), .B3(n_1415), .Y(n_1405) );
INVx2_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1925 ( .A(n_1415), .Y(n_1925) );
OAI22xp33_ASAP7_75t_L g1421 ( .A1(n_1422), .A2(n_1468), .B1(n_1648), .B2(n_1649), .Y(n_1421) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1422), .Y(n_1648) );
XNOR2x1_ASAP7_75t_L g1422 ( .A(n_1423), .B(n_1424), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1454), .Y(n_1424) );
NOR3xp33_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1433), .C(n_1434), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_1427), .B(n_1430), .Y(n_1426) );
OAI22xp5_ASAP7_75t_SL g1443 ( .A1(n_1444), .A2(n_1445), .B1(n_1446), .B2(n_1447), .Y(n_1443) );
AOI221xp5_ASAP7_75t_L g1456 ( .A1(n_1444), .A2(n_1457), .B1(n_1458), .B2(n_1459), .C(n_1460), .Y(n_1456) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
HB1xp67_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
INVx2_ASAP7_75t_L g1549 ( .A(n_1450), .Y(n_1549) );
NAND3xp33_ASAP7_75t_L g1455 ( .A(n_1456), .B(n_1461), .C(n_1465), .Y(n_1455) );
INVx2_ASAP7_75t_L g1649 ( .A(n_1468), .Y(n_1649) );
XNOR2x1_ASAP7_75t_L g1468 ( .A(n_1469), .B(n_1557), .Y(n_1468) );
NAND3xp33_ASAP7_75t_L g1470 ( .A(n_1471), .B(n_1512), .C(n_1520), .Y(n_1470) );
NOR2xp33_ASAP7_75t_L g1471 ( .A(n_1472), .B(n_1487), .Y(n_1471) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1473), .B(n_1481), .Y(n_1472) );
AOI22xp33_ASAP7_75t_L g1473 ( .A1(n_1474), .A2(n_1475), .B1(n_1478), .B2(n_1479), .Y(n_1473) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
CKINVDCx6p67_ASAP7_75t_R g1479 ( .A(n_1480), .Y(n_1479) );
AOI22xp33_ASAP7_75t_L g1481 ( .A1(n_1482), .A2(n_1483), .B1(n_1484), .B2(n_1485), .Y(n_1481) );
CKINVDCx6p67_ASAP7_75t_R g1485 ( .A(n_1486), .Y(n_1485) );
NAND3xp33_ASAP7_75t_SL g1487 ( .A(n_1488), .B(n_1498), .C(n_1508), .Y(n_1487) );
AOI22xp33_ASAP7_75t_L g1488 ( .A1(n_1489), .A2(n_1490), .B1(n_1495), .B2(n_1496), .Y(n_1488) );
AOI22xp33_ASAP7_75t_L g1531 ( .A1(n_1489), .A2(n_1495), .B1(n_1532), .B2(n_1534), .Y(n_1531) );
INVx2_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
NAND2x1p5_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1493), .Y(n_1491) );
INVx2_ASAP7_75t_SL g1493 ( .A(n_1494), .Y(n_1493) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1494), .Y(n_1511) );
INVx2_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
AOI33xp33_ASAP7_75t_L g1498 ( .A1(n_1499), .A2(n_1501), .A3(n_1503), .B1(n_1505), .B2(n_1506), .B3(n_1507), .Y(n_1498) );
CKINVDCx5p33_ASAP7_75t_R g1499 ( .A(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1510), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1512 ( .A(n_1513), .B(n_1514), .Y(n_1512) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1518), .Y(n_1517) );
INVx2_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
INVx8_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
AND2x4_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1526), .Y(n_1523) );
AND2x4_ASAP7_75t_L g1556 ( .A(n_1524), .B(n_1549), .Y(n_1556) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
HB1xp67_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
CKINVDCx11_ASAP7_75t_R g1534 ( .A(n_1535), .Y(n_1534) );
CKINVDCx6p67_ASAP7_75t_R g1537 ( .A(n_1538), .Y(n_1537) );
INVx2_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
INVx3_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
INVx3_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
AO22x2_ASAP7_75t_L g1557 ( .A1(n_1558), .A2(n_1597), .B1(n_1646), .B2(n_1647), .Y(n_1557) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1558), .Y(n_1647) );
XOR2x2_ASAP7_75t_L g1558 ( .A(n_1559), .B(n_1596), .Y(n_1558) );
NAND2xp5_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1578), .Y(n_1559) );
NAND3xp33_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1568), .C(n_1574), .Y(n_1561) );
NOR3xp33_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1586), .C(n_1587), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1583), .Y(n_1579) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1597), .Y(n_1646) );
XNOR2xp5_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1599), .Y(n_1597) );
NAND2xp5_ASAP7_75t_L g1599 ( .A(n_1600), .B(n_1627), .Y(n_1599) );
NOR3xp33_ASAP7_75t_SL g1600 ( .A(n_1601), .B(n_1609), .C(n_1610), .Y(n_1600) );
NAND2xp5_ASAP7_75t_L g1601 ( .A(n_1602), .B(n_1605), .Y(n_1601) );
OAI33xp33_ASAP7_75t_L g1911 ( .A1(n_1611), .A2(n_1912), .A3(n_1916), .B1(n_1919), .B2(n_1922), .B3(n_1925), .Y(n_1911) );
INVx2_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
AOI31xp33_ASAP7_75t_L g1632 ( .A1(n_1633), .A2(n_1634), .A3(n_1635), .B(n_1636), .Y(n_1632) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
OAI221xp5_ASAP7_75t_L g1653 ( .A1(n_1654), .A2(n_1896), .B1(n_1898), .B2(n_1947), .C(n_1951), .Y(n_1653) );
AND4x1_ASAP7_75t_L g1654 ( .A(n_1655), .B(n_1823), .C(n_1837), .D(n_1869), .Y(n_1654) );
AOI211xp5_ASAP7_75t_L g1655 ( .A1(n_1656), .A2(n_1684), .B(n_1785), .C(n_1799), .Y(n_1655) );
NAND2xp5_ASAP7_75t_L g1800 ( .A(n_1656), .B(n_1801), .Y(n_1800) );
NAND2xp5_ASAP7_75t_L g1846 ( .A(n_1656), .B(n_1758), .Y(n_1846) );
AOI221xp5_ASAP7_75t_L g1864 ( .A1(n_1656), .A2(n_1734), .B1(n_1762), .B2(n_1865), .C(n_1866), .Y(n_1864) );
OAI333xp33_ASAP7_75t_L g1888 ( .A1(n_1656), .A2(n_1732), .A3(n_1790), .B1(n_1825), .B2(n_1889), .B3(n_1891), .C1(n_1892), .C2(n_1894), .C3(n_1895), .Y(n_1888) );
CKINVDCx5p33_ASAP7_75t_R g1656 ( .A(n_1657), .Y(n_1656) );
NAND2xp5_ASAP7_75t_L g1825 ( .A(n_1657), .B(n_1792), .Y(n_1825) );
OAI32xp33_ASAP7_75t_L g1845 ( .A1(n_1657), .A2(n_1697), .A3(n_1758), .B1(n_1817), .B2(n_1846), .Y(n_1845) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1657), .Y(n_1879) );
NAND2xp5_ASAP7_75t_L g1894 ( .A(n_1657), .B(n_1717), .Y(n_1894) );
OR2x6_ASAP7_75t_SL g1657 ( .A(n_1658), .B(n_1670), .Y(n_1657) );
OAI22xp5_ASAP7_75t_L g1658 ( .A1(n_1659), .A2(n_1660), .B1(n_1667), .B2(n_1668), .Y(n_1658) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1661), .Y(n_1660) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1661), .Y(n_1724) );
AND2x4_ASAP7_75t_L g1661 ( .A(n_1662), .B(n_1665), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1662), .B(n_1665), .Y(n_1691) );
HB1xp67_ASAP7_75t_L g1961 ( .A(n_1662), .Y(n_1961) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
AND2x4_ASAP7_75t_L g1669 ( .A(n_1663), .B(n_1665), .Y(n_1669) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
NAND2xp5_ASAP7_75t_L g1676 ( .A(n_1664), .B(n_1677), .Y(n_1676) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1666), .Y(n_1677) );
INVx2_ASAP7_75t_L g1707 ( .A(n_1668), .Y(n_1707) );
INVx1_ASAP7_75t_L g1897 ( .A(n_1668), .Y(n_1897) );
INVx2_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
INVx1_ASAP7_75t_SL g1693 ( .A(n_1669), .Y(n_1693) );
OAI22xp5_ASAP7_75t_L g1670 ( .A1(n_1671), .A2(n_1672), .B1(n_1678), .B2(n_1679), .Y(n_1670) );
BUFx3_ASAP7_75t_L g1672 ( .A(n_1673), .Y(n_1672) );
OAI22xp5_ASAP7_75t_L g1694 ( .A1(n_1673), .A2(n_1682), .B1(n_1695), .B2(n_1696), .Y(n_1694) );
OAI22xp33_ASAP7_75t_L g1719 ( .A1(n_1673), .A2(n_1680), .B1(n_1720), .B2(n_1721), .Y(n_1719) );
OAI22xp33_ASAP7_75t_L g1736 ( .A1(n_1673), .A2(n_1682), .B1(n_1737), .B2(n_1738), .Y(n_1736) );
BUFx6f_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
OAI22xp5_ASAP7_75t_L g1713 ( .A1(n_1674), .A2(n_1682), .B1(n_1714), .B2(n_1715), .Y(n_1713) );
OR2x2_ASAP7_75t_L g1674 ( .A(n_1675), .B(n_1676), .Y(n_1674) );
OR2x2_ASAP7_75t_L g1682 ( .A(n_1675), .B(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1675), .Y(n_1703) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1676), .Y(n_1702) );
HB1xp67_ASAP7_75t_L g1963 ( .A(n_1677), .Y(n_1963) );
HB1xp67_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1683), .Y(n_1705) );
NAND5xp2_ASAP7_75t_L g1684 ( .A(n_1685), .B(n_1753), .C(n_1766), .D(n_1774), .E(n_1778), .Y(n_1684) );
AOI211xp5_ASAP7_75t_SL g1685 ( .A1(n_1686), .A2(n_1716), .B(n_1728), .C(n_1749), .Y(n_1685) );
INVx1_ASAP7_75t_L g1835 ( .A(n_1686), .Y(n_1835) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_1687), .B(n_1697), .Y(n_1686) );
AND2x2_ASAP7_75t_L g1730 ( .A(n_1687), .B(n_1731), .Y(n_1730) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1687), .B(n_1732), .Y(n_1748) );
AND2x2_ASAP7_75t_L g1765 ( .A(n_1687), .B(n_1699), .Y(n_1765) );
NOR2xp33_ASAP7_75t_L g1777 ( .A(n_1687), .B(n_1699), .Y(n_1777) );
NAND2xp5_ASAP7_75t_L g1808 ( .A(n_1687), .B(n_1809), .Y(n_1808) );
AND2x2_ASAP7_75t_L g1820 ( .A(n_1687), .B(n_1743), .Y(n_1820) );
OR2x2_ASAP7_75t_L g1822 ( .A(n_1687), .B(n_1743), .Y(n_1822) );
AND2x2_ASAP7_75t_L g1844 ( .A(n_1687), .B(n_1742), .Y(n_1844) );
AND2x2_ASAP7_75t_L g1849 ( .A(n_1687), .B(n_1708), .Y(n_1849) );
NOR2xp33_ASAP7_75t_L g1860 ( .A(n_1687), .B(n_1760), .Y(n_1860) );
NOR2xp33_ASAP7_75t_L g1890 ( .A(n_1687), .B(n_1712), .Y(n_1890) );
CKINVDCx6p67_ASAP7_75t_R g1687 ( .A(n_1688), .Y(n_1687) );
OR2x2_ASAP7_75t_L g1780 ( .A(n_1688), .B(n_1732), .Y(n_1780) );
AND2x2_ASAP7_75t_L g1803 ( .A(n_1688), .B(n_1767), .Y(n_1803) );
AND2x2_ASAP7_75t_L g1815 ( .A(n_1688), .B(n_1732), .Y(n_1815) );
AND2x2_ASAP7_75t_L g1817 ( .A(n_1688), .B(n_1708), .Y(n_1817) );
NAND2xp5_ASAP7_75t_L g1829 ( .A(n_1688), .B(n_1830), .Y(n_1829) );
AND2x2_ASAP7_75t_L g1833 ( .A(n_1688), .B(n_1731), .Y(n_1833) );
AND2x2_ASAP7_75t_L g1863 ( .A(n_1688), .B(n_1742), .Y(n_1863) );
OR2x2_ASAP7_75t_L g1872 ( .A(n_1688), .B(n_1768), .Y(n_1872) );
OR2x6_ASAP7_75t_SL g1688 ( .A(n_1689), .B(n_1694), .Y(n_1688) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
AND2x2_ASAP7_75t_L g1697 ( .A(n_1698), .B(n_1708), .Y(n_1697) );
NAND2xp5_ASAP7_75t_L g1729 ( .A(n_1698), .B(n_1730), .Y(n_1729) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1698), .Y(n_1741) );
NOR2xp33_ASAP7_75t_L g1793 ( .A(n_1698), .B(n_1794), .Y(n_1793) );
NOR2xp33_ASAP7_75t_L g1830 ( .A(n_1698), .B(n_1768), .Y(n_1830) );
INVx4_ASAP7_75t_L g1698 ( .A(n_1699), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1747 ( .A(n_1699), .B(n_1748), .Y(n_1747) );
NAND2xp5_ASAP7_75t_L g1760 ( .A(n_1699), .B(n_1708), .Y(n_1760) );
INVx2_ASAP7_75t_L g1772 ( .A(n_1699), .Y(n_1772) );
AND2x2_ASAP7_75t_L g1809 ( .A(n_1699), .B(n_1718), .Y(n_1809) );
OR2x2_ASAP7_75t_L g1856 ( .A(n_1699), .B(n_1783), .Y(n_1856) );
NAND2xp5_ASAP7_75t_L g1862 ( .A(n_1699), .B(n_1863), .Y(n_1862) );
OR2x2_ASAP7_75t_L g1867 ( .A(n_1699), .B(n_1768), .Y(n_1867) );
OR2x2_ASAP7_75t_L g1871 ( .A(n_1699), .B(n_1872), .Y(n_1871) );
NAND2xp5_ASAP7_75t_L g1891 ( .A(n_1699), .B(n_1784), .Y(n_1891) );
AND2x2_ASAP7_75t_L g1893 ( .A(n_1699), .B(n_1762), .Y(n_1893) );
AND2x6_ASAP7_75t_L g1699 ( .A(n_1700), .B(n_1706), .Y(n_1699) );
AND2x4_ASAP7_75t_L g1701 ( .A(n_1702), .B(n_1703), .Y(n_1701) );
AND2x4_ASAP7_75t_L g1704 ( .A(n_1703), .B(n_1705), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1708 ( .A(n_1709), .B(n_1712), .Y(n_1708) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1709), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1742 ( .A(n_1709), .B(n_1743), .Y(n_1742) );
OR2x2_ASAP7_75t_L g1768 ( .A(n_1709), .B(n_1712), .Y(n_1768) );
AND2x2_ASAP7_75t_L g1709 ( .A(n_1710), .B(n_1711), .Y(n_1709) );
AND2x2_ASAP7_75t_L g1731 ( .A(n_1712), .B(n_1732), .Y(n_1731) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1712), .Y(n_1743) );
NAND2xp5_ASAP7_75t_L g1797 ( .A(n_1716), .B(n_1798), .Y(n_1797) );
AND2x2_ASAP7_75t_L g1876 ( .A(n_1716), .B(n_1865), .Y(n_1876) );
AND2x2_ASAP7_75t_L g1716 ( .A(n_1717), .B(n_1725), .Y(n_1716) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1717), .B(n_1734), .Y(n_1744) );
AND2x2_ASAP7_75t_L g1745 ( .A(n_1717), .B(n_1746), .Y(n_1745) );
AND2x2_ASAP7_75t_L g1757 ( .A(n_1717), .B(n_1758), .Y(n_1757) );
OR2x2_ASAP7_75t_L g1790 ( .A(n_1717), .B(n_1725), .Y(n_1790) );
INVx3_ASAP7_75t_L g1792 ( .A(n_1717), .Y(n_1792) );
AOI21xp5_ASAP7_75t_L g1884 ( .A1(n_1717), .A2(n_1885), .B(n_1888), .Y(n_1884) );
INVx3_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
OR2x2_ASAP7_75t_L g1751 ( .A(n_1718), .B(n_1752), .Y(n_1751) );
AND2x2_ASAP7_75t_L g1883 ( .A(n_1718), .B(n_1725), .Y(n_1883) );
OR2x2_ASAP7_75t_L g1718 ( .A(n_1719), .B(n_1722), .Y(n_1718) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_1725), .B(n_1735), .Y(n_1734) );
OR2x2_ASAP7_75t_L g1752 ( .A(n_1725), .B(n_1735), .Y(n_1752) );
INVx2_ASAP7_75t_L g1758 ( .A(n_1725), .Y(n_1758) );
AND2x2_ASAP7_75t_L g1762 ( .A(n_1725), .B(n_1746), .Y(n_1762) );
OR2x2_ASAP7_75t_L g1773 ( .A(n_1725), .B(n_1746), .Y(n_1773) );
AOI22xp5_ASAP7_75t_L g1826 ( .A1(n_1725), .A2(n_1794), .B1(n_1827), .B2(n_1831), .Y(n_1826) );
OAI221xp5_ASAP7_75t_L g1853 ( .A1(n_1725), .A2(n_1852), .B1(n_1854), .B2(n_1862), .C(n_1864), .Y(n_1853) );
AND2x4_ASAP7_75t_L g1725 ( .A(n_1726), .B(n_1727), .Y(n_1725) );
OAI21xp5_ASAP7_75t_SL g1728 ( .A1(n_1729), .A2(n_1733), .B(n_1739), .Y(n_1728) );
NAND2xp5_ASAP7_75t_L g1791 ( .A(n_1730), .B(n_1792), .Y(n_1791) );
A2O1A1Ixp33_ASAP7_75t_SL g1823 ( .A1(n_1730), .A2(n_1824), .B(n_1826), .C(n_1834), .Y(n_1823) );
AOI211xp5_ASAP7_75t_L g1854 ( .A1(n_1730), .A2(n_1855), .B(n_1857), .C(n_1861), .Y(n_1854) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1731), .Y(n_1750) );
NAND2xp5_ASAP7_75t_L g1764 ( .A(n_1731), .B(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1734), .Y(n_1733) );
AOI322xp5_ASAP7_75t_L g1804 ( .A1(n_1734), .A2(n_1757), .A3(n_1805), .B1(n_1807), .B2(n_1810), .C1(n_1813), .C2(n_1818), .Y(n_1804) );
INVx2_ASAP7_75t_SL g1746 ( .A(n_1735), .Y(n_1746) );
HB1xp67_ASAP7_75t_L g1756 ( .A(n_1735), .Y(n_1756) );
AOI22xp5_ASAP7_75t_L g1739 ( .A1(n_1740), .A2(n_1744), .B1(n_1745), .B2(n_1747), .Y(n_1739) );
INVxp67_ASAP7_75t_L g1895 ( .A(n_1740), .Y(n_1895) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1741), .B(n_1742), .Y(n_1740) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1742), .Y(n_1806) );
NOR2xp33_ASAP7_75t_L g1889 ( .A(n_1742), .B(n_1890), .Y(n_1889) );
INVx1_ASAP7_75t_L g1873 ( .A(n_1745), .Y(n_1873) );
INVx2_ASAP7_75t_SL g1784 ( .A(n_1746), .Y(n_1784) );
NOR2xp33_ASAP7_75t_L g1749 ( .A(n_1750), .B(n_1751), .Y(n_1749) );
AND2x2_ASAP7_75t_L g1805 ( .A(n_1750), .B(n_1806), .Y(n_1805) );
INVx1_ASAP7_75t_L g1818 ( .A(n_1751), .Y(n_1818) );
INVx1_ASAP7_75t_L g1836 ( .A(n_1752), .Y(n_1836) );
OAI21xp33_ASAP7_75t_SL g1847 ( .A1(n_1752), .A2(n_1848), .B(n_1850), .Y(n_1847) );
AOI21xp5_ASAP7_75t_L g1753 ( .A1(n_1754), .A2(n_1759), .B(n_1761), .Y(n_1753) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
NAND2xp5_ASAP7_75t_L g1755 ( .A(n_1756), .B(n_1757), .Y(n_1755) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1756), .Y(n_1787) );
NAND2xp5_ASAP7_75t_L g1802 ( .A(n_1756), .B(n_1803), .Y(n_1802) );
NAND2xp5_ASAP7_75t_L g1831 ( .A(n_1756), .B(n_1832), .Y(n_1831) );
INVx1_ASAP7_75t_L g1852 ( .A(n_1756), .Y(n_1852) );
INVx1_ASAP7_75t_L g1859 ( .A(n_1756), .Y(n_1859) );
AOI211xp5_ASAP7_75t_SL g1874 ( .A1(n_1757), .A2(n_1875), .B(n_1876), .C(n_1877), .Y(n_1874) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
A2O1A1Ixp33_ASAP7_75t_L g1870 ( .A1(n_1760), .A2(n_1871), .B(n_1873), .C(n_1874), .Y(n_1870) );
AND2x2_ASAP7_75t_L g1761 ( .A(n_1762), .B(n_1763), .Y(n_1761) );
NAND2xp5_ASAP7_75t_L g1774 ( .A(n_1762), .B(n_1775), .Y(n_1774) );
AOI21xp5_ASAP7_75t_L g1834 ( .A1(n_1762), .A2(n_1835), .B(n_1836), .Y(n_1834) );
INVx1_ASAP7_75t_L g1840 ( .A(n_1762), .Y(n_1840) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
NOR2xp33_ASAP7_75t_L g1796 ( .A(n_1764), .B(n_1797), .Y(n_1796) );
NAND2xp5_ASAP7_75t_L g1789 ( .A(n_1765), .B(n_1767), .Y(n_1789) );
NAND2xp5_ASAP7_75t_L g1766 ( .A(n_1767), .B(n_1769), .Y(n_1766) );
NAND2xp5_ASAP7_75t_L g1776 ( .A(n_1767), .B(n_1777), .Y(n_1776) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1768), .Y(n_1767) );
OAI211xp5_ASAP7_75t_L g1819 ( .A1(n_1769), .A2(n_1792), .B(n_1820), .C(n_1821), .Y(n_1819) );
INVx1_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
OR2x2_ASAP7_75t_L g1770 ( .A(n_1771), .B(n_1773), .Y(n_1770) );
NAND2xp5_ASAP7_75t_L g1814 ( .A(n_1771), .B(n_1815), .Y(n_1814) );
AND2x2_ASAP7_75t_L g1832 ( .A(n_1771), .B(n_1833), .Y(n_1832) );
NOR2x1_ASAP7_75t_L g1865 ( .A(n_1771), .B(n_1822), .Y(n_1865) );
INVx2_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
NAND2xp5_ASAP7_75t_L g1782 ( .A(n_1772), .B(n_1783), .Y(n_1782) );
AND2x2_ASAP7_75t_L g1875 ( .A(n_1772), .B(n_1779), .Y(n_1875) );
INVx2_ASAP7_75t_L g1794 ( .A(n_1773), .Y(n_1794) );
AND2x2_ASAP7_75t_L g1851 ( .A(n_1775), .B(n_1852), .Y(n_1851) );
INVx1_ASAP7_75t_L g1775 ( .A(n_1776), .Y(n_1775) );
NOR2xp33_ASAP7_75t_L g1887 ( .A(n_1776), .B(n_1852), .Y(n_1887) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1777), .Y(n_1812) );
NAND2xp5_ASAP7_75t_L g1778 ( .A(n_1779), .B(n_1781), .Y(n_1778) );
INVx1_ASAP7_75t_L g1779 ( .A(n_1780), .Y(n_1779) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1782), .Y(n_1781) );
INVx1_ASAP7_75t_L g1783 ( .A(n_1784), .Y(n_1783) );
INVx1_ASAP7_75t_L g1798 ( .A(n_1784), .Y(n_1798) );
OAI21xp33_ASAP7_75t_L g1885 ( .A1(n_1784), .A2(n_1811), .B(n_1886), .Y(n_1885) );
OAI221xp5_ASAP7_75t_L g1785 ( .A1(n_1786), .A2(n_1790), .B1(n_1791), .B2(n_1793), .C(n_1795), .Y(n_1785) );
NAND2xp5_ASAP7_75t_L g1786 ( .A(n_1787), .B(n_1788), .Y(n_1786) );
INVx1_ASAP7_75t_L g1788 ( .A(n_1789), .Y(n_1788) );
INVx1_ASAP7_75t_SL g1801 ( .A(n_1792), .Y(n_1801) );
NOR3xp33_ASAP7_75t_L g1877 ( .A(n_1792), .B(n_1806), .C(n_1856), .Y(n_1877) );
INVxp67_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
NOR2xp33_ASAP7_75t_L g1828 ( .A(n_1798), .B(n_1829), .Y(n_1828) );
OAI211xp5_ASAP7_75t_SL g1799 ( .A1(n_1800), .A2(n_1802), .B(n_1804), .C(n_1819), .Y(n_1799) );
OAI311xp33_ASAP7_75t_L g1837 ( .A1(n_1800), .A2(n_1838), .A3(n_1839), .B1(n_1847), .C1(n_1853), .Y(n_1837) );
INVx1_ASAP7_75t_L g1842 ( .A(n_1803), .Y(n_1842) );
OR2x2_ASAP7_75t_L g1811 ( .A(n_1806), .B(n_1812), .Y(n_1811) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1808), .Y(n_1807) );
INVx1_ASAP7_75t_L g1810 ( .A(n_1811), .Y(n_1810) );
NAND2xp33_ASAP7_75t_L g1813 ( .A(n_1814), .B(n_1816), .Y(n_1813) );
INVx1_ASAP7_75t_L g1816 ( .A(n_1817), .Y(n_1816) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1822), .Y(n_1821) );
INVx1_ASAP7_75t_L g1824 ( .A(n_1825), .Y(n_1824) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1828), .Y(n_1827) );
INVx1_ASAP7_75t_L g1861 ( .A(n_1829), .Y(n_1861) );
INVx1_ASAP7_75t_L g1838 ( .A(n_1831), .Y(n_1838) );
INVxp67_ASAP7_75t_L g1881 ( .A(n_1832), .Y(n_1881) );
OAI21xp33_ASAP7_75t_L g1839 ( .A1(n_1840), .A2(n_1841), .B(n_1845), .Y(n_1839) );
AND2x2_ASAP7_75t_L g1841 ( .A(n_1842), .B(n_1843), .Y(n_1841) );
INVx1_ASAP7_75t_L g1843 ( .A(n_1844), .Y(n_1843) );
INVx1_ASAP7_75t_L g1848 ( .A(n_1849), .Y(n_1848) );
A2O1A1Ixp33_ASAP7_75t_L g1880 ( .A1(n_1850), .A2(n_1881), .B(n_1882), .C(n_1884), .Y(n_1880) );
INVx1_ASAP7_75t_L g1850 ( .A(n_1851), .Y(n_1850) );
INVx1_ASAP7_75t_L g1855 ( .A(n_1856), .Y(n_1855) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1858), .Y(n_1857) );
NAND2xp5_ASAP7_75t_L g1858 ( .A(n_1859), .B(n_1860), .Y(n_1858) );
INVx1_ASAP7_75t_L g1868 ( .A(n_1863), .Y(n_1868) );
NAND2xp5_ASAP7_75t_L g1866 ( .A(n_1867), .B(n_1868), .Y(n_1866) );
AOI21xp5_ASAP7_75t_L g1869 ( .A1(n_1870), .A2(n_1878), .B(n_1880), .Y(n_1869) );
CKINVDCx14_ASAP7_75t_R g1878 ( .A(n_1879), .Y(n_1878) );
INVx1_ASAP7_75t_L g1882 ( .A(n_1883), .Y(n_1882) );
INVxp33_ASAP7_75t_L g1886 ( .A(n_1887), .Y(n_1886) );
INVx1_ASAP7_75t_L g1892 ( .A(n_1893), .Y(n_1892) );
INVx1_ASAP7_75t_L g1896 ( .A(n_1897), .Y(n_1896) );
INVx2_ASAP7_75t_L g1898 ( .A(n_1899), .Y(n_1898) );
XNOR2x1_ASAP7_75t_L g1899 ( .A(n_1900), .B(n_1901), .Y(n_1899) );
AND2x2_ASAP7_75t_L g1901 ( .A(n_1902), .B(n_1926), .Y(n_1901) );
NOR3xp33_ASAP7_75t_SL g1902 ( .A(n_1903), .B(n_1909), .C(n_1911), .Y(n_1902) );
AOI221xp5_ASAP7_75t_L g1937 ( .A1(n_1924), .A2(n_1938), .B1(n_1940), .B2(n_1943), .C(n_1944), .Y(n_1937) );
AOI21xp5_ASAP7_75t_L g1926 ( .A1(n_1927), .A2(n_1929), .B(n_1930), .Y(n_1926) );
INVx1_ASAP7_75t_L g1927 ( .A(n_1928), .Y(n_1927) );
INVx1_ASAP7_75t_L g1938 ( .A(n_1939), .Y(n_1938) );
INVx1_ASAP7_75t_L g1944 ( .A(n_1945), .Y(n_1944) );
INVx4_ASAP7_75t_SL g1947 ( .A(n_1948), .Y(n_1947) );
BUFx3_ASAP7_75t_L g1948 ( .A(n_1949), .Y(n_1948) );
BUFx2_ASAP7_75t_L g1949 ( .A(n_1950), .Y(n_1949) );
BUFx2_ASAP7_75t_L g1952 ( .A(n_1953), .Y(n_1952) );
A2O1A1Ixp33_ASAP7_75t_L g1959 ( .A1(n_1954), .A2(n_1960), .B(n_1962), .C(n_1964), .Y(n_1959) );
INVxp33_ASAP7_75t_SL g1955 ( .A(n_1956), .Y(n_1955) );
BUFx2_ASAP7_75t_L g1957 ( .A(n_1958), .Y(n_1957) );
HB1xp67_ASAP7_75t_L g1958 ( .A(n_1959), .Y(n_1958) );
INVx1_ASAP7_75t_L g1960 ( .A(n_1961), .Y(n_1960) );
INVx1_ASAP7_75t_L g1962 ( .A(n_1963), .Y(n_1962) );
endmodule