module fake_jpeg_23376_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_21),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_37),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_33),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_21),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_23),
.B1(n_25),
.B2(n_28),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_23),
.B1(n_25),
.B2(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_51),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_65),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_68),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_81),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_72),
.B1(n_75),
.B2(n_79),
.Y(n_99)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_67),
.Y(n_96)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_47),
.Y(n_109)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_48),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_38),
.B1(n_57),
.B2(n_23),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_38),
.B1(n_26),
.B2(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_17),
.Y(n_78)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_34),
.C(n_36),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_34),
.C(n_27),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_17),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_25),
.B1(n_31),
.B2(n_29),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_29),
.B1(n_51),
.B2(n_27),
.Y(n_91)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_89),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_58),
.B(n_32),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_32),
.B(n_17),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_70),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_106),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_98),
.B1(n_104),
.B2(n_65),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_62),
.CI(n_72),
.CON(n_94),
.SN(n_94)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_102),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_32),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_97),
.B(n_9),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_37),
.B1(n_34),
.B2(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_47),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_58),
.A2(n_37),
.B1(n_34),
.B2(n_30),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_34),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_76),
.B(n_34),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_71),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_58),
.A2(n_30),
.B1(n_27),
.B2(n_48),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_110),
.A2(n_111),
.B1(n_76),
.B2(n_82),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_68),
.A2(n_16),
.B1(n_24),
.B2(n_22),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_69),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_117),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_122),
.B1(n_89),
.B2(n_102),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_81),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_118),
.B(n_120),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_70),
.B1(n_83),
.B2(n_73),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_119),
.A2(n_107),
.B1(n_1),
.B2(n_3),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_83),
.B1(n_74),
.B2(n_73),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_137),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_127),
.B(n_101),
.Y(n_160)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_125),
.B(n_131),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_22),
.B(n_19),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_74),
.B1(n_60),
.B2(n_19),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_18),
.B1(n_16),
.B2(n_32),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_97),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_136),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_86),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_111),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_90),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_10),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_10),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_100),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_88),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_142),
.C(n_151),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_162),
.B1(n_165),
.B2(n_3),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_105),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_106),
.B(n_94),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_145),
.A2(n_146),
.B(n_163),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_110),
.B(n_90),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_148),
.B(n_162),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_94),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_161),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_103),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_152),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_113),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_154),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_103),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_101),
.Y(n_157)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_112),
.B(n_10),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_122),
.B(n_126),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_129),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_0),
.B(n_1),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_142),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_175),
.C(n_176),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_150),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_141),
.B1(n_164),
.B2(n_154),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_163),
.A2(n_135),
.B1(n_115),
.B2(n_121),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_158),
.B1(n_149),
.B2(n_153),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_183),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_137),
.C(n_121),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_127),
.C(n_5),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_8),
.B(n_11),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_3),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_SL g194 ( 
.A(n_179),
.B(n_180),
.C(n_140),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_181),
.A2(n_144),
.B1(n_165),
.B2(n_148),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_157),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_159),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_161),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_188),
.B(n_205),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_144),
.B1(n_146),
.B2(n_155),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_191),
.B1(n_196),
.B2(n_177),
.Y(n_215)
);

FAx1_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_153),
.CI(n_160),
.CON(n_192),
.SN(n_192)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_198),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_202),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_179),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_199),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_151),
.B(n_8),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_7),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_204),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_11),
.B(n_12),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_171),
.B(n_12),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_187),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_12),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_209),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_211),
.Y(n_222)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_173),
.C(n_175),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_212),
.C(n_213),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_173),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_186),
.C(n_166),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_186),
.C(n_166),
.Y(n_213)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_168),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_225),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_192),
.B1(n_200),
.B2(n_203),
.Y(n_223)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_189),
.B1(n_192),
.B2(n_174),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_224),
.Y(n_232)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_217),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_219),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_174),
.C(n_193),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_230),
.C(n_207),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_205),
.C(n_184),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_231),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_235),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_220),
.A2(n_207),
.B1(n_206),
.B2(n_201),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_237),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_226),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_228),
.A2(n_211),
.B(n_202),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_228),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_223),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_241),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_243),
.B(n_245),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_230),
.B(n_222),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_236),
.B(n_234),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_248),
.B(n_249),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_238),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_240),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_242),
.C(n_14),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_247),
.B(n_235),
.Y(n_252)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_252),
.A2(n_13),
.B(n_15),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_253),
.A2(n_254),
.B(n_251),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_15),
.Y(n_256)
);


endmodule