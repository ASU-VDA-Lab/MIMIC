module fake_jpeg_32044_n_533 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_533);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_533;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_6),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_52),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_22),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_53),
.B(n_56),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_57),
.B(n_69),
.Y(n_152)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_61),
.B(n_90),
.Y(n_164)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_17),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_74),
.B(n_81),
.Y(n_107)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_24),
.B(n_17),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_39),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_91),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_24),
.B(n_50),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_96),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_19),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_100),
.A2(n_31),
.B1(n_36),
.B2(n_49),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_39),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_101),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_64),
.B1(n_59),
.B2(n_63),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_103),
.A2(n_124),
.B1(n_142),
.B2(n_104),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_104),
.A2(n_142),
.B1(n_88),
.B2(n_80),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_54),
.A2(n_34),
.B1(n_47),
.B2(n_46),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

BUFx4f_ASAP7_75t_L g137 ( 
.A(n_55),
.Y(n_137)
);

BUFx24_ASAP7_75t_L g210 ( 
.A(n_137),
.Y(n_210)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_75),
.A2(n_72),
.B1(n_19),
.B2(n_48),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

BUFx16f_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_89),
.B(n_28),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_37),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_60),
.Y(n_155)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_77),
.Y(n_156)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_99),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_159),
.B(n_25),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_91),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_163),
.Y(n_178)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_166),
.A2(n_215),
.B1(n_0),
.B2(n_1),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_167),
.B(n_168),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_49),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_169),
.Y(n_236)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_170),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_37),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_172),
.B(n_179),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_173),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_177),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_108),
.Y(n_179)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_181),
.Y(n_271)
);

OR2x2_ASAP7_75t_SL g182 ( 
.A(n_144),
.B(n_100),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_182),
.A2(n_192),
.B(n_205),
.Y(n_276)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_127),
.Y(n_186)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_108),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_189),
.B(n_191),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_40),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_204),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_126),
.B(n_40),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_148),
.B(n_32),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_194),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_195),
.A2(n_103),
.B1(n_117),
.B2(n_150),
.Y(n_226)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_111),
.Y(n_197)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_197),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_126),
.B(n_152),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_218),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_152),
.A2(n_71),
.B(n_85),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_199),
.A2(n_145),
.B(n_151),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_109),
.A2(n_71),
.B1(n_85),
.B2(n_55),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_200),
.A2(n_223),
.B1(n_43),
.B2(n_147),
.Y(n_265)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_105),
.Y(n_201)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_202),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_132),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_203),
.Y(n_248)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_149),
.B(n_31),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_114),
.B(n_123),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_207),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_137),
.Y(n_207)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_133),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_208),
.B(n_209),
.Y(n_270)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_135),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_211),
.B(n_213),
.Y(n_273)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

NAND2x1_ASAP7_75t_SL g238 ( 
.A(n_212),
.B(n_115),
.Y(n_238)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_136),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_110),
.B(n_128),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_221),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_121),
.A2(n_67),
.B1(n_65),
.B2(n_97),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_SL g216 ( 
.A1(n_124),
.A2(n_92),
.B(n_48),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_94),
.C(n_131),
.Y(n_255)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_217),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_110),
.B(n_36),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_133),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_143),
.B(n_27),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_119),
.B(n_44),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_48),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_115),
.A2(n_66),
.B1(n_48),
.B2(n_43),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_224),
.Y(n_264)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_138),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_225),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_226),
.B(n_238),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_162),
.B(n_157),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_231),
.A2(n_243),
.B(n_244),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_166),
.A2(n_125),
.B1(n_150),
.B2(n_138),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_235),
.A2(n_258),
.B1(n_210),
.B2(n_3),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_41),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_237),
.B(n_241),
.C(n_263),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_47),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_41),
.B(n_44),
.C(n_46),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_178),
.A2(n_180),
.B(n_171),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_255),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_183),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_251),
.B(n_253),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_215),
.A2(n_131),
.B1(n_25),
.B2(n_27),
.Y(n_254)
);

AOI32xp33_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_208),
.A3(n_169),
.B1(n_170),
.B2(n_185),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_223),
.A2(n_66),
.B1(n_48),
.B2(n_43),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_261),
.A2(n_186),
.B1(n_219),
.B2(n_203),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_165),
.B(n_43),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_220),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_183),
.B(n_163),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_265),
.A2(n_266),
.B1(n_2),
.B2(n_4),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_181),
.A2(n_43),
.B1(n_27),
.B2(n_25),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_183),
.B(n_27),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_275),
.C(n_201),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_175),
.B(n_176),
.Y(n_275)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_274),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_277),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_SL g326 ( 
.A1(n_278),
.A2(n_238),
.B(n_263),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_279),
.B(n_283),
.Y(n_325)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_282),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_187),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_285),
.B(n_272),
.Y(n_343)
);

OR2x4_ASAP7_75t_L g286 ( 
.A(n_231),
.B(n_200),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g360 ( 
.A1(n_286),
.A2(n_283),
.B(n_320),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_256),
.B(n_212),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_288),
.B(n_291),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_289),
.A2(n_290),
.B1(n_300),
.B2(n_320),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_261),
.A2(n_173),
.B1(n_202),
.B2(n_174),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_234),
.B(n_197),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_232),
.B(n_220),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_293),
.B(n_295),
.Y(n_361)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_294),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_250),
.B(n_15),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_296),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_228),
.B(n_1),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_297),
.B(n_302),
.Y(n_362)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_298),
.Y(n_329)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_299),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_264),
.A2(n_174),
.B1(n_210),
.B2(n_27),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_239),
.Y(n_301)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_301),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_228),
.B(n_25),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_227),
.B(n_25),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_307),
.Y(n_355)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_304),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_255),
.B(n_210),
.C(n_14),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_305),
.B(n_267),
.C(n_262),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_306),
.A2(n_308),
.B1(n_286),
.B2(n_318),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_242),
.B(n_11),
.Y(n_307)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_309),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_273),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_319),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g311 ( 
.A(n_276),
.B(n_10),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_311),
.A2(n_323),
.B(n_7),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_242),
.B(n_268),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_312),
.Y(n_324)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_271),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_314),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_241),
.B(n_2),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g336 ( 
.A(n_315),
.B(n_318),
.CI(n_260),
.CON(n_336),
.SN(n_336)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_235),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_316),
.A2(n_249),
.B1(n_236),
.B2(n_260),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_247),
.B(n_5),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_317),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_264),
.B(n_5),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_252),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_226),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_244),
.B(n_6),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_321),
.B(n_237),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_249),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_322),
.A2(n_248),
.B1(n_236),
.B2(n_257),
.Y(n_350)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_243),
.B(n_7),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_326),
.A2(n_346),
.B1(n_352),
.B2(n_313),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_327),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_292),
.A2(n_258),
.B(n_254),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_330),
.A2(n_337),
.B(n_339),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_335),
.B(n_336),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_280),
.A2(n_245),
.B(n_246),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_280),
.A2(n_246),
.B(n_259),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_292),
.A2(n_290),
.B1(n_289),
.B2(n_281),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_340),
.A2(n_342),
.B1(n_351),
.B2(n_285),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_292),
.A2(n_233),
.B1(n_230),
.B2(n_229),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_349),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_345),
.A2(n_350),
.B1(n_298),
.B2(n_309),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_284),
.B(n_259),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_281),
.A2(n_233),
.B1(n_248),
.B2(n_257),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_306),
.A2(n_248),
.B1(n_252),
.B2(n_10),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_311),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_284),
.A2(n_9),
.B(n_305),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_356),
.B(n_359),
.Y(n_375)
);

OA22x2_ASAP7_75t_L g357 ( 
.A1(n_294),
.A2(n_9),
.B1(n_296),
.B2(n_287),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_360),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_279),
.A2(n_9),
.B(n_323),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_365),
.B(n_378),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_366),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_334),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_368),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_325),
.B(n_297),
.Y(n_371)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_371),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_315),
.C(n_299),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_372),
.B(n_389),
.C(n_336),
.Y(n_406)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_358),
.Y(n_374)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_310),
.Y(n_376)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_347),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_377),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_324),
.B(n_301),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_304),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_391),
.Y(n_413)
);

CKINVDCx12_ASAP7_75t_R g380 ( 
.A(n_344),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_380),
.B(n_393),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_381),
.B(n_394),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_382),
.A2(n_332),
.B1(n_337),
.B2(n_330),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_319),
.Y(n_383)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_383),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_322),
.Y(n_385)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_385),
.Y(n_423)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_386),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_314),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_388),
.Y(n_400)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_344),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_335),
.B(n_277),
.C(n_282),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_333),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_390),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_336),
.B(n_356),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_340),
.A2(n_332),
.B1(n_339),
.B2(n_351),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_396),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_324),
.B(n_331),
.Y(n_393)
);

INVx13_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_331),
.B(n_362),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_395),
.B(n_355),
.Y(n_409)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_338),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_334),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_397),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_357),
.B(n_341),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_357),
.Y(n_422)
);

BUFx10_ASAP7_75t_L g399 ( 
.A(n_354),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_399),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_403),
.A2(n_414),
.B1(n_384),
.B2(n_352),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_406),
.B(n_391),
.Y(n_439)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_409),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_377),
.A2(n_364),
.B1(n_329),
.B2(n_354),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_410),
.A2(n_354),
.B1(n_363),
.B2(n_387),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_390),
.B(n_361),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_411),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_382),
.A2(n_338),
.B1(n_341),
.B2(n_342),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_367),
.B(n_327),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_416),
.B(n_370),
.Y(n_445)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_422),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_367),
.B(n_389),
.C(n_372),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_428),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_376),
.B(n_348),
.Y(n_425)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_425),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_384),
.A2(n_359),
.B(n_353),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_427),
.A2(n_388),
.B(n_396),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_379),
.B(n_363),
.C(n_364),
.Y(n_428)
);

OAI21xp33_ASAP7_75t_L g430 ( 
.A1(n_412),
.A2(n_385),
.B(n_383),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_435),
.Y(n_465)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_425),
.Y(n_433)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_433),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_413),
.B(n_373),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_436),
.A2(n_440),
.B1(n_448),
.B2(n_423),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_421),
.B(n_392),
.Y(n_437)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_437),
.Y(n_475)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_402),
.Y(n_438)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_427),
.C(n_414),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_423),
.A2(n_370),
.B1(n_398),
.B2(n_375),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_426),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_441),
.B(n_443),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_365),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_445),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_400),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_446),
.A2(n_454),
.B1(n_417),
.B2(n_443),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_413),
.B(n_371),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_449),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_417),
.A2(n_419),
.B1(n_412),
.B2(n_401),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_406),
.B(n_369),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_408),
.Y(n_450)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_450),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_422),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_419),
.B(n_374),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_415),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_403),
.A2(n_386),
.B1(n_368),
.B2(n_397),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_404),
.B(n_329),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_455),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_428),
.C(n_416),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_463),
.C(n_466),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_457),
.B(n_394),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_458),
.A2(n_446),
.B1(n_431),
.B2(n_415),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_404),
.C(n_400),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_471),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_407),
.C(n_418),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_407),
.C(n_418),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_470),
.C(n_476),
.Y(n_491)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_439),
.B(n_447),
.C(n_437),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_429),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_473),
.A2(n_440),
.B1(n_444),
.B2(n_408),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_455),
.C(n_432),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_488),
.Y(n_500)
);

AO21x1_ASAP7_75t_L g478 ( 
.A1(n_475),
.A2(n_430),
.B(n_434),
.Y(n_478)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_478),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_481),
.A2(n_459),
.B1(n_399),
.B2(n_460),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_461),
.B(n_450),
.Y(n_482)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_482),
.Y(n_505)
);

INVx13_ASAP7_75t_L g483 ( 
.A(n_474),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_483),
.B(n_485),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_474),
.A2(n_429),
.B(n_411),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_484),
.A2(n_492),
.B(n_482),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_467),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_476),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_487),
.Y(n_504)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_472),
.Y(n_487)
);

INVx13_ASAP7_75t_L g490 ( 
.A(n_462),
.Y(n_490)
);

NAND3xp33_ASAP7_75t_SL g497 ( 
.A(n_490),
.B(n_493),
.C(n_399),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_463),
.A2(n_405),
.B(n_420),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_468),
.Y(n_493)
);

FAx1_ASAP7_75t_SL g494 ( 
.A(n_481),
.B(n_465),
.CI(n_466),
.CON(n_494),
.SN(n_494)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_497),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_486),
.A2(n_470),
.B(n_465),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_496),
.A2(n_480),
.B(n_479),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_491),
.A2(n_456),
.B(n_409),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_498),
.B(n_480),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_478),
.A2(n_405),
.B(n_420),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_506),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_501),
.A2(n_477),
.B1(n_485),
.B2(n_482),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_399),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_492),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_503),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_491),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_509),
.B(n_512),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_510),
.B(n_511),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_504),
.B(n_489),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_514),
.B(n_515),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_484),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_502),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_519),
.B(n_509),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_508),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_507),
.A2(n_506),
.B(n_495),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_521),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_523),
.B(n_524),
.Y(n_527)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_516),
.Y(n_525)
);

NOR3xp33_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_518),
.C(n_517),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_526),
.B(n_522),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_527),
.B(n_499),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_513),
.Y(n_530)
);

AO21x1_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_487),
.B(n_505),
.Y(n_531)
);

MAJx2_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_490),
.C(n_483),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_494),
.B1(n_524),
.B2(n_525),
.Y(n_533)
);


endmodule