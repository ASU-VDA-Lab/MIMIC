module real_jpeg_30832_n_19 (n_17, n_8, n_0, n_141, n_2, n_142, n_143, n_10, n_9, n_12, n_147, n_146, n_6, n_151, n_11, n_14, n_7, n_18, n_3, n_145, n_144, n_5, n_4, n_150, n_1, n_148, n_149, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_141;
input n_2;
input n_142;
input n_143;
input n_10;
input n_9;
input n_12;
input n_147;
input n_146;
input n_6;
input n_151;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_145;
input n_144;
input n_5;
input n_4;
input n_150;
input n_1;
input n_148;
input n_149;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx1_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_0),
.B(n_63),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_2),
.B(n_69),
.Y(n_68)
);

HAxp5_ASAP7_75t_SL g119 ( 
.A(n_2),
.B(n_69),
.CON(n_119),
.SN(n_119)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_4),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_5),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_5),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_6),
.B(n_36),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_7),
.B(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_8),
.B(n_35),
.Y(n_127)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_10),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_10),
.Y(n_134)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

AOI322xp5_ASAP7_75t_L g121 ( 
.A1(n_11),
.A2(n_52),
.A3(n_54),
.B1(n_61),
.B2(n_122),
.C1(n_124),
.C2(n_151),
.Y(n_121)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_13),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_13),
.B(n_113),
.Y(n_123)
);

AOI221xp5_ASAP7_75t_L g83 ( 
.A1(n_14),
.A2(n_16),
.B1(n_84),
.B2(n_89),
.C(n_93),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_14),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_16),
.B(n_84),
.C(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_18),
.B(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_136),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_130),
.B(n_133),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_32),
.B(n_128),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_31),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_24),
.B(n_31),
.Y(n_129)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_27),
.Y(n_138)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_40),
.B(n_127),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_39),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI31xp67_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_74),
.A3(n_111),
.B(n_117),
.Y(n_41)
);

NOR3xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_60),
.C(n_68),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_43),
.A2(n_118),
.B(n_121),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_52),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_45),
.B(n_68),
.C(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_46),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_142),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

OA21x2_ASAP7_75t_SL g118 ( 
.A1(n_60),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_67),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_105),
.C(n_106),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_97),
.B(n_104),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_83),
.B1(n_95),
.B2(n_96),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_147),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_103),
.Y(n_104)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_141),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_143),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_144),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_145),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_146),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_148),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_149),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_150),
.Y(n_114)
);


endmodule