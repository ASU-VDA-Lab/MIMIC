module fake_jpeg_10675_n_75 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_75);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_75;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_3),
.B(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_21),
.B(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_0),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_9),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_11),
.B1(n_19),
.B2(n_18),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_11),
.B1(n_13),
.B2(n_6),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_10),
.B(n_16),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_29),
.A2(n_31),
.B(n_5),
.Y(n_45)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_21),
.A2(n_10),
.B(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_9),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_14),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_47),
.Y(n_55)
);

OAI21x1_ASAP7_75t_SL g47 ( 
.A1(n_28),
.A2(n_34),
.B(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_53),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_58),
.Y(n_65)
);

AND2x6_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_45),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_60),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_33),
.C(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_60),
.C(n_51),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_68),
.C(n_63),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_67),
.B(n_65),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_70),
.B(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_53),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_7),
.Y(n_75)
);


endmodule