module fake_jpeg_1331_n_262 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_17),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_24),
.B(n_19),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_43),
.A2(n_32),
.B(n_30),
.Y(n_86)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_20),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_65),
.Y(n_69)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_1),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_31),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_38),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_79),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_43),
.A2(n_36),
.B1(n_23),
.B2(n_34),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_68),
.B1(n_49),
.B2(n_47),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_36),
.B1(n_23),
.B2(n_34),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_80),
.B(n_81),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_87),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_38),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_91),
.B(n_51),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_66),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_93),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_46),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_63),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_57),
.A2(n_28),
.B1(n_22),
.B2(n_32),
.Y(n_101)
);

AO22x1_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_58),
.B1(n_61),
.B2(n_56),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_28),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_104),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_129),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_26),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_73),
.B1(n_95),
.B2(n_90),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

BUFx4f_ASAP7_75t_SL g141 ( 
.A(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_108),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_26),
.B1(n_30),
.B2(n_59),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_56),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_132),
.C(n_77),
.Y(n_143)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_128),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_123),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_70),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_122),
.B(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_60),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_55),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_89),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_76),
.B(n_12),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_73),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_88),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_133),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_56),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_95),
.B(n_15),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_149),
.C(n_109),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_143),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_71),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_126),
.B(n_89),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_74),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_145),
.Y(n_162)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_113),
.A2(n_132),
.B(n_111),
.Y(n_158)
);

AOI21x1_ASAP7_75t_SL g177 ( 
.A1(n_158),
.A2(n_128),
.B(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_162),
.B(n_179),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_113),
.C(n_103),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_166),
.C(n_174),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_134),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_165),
.B(n_183),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_142),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_145),
.A2(n_119),
.B1(n_123),
.B2(n_124),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_136),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_113),
.B1(n_109),
.B2(n_104),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_175),
.B1(n_181),
.B2(n_144),
.Y(n_187)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_184),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_109),
.C(n_130),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_128),
.B1(n_106),
.B2(n_74),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_164),
.Y(n_202)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_159),
.A2(n_72),
.B1(n_117),
.B2(n_112),
.Y(n_181)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_182),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_161),
.A2(n_151),
.B1(n_140),
.B2(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_186),
.B(n_187),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_201),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_177),
.B(n_181),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_163),
.B(n_170),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_144),
.B1(n_139),
.B2(n_154),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_139),
.C(n_147),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_96),
.C(n_83),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_176),
.B(n_138),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_152),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_147),
.Y(n_203)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

AOI21x1_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_187),
.B(n_194),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_169),
.B(n_178),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_205),
.B(n_211),
.Y(n_224)
);

A2O1A1O1Ixp25_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_152),
.B(n_156),
.C(n_137),
.D(n_182),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_SL g222 ( 
.A(n_208),
.B(n_212),
.C(n_193),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_215),
.C(n_185),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_172),
.Y(n_211)
);

OAI322xp33_ASAP7_75t_L g212 ( 
.A1(n_198),
.A2(n_153),
.A3(n_184),
.B1(n_83),
.B2(n_141),
.C1(n_22),
.C2(n_96),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_153),
.B(n_14),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_200),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_197),
.A2(n_189),
.B1(n_202),
.B2(n_203),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_217),
.A2(n_216),
.B1(n_210),
.B2(n_206),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_218),
.B(n_219),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_14),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_222),
.B1(n_225),
.B2(n_231),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_226),
.Y(n_234)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_212),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_185),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_204),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_217),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_200),
.B1(n_193),
.B2(n_191),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_230),
.B(n_207),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_233),
.B(n_238),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_231),
.B(n_223),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_228),
.Y(n_241)
);

NOR3xp33_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_206),
.C(n_210),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_225),
.A2(n_209),
.B1(n_215),
.B2(n_191),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_227),
.B1(n_222),
.B2(n_224),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_242),
.C(n_237),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_236),
.B1(n_232),
.B2(n_238),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_223),
.B(n_188),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_246),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_239),
.A2(n_188),
.B1(n_13),
.B2(n_4),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_252),
.Y(n_255)
);

AOI322xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_22),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_247),
.B(n_83),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_256),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_252),
.A2(n_1),
.B(n_2),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_1),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_257),
.Y(n_260)
);

AOI322xp5_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_253),
.A3(n_22),
.B1(n_5),
.B2(n_9),
.C1(n_4),
.C2(n_2),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_253),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_260),
.Y(n_262)
);


endmodule