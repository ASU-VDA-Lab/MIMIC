module fake_jpeg_15563_n_353 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_21),
.B1(n_32),
.B2(n_36),
.Y(n_69)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_16),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_38),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_68),
.Y(n_104)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_32),
.B1(n_46),
.B2(n_44),
.Y(n_90)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_34),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_21),
.B1(n_36),
.B2(n_18),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_81),
.A2(n_24),
.B1(n_49),
.B2(n_48),
.Y(n_138)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx2_ASAP7_75t_SL g124 ( 
.A(n_82),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_51),
.A3(n_21),
.B1(n_39),
.B2(n_42),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_83),
.A2(n_28),
.A3(n_27),
.B1(n_20),
.B2(n_37),
.Y(n_144)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_88),
.B(n_97),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_42),
.B1(n_46),
.B2(n_41),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_94),
.B1(n_112),
.B2(n_17),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_95),
.B1(n_17),
.B2(n_30),
.Y(n_122)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_96),
.Y(n_119)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_41),
.B1(n_18),
.B2(n_47),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_47),
.B1(n_18),
.B2(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_26),
.Y(n_97)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_32),
.B1(n_52),
.B2(n_50),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_53),
.Y(n_117)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_105),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_27),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_33),
.C(n_29),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_26),
.B(n_17),
.C(n_30),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_101),
.A2(n_102),
.B1(n_24),
.B2(n_33),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_40),
.B1(n_38),
.B2(n_35),
.Y(n_102)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_66),
.B(n_25),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_109),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_40),
.B1(n_22),
.B2(n_38),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_26),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_114),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_68),
.A2(n_22),
.B1(n_35),
.B2(n_34),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_22),
.B1(n_35),
.B2(n_34),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_126),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_144),
.B1(n_84),
.B2(n_103),
.Y(n_155)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_128),
.B1(n_139),
.B2(n_96),
.Y(n_151)
);

NAND2x1_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_53),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_52),
.B1(n_50),
.B2(n_49),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_134),
.C(n_117),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_30),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_98),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_25),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_135),
.B(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_25),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_137),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_138),
.A2(n_91),
.B1(n_99),
.B2(n_84),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_90),
.A2(n_52),
.B1(n_49),
.B2(n_28),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_95),
.A2(n_28),
.B1(n_24),
.B2(n_29),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_140),
.A2(n_79),
.B1(n_37),
.B2(n_33),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_107),
.Y(n_154)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_158),
.Y(n_180)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_151),
.B1(n_155),
.B2(n_159),
.Y(n_194)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_124),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_154),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_104),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_80),
.B1(n_78),
.B2(n_105),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_80),
.B1(n_78),
.B2(n_93),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_161),
.B1(n_171),
.B2(n_173),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_101),
.B1(n_82),
.B2(n_79),
.Y(n_161)
);

BUFx4f_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_167),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_129),
.C(n_130),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_147),
.B(n_162),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_37),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_168),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_27),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_29),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_133),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_136),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_15),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_175),
.Y(n_178)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_170),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_182),
.B(n_196),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_183),
.B(n_192),
.C(n_193),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_176),
.A2(n_137),
.B1(n_140),
.B2(n_120),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_184),
.A2(n_190),
.B1(n_195),
.B2(n_208),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_133),
.B(n_135),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_187),
.A2(n_197),
.B(n_199),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_172),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_120),
.B1(n_146),
.B2(n_119),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_119),
.A3(n_125),
.B1(n_132),
.B2(n_146),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_206),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_123),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_142),
.C(n_118),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_155),
.A2(n_118),
.B1(n_142),
.B2(n_143),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_157),
.A2(n_15),
.B1(n_13),
.B2(n_11),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_0),
.B(n_3),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_162),
.Y(n_200)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_205),
.B1(n_153),
.B2(n_6),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_161),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_15),
.C(n_13),
.Y(n_206)
);

OAI32xp33_ASAP7_75t_L g207 ( 
.A1(n_173),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_207),
.B(n_4),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_157),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_151),
.A2(n_9),
.B1(n_10),
.B2(n_7),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_209),
.A2(n_197),
.B(n_199),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_166),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_183),
.C(n_187),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_186),
.Y(n_245)
);

AOI221xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_174),
.B1(n_172),
.B2(n_168),
.C(n_165),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_150),
.Y(n_214)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_215),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_188),
.B(n_160),
.Y(n_216)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_218),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_156),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_156),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_180),
.A2(n_152),
.B(n_163),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_221),
.A2(n_231),
.B(n_240),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_189),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_223),
.B(n_227),
.C(n_233),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_225),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_180),
.A2(n_153),
.B(n_7),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_189),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

NAND2xp33_ASAP7_75t_SL g238 ( 
.A(n_204),
.B(n_7),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_238),
.A2(n_240),
.B1(n_207),
.B2(n_208),
.Y(n_243)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_243),
.A2(n_251),
.B1(n_228),
.B2(n_231),
.Y(n_276)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_263),
.C(n_222),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_229),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_253),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_194),
.B1(n_179),
.B2(n_193),
.Y(n_251)
);

AOI22x1_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_204),
.B1(n_190),
.B2(n_184),
.Y(n_252)
);

OA21x2_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_244),
.B(n_224),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_235),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_186),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_224),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_215),
.Y(n_257)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_195),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_211),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_206),
.C(n_182),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_228),
.B(n_227),
.Y(n_277)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_221),
.C(n_226),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_269),
.B(n_270),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_265),
.B(n_226),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_216),
.B1(n_205),
.B2(n_233),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_274),
.B1(n_282),
.B2(n_285),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_248),
.B(n_198),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_273),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_277),
.Y(n_292)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_266),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_201),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_281),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_284),
.C(n_286),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_234),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_242),
.A2(n_236),
.B1(n_237),
.B2(n_235),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_251),
.B(n_196),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_252),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_210),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_241),
.A2(n_230),
.B1(n_239),
.B2(n_210),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_245),
.B(n_230),
.C(n_200),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_8),
.C(n_9),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_243),
.C(n_249),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_301),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_264),
.Y(n_294)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_272),
.Y(n_298)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_286),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_303),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_257),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_304),
.C(n_281),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_241),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_305),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_262),
.B1(n_283),
.B2(n_274),
.Y(n_306)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

NAND3xp33_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_269),
.C(n_270),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_316),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_290),
.A2(n_274),
.B1(n_278),
.B2(n_249),
.Y(n_308)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_300),
.A2(n_244),
.B(n_255),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_309),
.A2(n_261),
.B(n_295),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_284),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_255),
.B(n_259),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_295),
.C(n_297),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_258),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_258),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_320),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_248),
.B1(n_246),
.B2(n_256),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_256),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_314),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_324),
.A2(n_317),
.B(n_315),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_326),
.B(n_329),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_296),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_331),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_312),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_324),
.C(n_292),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_337),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_328),
.A2(n_319),
.B1(n_313),
.B2(n_311),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_334),
.B(n_339),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_327),
.A2(n_325),
.B1(n_321),
.B2(n_322),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_306),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_331),
.A2(n_316),
.B(n_309),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_308),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_338),
.B(n_330),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_340),
.A2(n_332),
.B(n_335),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_342),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_343),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_345),
.B(n_343),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_348),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_344),
.C(n_346),
.Y(n_350)
);

AOI321xp33_ASAP7_75t_SL g351 ( 
.A1(n_350),
.A2(n_341),
.A3(n_347),
.B1(n_336),
.B2(n_292),
.C(n_296),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_275),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_352),
.Y(n_353)
);


endmodule