module fake_jpeg_4834_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_26),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_1),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_37),
.Y(n_48)
);

BUFx12f_ASAP7_75t_SL g36 ( 
.A(n_23),
.Y(n_36)
);

AND2x4_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx2_ASAP7_75t_SL g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_52),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_58),
.Y(n_61)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_40),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_56),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_35),
.B1(n_32),
.B2(n_21),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_52),
.C(n_20),
.Y(n_74)
);

CKINVDCx9p33_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_75),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_39),
.B(n_38),
.C(n_30),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_74),
.B(n_20),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_25),
.B1(n_21),
.B2(n_29),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_25),
.B1(n_21),
.B2(n_27),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_15),
.B1(n_27),
.B2(n_28),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_26),
.B1(n_28),
.B2(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_16),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_81),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_44),
.B1(n_59),
.B2(n_50),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_80),
.B1(n_49),
.B2(n_42),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_44),
.B1(n_59),
.B2(n_57),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_66),
.B1(n_22),
.B2(n_24),
.Y(n_103)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_48),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_38),
.B(n_39),
.C(n_46),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_91),
.B1(n_45),
.B2(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_16),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_92),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_61),
.Y(n_106)
);

AO21x1_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_41),
.B(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_16),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_96),
.B(n_106),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_76),
.Y(n_98)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_110),
.B(n_106),
.C(n_80),
.D(n_104),
.Y(n_128)
);

XNOR2x1_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_66),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_102),
.C(n_79),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_74),
.C(n_61),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_113),
.B1(n_82),
.B2(n_95),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_83),
.B1(n_84),
.B2(n_88),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_77),
.B(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_87),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_66),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_99),
.B(n_77),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_88),
.B1(n_66),
.B2(n_91),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_126),
.C(n_60),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_120),
.B(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_117),
.B(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_125),
.Y(n_137)
);

XNOR2x2_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_90),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_60),
.B1(n_16),
.B2(n_19),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_62),
.B1(n_16),
.B2(n_19),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_102),
.C(n_85),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_80),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_96),
.A2(n_97),
.B(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_82),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_81),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_91),
.B(n_68),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_91),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_133),
.B(n_135),
.CI(n_145),
.CON(n_158),
.SN(n_158)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_141),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_147),
.C(n_118),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_114),
.B1(n_117),
.B2(n_129),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_4),
.B(n_5),
.Y(n_159)
);

OAI322xp33_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_16),
.A3(n_81),
.B1(n_62),
.B2(n_56),
.C1(n_13),
.C2(n_14),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_122),
.Y(n_149)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

AOI221x1_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_19),
.B1(n_17),
.B2(n_56),
.C(n_13),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_56),
.B1(n_2),
.B2(n_3),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_146),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_12),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_126),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_150),
.C(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_152),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_116),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_124),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_154),
.A2(n_160),
.B1(n_152),
.B2(n_158),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_131),
.C(n_114),
.Y(n_156)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_134),
.B1(n_137),
.B2(n_133),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_5),
.C(n_6),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_12),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_135),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_162),
.B(n_150),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_155),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_153),
.A2(n_144),
.B1(n_140),
.B2(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_143),
.B1(n_7),
.B2(n_8),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_169),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_162),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_162),
.B1(n_163),
.B2(n_171),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_151),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_180),
.C(n_181),
.Y(n_182)
);

NAND2x1p5_ASAP7_75t_R g177 ( 
.A(n_167),
.B(n_158),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_181),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_148),
.C(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_186),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_173),
.B(n_169),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_183),
.B(n_187),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_179),
.B(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_177),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_165),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_175),
.B(n_166),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_182),
.C(n_176),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_175),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_184),
.Y(n_194)
);

NOR5xp2_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.C(n_196),
.D(n_197),
.E(n_193),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_180),
.C(n_166),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_6),
.C(n_7),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_199),
.B(n_6),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_191),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_10),
.Y(n_201)
);


endmodule