module fake_jpeg_21641_n_145 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_1),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_1),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_15),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_37),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_78),
.Y(n_84)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_77),
.Y(n_89)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_49),
.B1(n_66),
.B2(n_61),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_86),
.B(n_50),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_78),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_87),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_68),
.C(n_54),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_67),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_57),
.B1(n_56),
.B2(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_69),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_95),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_93),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_77),
.B(n_73),
.C(n_54),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_52),
.B(n_62),
.C(n_51),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_63),
.A3(n_55),
.B1(n_59),
.B2(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_101),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_99),
.B(n_102),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_48),
.Y(n_113)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_58),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_64),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_110),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_77),
.B1(n_71),
.B2(n_70),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_114),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_67),
.B1(n_2),
.B2(n_3),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_116),
.Y(n_126)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_23),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_47),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_123),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_26),
.A3(n_43),
.B1(n_42),
.B2(n_39),
.C1(n_38),
.C2(n_10),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_112),
.B(n_108),
.Y(n_129)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_124),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_125),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_131),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_107),
.B1(n_109),
.B2(n_6),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_119),
.B1(n_117),
.B2(n_126),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_24),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_134),
.B(n_135),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_122),
.B1(n_4),
.B2(n_7),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_133),
.C(n_132),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_128),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_127),
.B(n_30),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_27),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_16),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_32),
.B(n_36),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_14),
.B1(n_34),
.B2(n_33),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_11),
.C(n_44),
.Y(n_145)
);


endmodule