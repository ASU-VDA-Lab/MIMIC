module real_jpeg_19181_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_0),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_0),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_0),
.A2(n_51),
.B1(n_52),
.B2(n_72),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_1),
.A2(n_36),
.B1(n_51),
.B2(n_52),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_1),
.A2(n_36),
.B1(n_66),
.B2(n_67),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_2),
.A2(n_66),
.B1(n_67),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_2),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_3),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_3),
.A2(n_29),
.B1(n_51),
.B2(n_52),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_3),
.A2(n_29),
.B1(n_66),
.B2(n_67),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_4),
.A2(n_66),
.B1(n_67),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_4),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_6),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_6),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_7),
.A2(n_32),
.B(n_63),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_7),
.B(n_100),
.Y(n_139)
);

A2O1A1O1Ixp25_ASAP7_75t_L g152 ( 
.A1(n_7),
.A2(n_52),
.B(n_83),
.C(n_153),
.D(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_7),
.B(n_52),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_7),
.B(n_50),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_7),
.A2(n_69),
.B(n_168),
.Y(n_186)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_7),
.A2(n_31),
.B(n_45),
.C(n_54),
.D(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_7),
.B(n_31),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_43),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_8),
.A2(n_43),
.B1(n_66),
.B2(n_67),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_8),
.A2(n_43),
.B1(n_51),
.B2(n_52),
.Y(n_198)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_10),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_81),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_81),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_12),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_12),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_12),
.A2(n_51),
.B1(n_52),
.B2(n_68),
.Y(n_88)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_104),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_21),
.B(n_104),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_73),
.C(n_90),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_22),
.B(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_58),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_40),
.B1(n_41),
.B2(n_57),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_25),
.A2(n_30),
.B1(n_38),
.B2(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_30),
.B(n_33),
.C(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_33),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_27),
.A2(n_33),
.B(n_61),
.C(n_62),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_46),
.B(n_49),
.C(n_50),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_46),
.Y(n_49)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_35),
.B(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_37),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_40),
.B(n_57),
.C(n_58),
.Y(n_125)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B(n_53),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_42),
.A2(n_44),
.B1(n_56),
.B2(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_45),
.B(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_46),
.B(n_52),
.Y(n_206)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_49),
.A2(n_51),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_84),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_56),
.A2(n_117),
.B(n_119),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_56),
.A2(n_103),
.B(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_59),
.A2(n_60),
.B1(n_64),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_61),
.B(n_89),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_61),
.B(n_143),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_64),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_65),
.A2(n_69),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_67),
.B1(n_84),
.B2(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_66),
.B(n_84),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_66),
.B(n_188),
.Y(n_187)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_67),
.A2(n_85),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_71),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_69),
.A2(n_75),
.B1(n_77),
.B2(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_69),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_69),
.Y(n_175)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_70),
.A2(n_174),
.B(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_73),
.B(n_90),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_79),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_75),
.A2(n_142),
.B(n_183),
.Y(n_207)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_88),
.B2(n_89),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_89),
.B(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_88),
.B1(n_89),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_82),
.A2(n_89),
.B1(n_165),
.B2(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_82),
.A2(n_198),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_94),
.Y(n_93)
);

CKINVDCx9p33_ASAP7_75t_R g87 ( 
.A(n_84),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_89),
.B(n_95),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_89),
.A2(n_93),
.B(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.C(n_101),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_91),
.A2(n_92),
.B1(n_101),
.B2(n_102),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_125),
.B2(n_126),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_113),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_116),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_125),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_146),
.B(n_230),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_144),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_130),
.B(n_144),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_135),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_131),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_133),
.A2(n_135),
.B1(n_136),
.B2(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_133),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.C(n_140),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_137),
.A2(n_138),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_139),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_224),
.B(n_229),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_210),
.B(n_223),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_192),
.B(n_209),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_170),
.B(n_191),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_159),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_151),
.B(n_159),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_152),
.A2(n_155),
.B1(n_156),
.B2(n_179),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_153),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_164),
.C(n_166),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_167),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_169),
.B(n_175),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_180),
.B(n_190),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_178),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_172),
.B(n_178),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_185),
.B(n_189),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_184),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_193),
.B(n_194),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_203),
.B2(n_208),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_197),
.Y(n_202)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_202),
.C(n_208),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_200),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_203),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_207),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_211),
.B(n_212),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_219),
.C(n_221),
.Y(n_225)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_218),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_219),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_225),
.B(n_226),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);


endmodule