module real_aes_2812_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_792;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_815;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g540 ( .A(n_0), .B(n_178), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_1), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g144 ( .A(n_2), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_3), .B(n_543), .Y(n_562) );
NAND2xp33_ASAP7_75t_SL g533 ( .A(n_4), .B(n_156), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_5), .B(n_163), .Y(n_169) );
INVx1_ASAP7_75t_L g525 ( .A(n_6), .Y(n_525) );
INVx1_ASAP7_75t_L g209 ( .A(n_7), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_8), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_9), .Y(n_248) );
AND2x2_ASAP7_75t_L g560 ( .A(n_10), .B(n_186), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_11), .A2(n_807), .B1(n_814), .B2(n_816), .Y(n_813) );
INVx2_ASAP7_75t_L g133 ( .A(n_12), .Y(n_133) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_13), .Y(n_115) );
INVx1_ASAP7_75t_L g179 ( .A(n_14), .Y(n_179) );
AOI221x1_ASAP7_75t_L g528 ( .A1(n_15), .A2(n_130), .B1(n_529), .B2(n_531), .C(n_532), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_16), .B(n_543), .Y(n_596) );
INVx1_ASAP7_75t_L g119 ( .A(n_17), .Y(n_119) );
INVx1_ASAP7_75t_L g176 ( .A(n_18), .Y(n_176) );
INVx1_ASAP7_75t_SL g191 ( .A(n_19), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_20), .B(n_150), .Y(n_276) );
AOI33xp33_ASAP7_75t_L g221 ( .A1(n_21), .A2(n_48), .A3(n_139), .B1(n_148), .B2(n_222), .B3(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_22), .A2(n_531), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_23), .B(n_178), .Y(n_565) );
AOI221xp5_ASAP7_75t_SL g605 ( .A1(n_24), .A2(n_39), .B1(n_531), .B2(n_543), .C(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g242 ( .A(n_25), .Y(n_242) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_26), .A2(n_90), .B(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g164 ( .A(n_26), .B(n_90), .Y(n_164) );
INVxp67_ASAP7_75t_L g527 ( .A(n_27), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_28), .B(n_181), .Y(n_600) );
AND2x2_ASAP7_75t_L g554 ( .A(n_29), .B(n_185), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_30), .B(n_158), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_31), .A2(n_531), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_32), .B(n_181), .Y(n_607) );
INVx1_ASAP7_75t_L g138 ( .A(n_33), .Y(n_138) );
AND2x2_ASAP7_75t_L g156 ( .A(n_33), .B(n_144), .Y(n_156) );
AND2x2_ASAP7_75t_L g162 ( .A(n_33), .B(n_141), .Y(n_162) );
OR2x6_ASAP7_75t_L g117 ( .A(n_34), .B(n_118), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_35), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_36), .B(n_158), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_37), .A2(n_131), .B1(n_163), .B2(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_38), .B(n_278), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_40), .A2(n_82), .B1(n_136), .B2(n_531), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_41), .B(n_150), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_42), .B(n_178), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_43), .B(n_206), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_44), .B(n_150), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_45), .Y(n_273) );
AND2x2_ASAP7_75t_L g544 ( .A(n_46), .B(n_185), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_47), .B(n_185), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_49), .B(n_150), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_50), .A2(n_62), .B1(n_484), .B2(n_485), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_50), .Y(n_485) );
INVx1_ASAP7_75t_L g143 ( .A(n_51), .Y(n_143) );
INVx1_ASAP7_75t_L g152 ( .A(n_51), .Y(n_152) );
AOI22x1_ASAP7_75t_L g807 ( .A1(n_52), .A2(n_808), .B1(n_809), .B2(n_810), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_52), .Y(n_808) );
AND2x2_ASAP7_75t_L g235 ( .A(n_53), .B(n_185), .Y(n_235) );
AOI221xp5_ASAP7_75t_L g207 ( .A1(n_54), .A2(n_75), .B1(n_136), .B2(n_158), .C(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_55), .B(n_158), .Y(n_157) );
AOI222xp33_ASAP7_75t_R g103 ( .A1(n_56), .A2(n_104), .B1(n_109), .B2(n_495), .C1(n_500), .C2(n_818), .Y(n_103) );
OAI21xp5_ASAP7_75t_L g109 ( .A1(n_56), .A2(n_110), .B(n_487), .Y(n_109) );
INVx1_ASAP7_75t_L g490 ( .A(n_56), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_57), .B(n_543), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_58), .B(n_131), .Y(n_250) );
AOI21xp5_ASAP7_75t_SL g135 ( .A1(n_59), .A2(n_136), .B(n_145), .Y(n_135) );
AND2x2_ASAP7_75t_L g581 ( .A(n_60), .B(n_185), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_61), .B(n_181), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_62), .Y(n_484) );
INVx1_ASAP7_75t_L g172 ( .A(n_63), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_64), .B(n_178), .Y(n_579) );
AND2x2_ASAP7_75t_SL g601 ( .A(n_65), .B(n_186), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_66), .A2(n_531), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g233 ( .A(n_67), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_68), .B(n_181), .Y(n_566) );
AND2x2_ASAP7_75t_SL g573 ( .A(n_69), .B(n_206), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_70), .A2(n_102), .B1(n_811), .B2(n_812), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_70), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_71), .A2(n_136), .B(n_232), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_72), .A2(n_482), .B1(n_483), .B2(n_486), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_72), .Y(n_482) );
INVx1_ASAP7_75t_L g141 ( .A(n_73), .Y(n_141) );
INVx1_ASAP7_75t_L g154 ( .A(n_73), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_74), .B(n_158), .Y(n_224) );
AND2x2_ASAP7_75t_L g193 ( .A(n_76), .B(n_130), .Y(n_193) );
INVx1_ASAP7_75t_L g173 ( .A(n_77), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_78), .A2(n_136), .B(n_190), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_79), .A2(n_136), .B(n_216), .C(n_275), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_80), .A2(n_85), .B1(n_158), .B2(n_543), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_81), .B(n_543), .Y(n_580) );
INVx1_ASAP7_75t_L g120 ( .A(n_83), .Y(n_120) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_84), .B(n_130), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_86), .A2(n_136), .B1(n_219), .B2(n_220), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_87), .B(n_178), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_88), .B(n_178), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_89), .A2(n_531), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g146 ( .A(n_91), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_92), .B(n_181), .Y(n_578) );
AND2x2_ASAP7_75t_L g225 ( .A(n_93), .B(n_130), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_94), .A2(n_240), .B(n_241), .C(n_243), .Y(n_239) );
INVxp67_ASAP7_75t_L g530 ( .A(n_95), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_96), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_97), .B(n_181), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_98), .A2(n_531), .B(n_598), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_99), .Y(n_494) );
BUFx2_ASAP7_75t_L g108 ( .A(n_100), .Y(n_108) );
BUFx2_ASAP7_75t_SL g822 ( .A(n_100), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_101), .B(n_150), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_102), .Y(n_812) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_SL g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx2_ASAP7_75t_L g498 ( .A(n_106), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_106), .A2(n_820), .B(n_823), .Y(n_819) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_108), .B(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_121), .Y(n_110) );
CKINVDCx11_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g492 ( .A(n_114), .Y(n_492) );
BUFx2_ASAP7_75t_L g499 ( .A(n_114), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x6_ASAP7_75t_SL g515 ( .A(n_115), .B(n_117), .Y(n_515) );
OR2x6_ASAP7_75t_SL g806 ( .A(n_115), .B(n_116), .Y(n_806) );
OR2x2_ASAP7_75t_L g817 ( .A(n_115), .B(n_117), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_121), .Y(n_488) );
XNOR2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_480), .Y(n_121) );
NAND3x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_367), .C(n_444), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_319), .Y(n_123) );
NAND5xp2_ASAP7_75t_L g505 ( .A(n_124), .B(n_319), .C(n_506), .D(n_507), .E(n_508), .Y(n_505) );
INVxp33_ASAP7_75t_L g512 ( .A(n_124), .Y(n_512) );
NOR2xp67_ASAP7_75t_L g124 ( .A(n_125), .B(n_259), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_194), .B1(n_201), .B2(n_252), .Y(n_125) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_165), .Y(n_126) );
NOR2xp67_ASAP7_75t_SL g302 ( .A(n_127), .B(n_303), .Y(n_302) );
AND2x4_ASAP7_75t_L g317 ( .A(n_127), .B(n_318), .Y(n_317) );
NOR2x1_ASAP7_75t_L g334 ( .A(n_127), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_SL g374 ( .A(n_127), .B(n_375), .Y(n_374) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_128), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_128), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g309 ( .A(n_128), .Y(n_309) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_128), .Y(n_314) );
AND2x2_ASAP7_75t_L g343 ( .A(n_128), .B(n_283), .Y(n_343) );
OR2x2_ASAP7_75t_L g347 ( .A(n_128), .B(n_183), .Y(n_347) );
AND2x4_ASAP7_75t_L g360 ( .A(n_128), .B(n_318), .Y(n_360) );
NOR2x1_ASAP7_75t_SL g362 ( .A(n_128), .B(n_168), .Y(n_362) );
AND2x2_ASAP7_75t_L g390 ( .A(n_128), .B(n_268), .Y(n_390) );
OR2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_134), .Y(n_128) );
INVx3_ASAP7_75t_L g228 ( .A(n_130), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_130), .A2(n_228), .B1(n_239), .B2(n_244), .Y(n_238) );
INVx4_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_131), .B(n_247), .Y(n_246) );
AOI21x1_ASAP7_75t_L g536 ( .A1(n_131), .A2(n_537), .B(n_544), .Y(n_536) );
INVx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx4f_ASAP7_75t_L g206 ( .A(n_132), .Y(n_206) );
AND2x4_ASAP7_75t_L g163 ( .A(n_133), .B(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_SL g186 ( .A(n_133), .B(n_164), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_157), .B(n_163), .Y(n_134) );
INVxp67_ASAP7_75t_L g249 ( .A(n_136), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_136), .A2(n_158), .B1(n_524), .B2(n_526), .Y(n_523) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_142), .Y(n_136) );
NOR2x1p5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
INVx1_ASAP7_75t_L g223 ( .A(n_139), .Y(n_223) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x6_ASAP7_75t_L g147 ( .A(n_140), .B(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x6_ASAP7_75t_L g178 ( .A(n_141), .B(n_151), .Y(n_178) );
AND2x6_ASAP7_75t_L g531 ( .A(n_142), .B(n_162), .Y(n_531) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
INVx2_ASAP7_75t_L g148 ( .A(n_143), .Y(n_148) );
AND2x4_ASAP7_75t_L g181 ( .A(n_143), .B(n_153), .Y(n_181) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_144), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_149), .C(n_155), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_147), .A2(n_172), .B1(n_173), .B2(n_174), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g190 ( .A1(n_147), .A2(n_155), .B(n_191), .C(n_192), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_SL g208 ( .A1(n_147), .A2(n_155), .B(n_209), .C(n_210), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_147), .A2(n_155), .B(n_233), .C(n_234), .Y(n_232) );
INVxp67_ASAP7_75t_L g240 ( .A(n_147), .Y(n_240) );
INVx2_ASAP7_75t_L g278 ( .A(n_147), .Y(n_278) );
AND2x2_ASAP7_75t_L g159 ( .A(n_148), .B(n_160), .Y(n_159) );
INVxp33_ASAP7_75t_L g222 ( .A(n_148), .Y(n_222) );
INVx1_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
AND2x4_ASAP7_75t_L g543 ( .A(n_150), .B(n_156), .Y(n_543) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_155), .B(n_163), .Y(n_182) );
INVx1_ASAP7_75t_L g219 ( .A(n_155), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_155), .A2(n_276), .B(n_277), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_155), .A2(n_540), .B(n_541), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_155), .A2(n_551), .B(n_552), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_155), .A2(n_565), .B(n_566), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_155), .A2(n_578), .B(n_579), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_155), .A2(n_599), .B(n_600), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_155), .A2(n_607), .B(n_608), .Y(n_606) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_156), .Y(n_243) );
INVx1_ASAP7_75t_L g251 ( .A(n_158), .Y(n_251) );
AND2x4_ASAP7_75t_L g158 ( .A(n_159), .B(n_161), .Y(n_158) );
INVx1_ASAP7_75t_L g271 ( .A(n_159), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_161), .Y(n_272) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_163), .B(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_163), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_163), .B(n_530), .Y(n_529) );
NOR3xp33_ASAP7_75t_L g532 ( .A(n_163), .B(n_174), .C(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_163), .A2(n_562), .B(n_563), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_165), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_166), .A2(n_448), .B1(n_450), .B2(n_453), .Y(n_447) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_183), .Y(n_166) );
INVx1_ASAP7_75t_L g200 ( .A(n_167), .Y(n_200) );
AND2x2_ASAP7_75t_L g305 ( .A(n_167), .B(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g310 ( .A(n_167), .B(n_268), .Y(n_310) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g267 ( .A(n_168), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g283 ( .A(n_168), .Y(n_283) );
AND2x2_ASAP7_75t_L g316 ( .A(n_168), .B(n_183), .Y(n_316) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_175), .B(n_182), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_174), .B(n_242), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B1(n_179), .B2(n_180), .Y(n_175) );
INVxp67_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVxp67_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g198 ( .A(n_183), .Y(n_198) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_183), .Y(n_285) );
INVx1_ASAP7_75t_L g304 ( .A(n_183), .Y(n_304) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_183), .Y(n_373) );
INVx1_ASAP7_75t_L g385 ( .A(n_183), .Y(n_385) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_187), .B(n_193), .Y(n_183) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_184), .A2(n_548), .B(n_554), .Y(n_547) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_184), .A2(n_575), .B(n_581), .Y(n_574) );
AO21x2_ASAP7_75t_L g612 ( .A1(n_184), .A2(n_548), .B(n_554), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
OA21x2_ASAP7_75t_L g604 ( .A1(n_185), .A2(n_605), .B(n_609), .Y(n_604) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OAI31xp33_ASAP7_75t_SL g439 ( .A1(n_195), .A2(n_440), .A3(n_441), .B(n_442), .Y(n_439) );
NOR2x1_ASAP7_75t_L g195 ( .A(n_196), .B(n_199), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g364 ( .A(n_197), .B(n_266), .Y(n_364) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g280 ( .A(n_198), .Y(n_280) );
AND2x4_ASAP7_75t_SL g400 ( .A(n_200), .B(n_304), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_201), .A2(n_321), .B(n_324), .Y(n_320) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_212), .Y(n_201) );
INVx2_ASAP7_75t_L g293 ( .A(n_202), .Y(n_293) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2x1p5_ASAP7_75t_L g420 ( .A(n_203), .B(n_328), .Y(n_420) );
BUFx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g330 ( .A(n_204), .B(n_236), .Y(n_330) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVxp67_ASAP7_75t_L g255 ( .A(n_205), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_205), .B(n_215), .Y(n_290) );
AND2x4_ASAP7_75t_L g300 ( .A(n_205), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g345 ( .A(n_205), .B(n_237), .Y(n_345) );
INVx2_ASAP7_75t_L g353 ( .A(n_205), .Y(n_353) );
INVx1_ASAP7_75t_L g452 ( .A(n_205), .Y(n_452) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_205), .Y(n_461) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_211), .Y(n_205) );
INVx2_ASAP7_75t_SL g216 ( .A(n_206), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_206), .A2(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g398 ( .A(n_212), .Y(n_398) );
NAND2x1p5_ASAP7_75t_L g212 ( .A(n_213), .B(n_226), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g254 ( .A(n_214), .B(n_255), .Y(n_254) );
AND2x4_ASAP7_75t_L g393 ( .A(n_214), .B(n_328), .Y(n_393) );
AND2x2_ASAP7_75t_L g410 ( .A(n_214), .B(n_227), .Y(n_410) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_215), .B(n_258), .Y(n_433) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_225), .Y(n_215) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_216), .A2(n_217), .B(n_225), .Y(n_263) );
AOI21x1_ASAP7_75t_L g569 ( .A1(n_216), .A2(n_570), .B(n_573), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_218), .B(n_224), .Y(n_217) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g356 ( .A(n_226), .B(n_254), .Y(n_356) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_236), .Y(n_226) );
INVx2_ASAP7_75t_L g262 ( .A(n_227), .Y(n_262) );
NOR2xp67_ASAP7_75t_L g443 ( .A(n_227), .B(n_236), .Y(n_443) );
NOR2x1_ASAP7_75t_L g451 ( .A(n_227), .B(n_452), .Y(n_451) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_235), .Y(n_227) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_228), .A2(n_229), .B(n_235), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AND2x2_ASAP7_75t_L g359 ( .A(n_236), .B(n_263), .Y(n_359) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_237), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g288 ( .A(n_237), .Y(n_288) );
AND2x4_ASAP7_75t_L g352 ( .A(n_237), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g382 ( .A(n_237), .Y(n_382) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_245), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_249), .B1(n_250), .B2(n_251), .Y(n_245) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OAI221xp5_ASAP7_75t_L g403 ( .A1(n_253), .A2(n_266), .B1(n_404), .B2(n_405), .C(n_406), .Y(n_403) );
NAND2x1p5_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
AND2x2_ASAP7_75t_L g380 ( .A(n_254), .B(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_L g423 ( .A(n_254), .Y(n_423) );
INVx2_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g366 ( .A(n_257), .B(n_290), .Y(n_366) );
INVx3_ASAP7_75t_L g328 ( .A(n_258), .Y(n_328) );
AND2x2_ASAP7_75t_L g460 ( .A(n_258), .B(n_461), .Y(n_460) );
NAND3xp33_ASAP7_75t_SL g259 ( .A(n_260), .B(n_291), .C(n_307), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_264), .B1(n_281), .B2(n_286), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_261), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g391 ( .A(n_261), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g402 ( .A(n_261), .B(n_297), .Y(n_402) );
AND2x2_ASAP7_75t_L g472 ( .A(n_261), .B(n_345), .Y(n_472) );
AND2x4_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g301 ( .A(n_263), .Y(n_301) );
INVx1_ASAP7_75t_L g350 ( .A(n_263), .Y(n_350) );
INVxp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OAI222xp33_ASAP7_75t_L g417 ( .A1(n_265), .A2(n_418), .B1(n_419), .B2(n_421), .C1(n_422), .C2(n_424), .Y(n_417) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_279), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_266), .B(n_293), .Y(n_292) );
NOR2x1_ASAP7_75t_L g425 ( .A(n_266), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g384 ( .A(n_267), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g440 ( .A(n_267), .B(n_314), .Y(n_440) );
INVx2_ASAP7_75t_L g306 ( .A(n_268), .Y(n_306) );
INVx1_ASAP7_75t_L g318 ( .A(n_268), .Y(n_318) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_268), .Y(n_375) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_274), .Y(n_268) );
NOR3xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .C(n_273), .Y(n_270) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_280), .Y(n_323) );
INVx3_ASAP7_75t_L g342 ( .A(n_280), .Y(n_342) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g408 ( .A(n_282), .Y(n_408) );
NAND2x1_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g395 ( .A(n_284), .Y(n_395) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g396 ( .A(n_287), .Y(n_396) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g297 ( .A(n_288), .Y(n_297) );
AND2x2_ASAP7_75t_L g415 ( .A(n_288), .B(n_300), .Y(n_415) );
AND2x2_ASAP7_75t_L g478 ( .A(n_288), .B(n_410), .Y(n_478) );
AND2x2_ASAP7_75t_L g407 ( .A(n_289), .B(n_327), .Y(n_407) );
INVx1_ASAP7_75t_L g418 ( .A(n_289), .Y(n_418) );
AND2x2_ASAP7_75t_L g435 ( .A(n_289), .B(n_382), .Y(n_435) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_294), .B1(n_298), .B2(n_302), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_294), .A2(n_308), .B(n_311), .Y(n_307) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g339 ( .A(n_297), .B(n_300), .Y(n_339) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g442 ( .A(n_300), .B(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g405 ( .A(n_303), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_304), .Y(n_333) );
AND2x2_ASAP7_75t_SL g313 ( .A(n_305), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g378 ( .A(n_305), .Y(n_378) );
AND2x2_ASAP7_75t_L g476 ( .A(n_305), .B(n_373), .Y(n_476) );
INVx1_ASAP7_75t_L g431 ( .A(n_306), .Y(n_431) );
INVx1_ASAP7_75t_L g337 ( .A(n_308), .Y(n_337) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g426 ( .A(n_309), .Y(n_426) );
INVx4_ASAP7_75t_L g335 ( .A(n_310), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI32xp33_ASAP7_75t_L g406 ( .A1(n_313), .A2(n_407), .A3(n_408), .B1(n_409), .B2(n_410), .Y(n_406) );
AND2x2_ASAP7_75t_L g401 ( .A(n_314), .B(n_316), .Y(n_401) );
O2A1O1Ixp33_ASAP7_75t_SL g464 ( .A1(n_314), .A2(n_465), .B(n_466), .C(n_468), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_SL g429 ( .A(n_316), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g468 ( .A(n_316), .Y(n_468) );
AND2x2_ASAP7_75t_L g322 ( .A(n_317), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g449 ( .A(n_317), .Y(n_449) );
AND2x2_ASAP7_75t_L g455 ( .A(n_317), .B(n_342), .Y(n_455) );
INVxp33_ASAP7_75t_SL g513 ( .A(n_319), .Y(n_513) );
NOR3x1_ASAP7_75t_L g319 ( .A(n_320), .B(n_336), .C(n_354), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_331), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
AND2x2_ASAP7_75t_L g344 ( .A(n_327), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g387 ( .A(n_327), .B(n_352), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_327), .B(n_373), .Y(n_414) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_335), .B(n_342), .Y(n_441) );
INVx2_ASAP7_75t_L g463 ( .A(n_335), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B(n_340), .Y(n_336) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_337), .A2(n_428), .B1(n_432), .B2(n_434), .C(n_439), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_338), .A2(n_458), .B1(n_459), .B2(n_462), .Y(n_457) );
INVx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B1(n_346), .B2(n_348), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
AND2x2_ASAP7_75t_L g386 ( .A(n_342), .B(n_362), .Y(n_386) );
INVx1_ASAP7_75t_L g392 ( .A(n_342), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_342), .B(n_360), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_345), .B(n_413), .Y(n_479) );
NAND2x1_ASAP7_75t_L g462 ( .A(n_346), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_347), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
NAND2x1_ASAP7_75t_SL g465 ( .A(n_350), .B(n_352), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_350), .B(n_450), .Y(n_471) );
OR2x2_ASAP7_75t_L g432 ( .A(n_351), .B(n_433), .Y(n_432) );
INVx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g467 ( .A(n_352), .B(n_393), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_355), .B(n_361), .Y(n_354) );
OAI21xp33_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_357), .B(n_360), .Y(n_355) );
OR2x2_ASAP7_75t_L g419 ( .A(n_358), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g453 ( .A(n_359), .B(n_451), .Y(n_453) );
AND2x2_ASAP7_75t_SL g399 ( .A(n_360), .B(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g409 ( .A(n_360), .Y(n_409) );
OAI21xp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_363), .B(n_365), .Y(n_361) );
AND2x2_ASAP7_75t_L g394 ( .A(n_362), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g506 ( .A(n_368), .Y(n_506) );
OAI21xp33_ASAP7_75t_L g510 ( .A1(n_368), .A2(n_445), .B(n_485), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_411), .Y(n_368) );
NOR3xp33_ASAP7_75t_SL g369 ( .A(n_370), .B(n_388), .C(n_403), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_376), .B(n_379), .C(n_383), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g437 ( .A(n_382), .Y(n_437) );
AND2x2_ASAP7_75t_L g450 ( .A(n_382), .B(n_451), .Y(n_450) );
OAI21xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .B(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g458 ( .A(n_384), .Y(n_458) );
OAI21xp5_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_396), .B(n_397), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_393), .B2(n_394), .Y(n_389) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_390), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_401), .B2(n_402), .Y(n_397) );
INVx1_ASAP7_75t_SL g404 ( .A(n_402), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_408), .B(n_449), .Y(n_448) );
OAI22xp33_ASAP7_75t_SL g474 ( .A1(n_409), .A2(n_475), .B1(n_477), .B2(n_479), .Y(n_474) );
AOI211x1_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_416), .B(n_417), .C(n_427), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_429), .A2(n_470), .B(n_472), .Y(n_469) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g438 ( .A(n_433), .Y(n_438) );
NOR2xp67_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_436), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND4xp25_ASAP7_75t_L g445 ( .A(n_446), .B(n_456), .C(n_469), .D(n_473), .Y(n_445) );
AND2x2_ASAP7_75t_L g507 ( .A(n_446), .B(n_456), .Y(n_507) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_454), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_464), .Y(n_456) );
INVxp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVxp67_ASAP7_75t_L g509 ( .A(n_469), .Y(n_509) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g508 ( .A(n_474), .B(n_485), .C(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g486 ( .A(n_483), .Y(n_486) );
OAI21xp33_ASAP7_75t_L g511 ( .A1(n_485), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B(n_493), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_492), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g823 ( .A(n_492), .Y(n_823) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_499), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_807), .B(n_813), .Y(n_500) );
INVxp67_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OAI22x1_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_514), .B1(n_516), .B2(n_804), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_504), .A2(n_514), .B1(n_517), .B2(n_815), .Y(n_814) );
AND3x1_ASAP7_75t_L g504 ( .A(n_505), .B(n_510), .C(n_511), .Y(n_504) );
CKINVDCx11_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_518), .B(n_681), .Y(n_517) );
NOR4xp25_ASAP7_75t_L g518 ( .A(n_519), .B(n_624), .C(n_663), .D(n_670), .Y(n_518) );
OAI221xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_545), .B1(n_582), .B2(n_591), .C(n_610), .Y(n_519) );
OR2x2_ASAP7_75t_L g754 ( .A(n_520), .B(n_616), .Y(n_754) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g669 ( .A(n_521), .B(n_594), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_521), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_SL g734 ( .A(n_521), .B(n_735), .Y(n_734) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_534), .Y(n_521) );
AND2x4_ASAP7_75t_SL g593 ( .A(n_522), .B(n_594), .Y(n_593) );
INVx3_ASAP7_75t_L g615 ( .A(n_522), .Y(n_615) );
AND2x2_ASAP7_75t_L g650 ( .A(n_522), .B(n_623), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_522), .B(n_535), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_522), .B(n_617), .Y(n_702) );
OR2x2_ASAP7_75t_L g780 ( .A(n_522), .B(n_594), .Y(n_780) );
AND2x4_ASAP7_75t_L g522 ( .A(n_523), .B(n_528), .Y(n_522) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g602 ( .A(n_535), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_535), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g628 ( .A(n_535), .Y(n_628) );
OR2x2_ASAP7_75t_L g633 ( .A(n_535), .B(n_617), .Y(n_633) );
AND2x2_ASAP7_75t_L g646 ( .A(n_535), .B(n_604), .Y(n_646) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_535), .Y(n_649) );
INVx1_ASAP7_75t_L g661 ( .A(n_535), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_535), .B(n_615), .Y(n_726) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_546), .B(n_555), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g590 ( .A(n_547), .B(n_574), .Y(n_590) );
AND2x4_ASAP7_75t_L g620 ( .A(n_547), .B(n_559), .Y(n_620) );
INVx2_ASAP7_75t_L g654 ( .A(n_547), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_547), .B(n_574), .Y(n_712) );
AND2x2_ASAP7_75t_L g759 ( .A(n_547), .B(n_588), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_553), .Y(n_548) );
AOI222xp33_ASAP7_75t_L g747 ( .A1(n_555), .A2(n_619), .B1(n_662), .B2(n_722), .C1(n_748), .C2(n_750), .Y(n_747) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_567), .Y(n_556) );
AND2x2_ASAP7_75t_L g666 ( .A(n_557), .B(n_586), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_557), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g795 ( .A(n_557), .B(n_635), .Y(n_795) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_558), .A2(n_626), .B(n_630), .Y(n_625) );
AND2x2_ASAP7_75t_L g706 ( .A(n_558), .B(n_589), .Y(n_706) );
OR2x2_ASAP7_75t_L g731 ( .A(n_558), .B(n_590), .Y(n_731) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx5_ASAP7_75t_L g585 ( .A(n_559), .Y(n_585) );
AND2x2_ASAP7_75t_L g672 ( .A(n_559), .B(n_654), .Y(n_672) );
AND2x2_ASAP7_75t_L g698 ( .A(n_559), .B(n_574), .Y(n_698) );
OR2x2_ASAP7_75t_L g701 ( .A(n_559), .B(n_588), .Y(n_701) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_559), .Y(n_719) );
AND2x4_ASAP7_75t_SL g776 ( .A(n_559), .B(n_653), .Y(n_776) );
OR2x2_ASAP7_75t_L g785 ( .A(n_559), .B(n_612), .Y(n_785) );
OR2x6_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g618 ( .A(n_567), .Y(n_618) );
AOI221xp5_ASAP7_75t_SL g736 ( .A1(n_567), .A2(n_620), .B1(n_737), .B2(n_739), .C(n_740), .Y(n_736) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_574), .Y(n_567) );
OR2x2_ASAP7_75t_L g675 ( .A(n_568), .B(n_645), .Y(n_675) );
OR2x2_ASAP7_75t_L g685 ( .A(n_568), .B(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g711 ( .A(n_568), .B(n_712), .Y(n_711) );
AND2x4_ASAP7_75t_L g717 ( .A(n_568), .B(n_636), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_568), .B(n_700), .Y(n_729) );
INVx2_ASAP7_75t_L g742 ( .A(n_568), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g763 ( .A(n_568), .B(n_620), .Y(n_763) );
AND2x2_ASAP7_75t_L g767 ( .A(n_568), .B(n_589), .Y(n_767) );
AND2x2_ASAP7_75t_L g775 ( .A(n_568), .B(n_776), .Y(n_775) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g588 ( .A(n_569), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_574), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g619 ( .A(n_574), .B(n_588), .Y(n_619) );
INVx2_ASAP7_75t_L g636 ( .A(n_574), .Y(n_636) );
AND2x4_ASAP7_75t_L g653 ( .A(n_574), .B(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_574), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_580), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_586), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g765 ( .A(n_584), .B(n_587), .Y(n_765) );
AND2x4_ASAP7_75t_L g611 ( .A(n_585), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g652 ( .A(n_585), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g679 ( .A(n_585), .B(n_619), .Y(n_679) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
AND2x2_ASAP7_75t_L g783 ( .A(n_587), .B(n_784), .Y(n_783) );
BUFx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g635 ( .A(n_588), .B(n_636), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g655 ( .A1(n_589), .A2(n_656), .B(n_662), .Y(n_655) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_602), .Y(n_592) );
INVx1_ASAP7_75t_SL g709 ( .A(n_593), .Y(n_709) );
AND2x2_ASAP7_75t_L g739 ( .A(n_593), .B(n_649), .Y(n_739) );
AND2x4_ASAP7_75t_L g750 ( .A(n_593), .B(n_751), .Y(n_750) );
OR2x2_ASAP7_75t_L g616 ( .A(n_594), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g623 ( .A(n_594), .Y(n_623) );
AND2x4_ASAP7_75t_L g629 ( .A(n_594), .B(n_615), .Y(n_629) );
INVx2_ASAP7_75t_L g640 ( .A(n_594), .Y(n_640) );
INVx1_ASAP7_75t_L g689 ( .A(n_594), .Y(n_689) );
OR2x2_ASAP7_75t_L g710 ( .A(n_594), .B(n_694), .Y(n_710) );
OR2x2_ASAP7_75t_L g724 ( .A(n_594), .B(n_604), .Y(n_724) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_594), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_594), .B(n_646), .Y(n_796) );
OR2x6_ASAP7_75t_L g594 ( .A(n_595), .B(n_601), .Y(n_594) );
INVx1_ASAP7_75t_L g641 ( .A(n_602), .Y(n_641) );
AND2x2_ASAP7_75t_L g774 ( .A(n_602), .B(n_640), .Y(n_774) );
AND2x2_ASAP7_75t_L g799 ( .A(n_602), .B(n_629), .Y(n_799) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g617 ( .A(n_604), .Y(n_617) );
BUFx3_ASAP7_75t_L g659 ( .A(n_604), .Y(n_659) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_604), .Y(n_686) );
INVx1_ASAP7_75t_L g695 ( .A(n_604), .Y(n_695) );
AOI33xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .A3(n_618), .B1(n_619), .B2(n_620), .B3(n_621), .Y(n_610) );
AOI21x1_ASAP7_75t_SL g713 ( .A1(n_611), .A2(n_635), .B(n_697), .Y(n_713) );
INVx2_ASAP7_75t_L g743 ( .A(n_611), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_611), .B(n_742), .Y(n_749) );
AND2x2_ASAP7_75t_L g697 ( .A(n_612), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g660 ( .A(n_615), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g761 ( .A(n_616), .Y(n_761) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_617), .Y(n_751) );
OAI32xp33_ASAP7_75t_L g800 ( .A1(n_618), .A2(n_620), .A3(n_796), .B1(n_801), .B2(n_803), .Y(n_800) );
AND2x2_ASAP7_75t_L g718 ( .A(n_619), .B(n_719), .Y(n_718) );
INVx2_ASAP7_75t_SL g708 ( .A(n_620), .Y(n_708) );
AND2x2_ASAP7_75t_L g773 ( .A(n_620), .B(n_717), .Y(n_773) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_634), .B1(n_637), .B2(n_651), .C(n_655), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_628), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_629), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_629), .B(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_629), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g678 ( .A(n_633), .Y(n_678) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NOR3xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_642), .C(n_647), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
OAI22xp33_ASAP7_75t_L g740 ( .A1(n_639), .A2(n_701), .B1(n_741), .B2(n_744), .Y(n_740) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g644 ( .A(n_640), .Y(n_644) );
NOR2x1p5_ASAP7_75t_L g658 ( .A(n_640), .B(n_659), .Y(n_658) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_640), .Y(n_680) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI322xp33_ASAP7_75t_L g707 ( .A1(n_643), .A2(n_685), .A3(n_708), .B1(n_709), .B2(n_710), .C1(n_711), .C2(n_713), .Y(n_707) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g663 ( .A1(n_645), .A2(n_664), .B(n_665), .C(n_667), .Y(n_663) );
OR2x2_ASAP7_75t_L g755 ( .A(n_645), .B(n_709), .Y(n_755) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g662 ( .A(n_646), .B(n_650), .Y(n_662) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g668 ( .A(n_652), .B(n_669), .Y(n_668) );
INVx3_ASAP7_75t_SL g700 ( .A(n_653), .Y(n_700) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_657), .B(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
INVx1_ASAP7_75t_SL g704 ( .A(n_660), .Y(n_704) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_661), .Y(n_746) );
OR2x6_ASAP7_75t_SL g801 ( .A(n_664), .B(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI211xp5_ASAP7_75t_L g791 ( .A1(n_669), .A2(n_792), .B(n_793), .C(n_800), .Y(n_791) );
O2A1O1Ixp33_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_673), .B(n_676), .C(n_680), .Y(n_670) );
OAI211xp5_ASAP7_75t_SL g682 ( .A1(n_671), .A2(n_683), .B(n_690), .C(n_714), .Y(n_682) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVxp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NOR3xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_727), .C(n_771), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_687), .Y(n_683) );
INVx1_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_686), .Y(n_778) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g733 ( .A(n_689), .Y(n_733) );
NOR3xp33_ASAP7_75t_SL g690 ( .A(n_691), .B(n_703), .C(n_707), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_696), .B1(n_699), .B2(n_702), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g735 ( .A(n_695), .Y(n_735) );
INVxp67_ASAP7_75t_SL g802 ( .A(n_695), .Y(n_802) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_SL g788 ( .A(n_701), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
OR2x2_ASAP7_75t_L g738 ( .A(n_704), .B(n_724), .Y(n_738) );
OR2x2_ASAP7_75t_L g789 ( .A(n_704), .B(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g787 ( .A(n_712), .Y(n_787) );
OR2x2_ASAP7_75t_L g803 ( .A(n_712), .B(n_742), .Y(n_803) );
OAI21xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_718), .B(n_720), .Y(n_714) );
OAI31xp33_ASAP7_75t_L g728 ( .A1(n_715), .A2(n_729), .A3(n_730), .B(n_732), .Y(n_728) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
AND2x4_ASAP7_75t_L g760 ( .A(n_725), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND4xp25_ASAP7_75t_SL g727 ( .A(n_728), .B(n_736), .C(n_747), .D(n_752), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_735), .Y(n_770) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVxp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_756), .B1(n_760), .B2(n_762), .C(n_764), .Y(n_752) );
NAND2xp33_ASAP7_75t_SL g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g797 ( .A(n_756), .Y(n_797) );
AND2x2_ASAP7_75t_SL g756 ( .A(n_757), .B(n_759), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AOI21xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B(n_768), .Y(n_764) );
INVx1_ASAP7_75t_L g792 ( .A(n_766), .Y(n_792) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g771 ( .A(n_772), .B(n_791), .Y(n_771) );
AOI221xp5_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B1(n_775), .B2(n_777), .C(n_781), .Y(n_772) );
AND2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
INVx1_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
AOI21xp33_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_786), .B(n_789), .Y(n_781) );
INVxp33_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_796), .B1(n_797), .B2(n_798), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_805), .Y(n_815) );
CKINVDCx11_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_SL g818 ( .A(n_819), .Y(n_818) );
CKINVDCx11_ASAP7_75t_R g820 ( .A(n_821), .Y(n_820) );
CKINVDCx8_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
endmodule