module fake_ariane_1860_n_2032 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2032);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2032;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_26),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_123),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_64),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_87),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_40),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_46),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_104),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_134),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_34),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_53),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_158),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_4),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_89),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_27),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_180),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_178),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_96),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_77),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_95),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_156),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_148),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_63),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_41),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_126),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_65),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_32),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_203),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_54),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_187),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_53),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_117),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_155),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_122),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_35),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_35),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_41),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_74),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_144),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_173),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_7),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_154),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_188),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_143),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_1),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_145),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_196),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_185),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_136),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_140),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_171),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_110),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_40),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_202),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_183),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_159),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_83),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_132),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_55),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_149),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_0),
.Y(n_275)
);

BUFx2_ASAP7_75t_R g276 ( 
.A(n_38),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_3),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_139),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_84),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_114),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_166),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_10),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_75),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_38),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_43),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_113),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_102),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_71),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_65),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_137),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_194),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_25),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_42),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_11),
.Y(n_294)
);

BUFx8_ASAP7_75t_SL g295 ( 
.A(n_197),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_182),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_100),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_129),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_25),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_74),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_109),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_28),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_115),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_75),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_24),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_69),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_167),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_20),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_195),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_49),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_52),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_169),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_31),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_10),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_31),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_174),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_55),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_138),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_91),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_46),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_49),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_11),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_79),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_172),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_170),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_105),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_153),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_165),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_121),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_131),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_85),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_181),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_192),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_29),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_93),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_142),
.Y(n_336)
);

HB1xp67_ASAP7_75t_SL g337 ( 
.A(n_1),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_3),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_24),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_17),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_128),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_98),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_67),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_2),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_103),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_59),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_73),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_108),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_19),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_2),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_22),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_92),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_124),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_64),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_45),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_36),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_116),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_150),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_27),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_80),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_130),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_20),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_78),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_168),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_198),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_37),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_9),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_193),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_8),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_17),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_54),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_99),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_59),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_43),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_86),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_15),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_175),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_0),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_21),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_177),
.Y(n_380)
);

BUFx8_ASAP7_75t_SL g381 ( 
.A(n_23),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_101),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_72),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_82),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_90),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_14),
.Y(n_386)
);

BUFx10_ASAP7_75t_L g387 ( 
.A(n_118),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_111),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_12),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_28),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_76),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_47),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_119),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_58),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_12),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_30),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_157),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_107),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_51),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_62),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_14),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_48),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_60),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_152),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_61),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_19),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_69),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_48),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_26),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_163),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_120),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_47),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_235),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_248),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_250),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_381),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_210),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_248),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_248),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_248),
.B(n_4),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_223),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_295),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_248),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_248),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_248),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_248),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_258),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_226),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_346),
.Y(n_429)
);

NOR2xp67_ASAP7_75t_L g430 ( 
.A(n_315),
.B(n_5),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_281),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_212),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_300),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_412),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g435 ( 
.A(n_315),
.B(n_5),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_277),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_253),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_223),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_266),
.B(n_6),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_375),
.Y(n_440)
);

NOR2xp67_ASAP7_75t_L g441 ( 
.A(n_322),
.B(n_6),
.Y(n_441)
);

INVxp33_ASAP7_75t_SL g442 ( 
.A(n_356),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_277),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_401),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_243),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_247),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_277),
.B(n_227),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_290),
.B(n_7),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_277),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_207),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_277),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_277),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g453 ( 
.A(n_337),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_207),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_275),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_282),
.Y(n_456)
);

CKINVDCx14_ASAP7_75t_R g457 ( 
.A(n_268),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_351),
.B(n_8),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_277),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_322),
.B(n_9),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_277),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_284),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_283),
.Y(n_463)
);

INVx4_ASAP7_75t_R g464 ( 
.A(n_375),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_284),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_284),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_351),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_240),
.B(n_13),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_274),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_284),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_284),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_285),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_216),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_216),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_234),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_234),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_367),
.B(n_13),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_264),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_288),
.Y(n_479)
);

INVxp33_ASAP7_75t_L g480 ( 
.A(n_205),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_209),
.B(n_15),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_289),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_218),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_292),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_218),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_264),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_213),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_293),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_294),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_329),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_299),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_329),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_363),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_354),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_302),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_363),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_217),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_221),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_233),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_361),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_268),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_304),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_382),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_237),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_268),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_241),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_272),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_382),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_308),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_365),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_311),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_305),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_221),
.Y(n_513)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_224),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_314),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_365),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_365),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_317),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_310),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_387),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_313),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_320),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_321),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_334),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_343),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_369),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_338),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_211),
.B(n_16),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_339),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_340),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_386),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_387),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_391),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_400),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_366),
.Y(n_535)
);

NOR2xp67_ASAP7_75t_L g536 ( 
.A(n_224),
.B(n_16),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_373),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_406),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_510),
.B(n_387),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_499),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_499),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_421),
.B(n_214),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_462),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_432),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_445),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_458),
.B(n_219),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_446),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_450),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_414),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_504),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_457),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_504),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_506),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_506),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_454),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_417),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_462),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_507),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_465),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_507),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_438),
.B(n_220),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_414),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_418),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_428),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_418),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_431),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_469),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_419),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_465),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_466),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_419),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_423),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_500),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_429),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_422),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_519),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_521),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_466),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_423),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_525),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_458),
.B(n_297),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_437),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_440),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_447),
.B(n_231),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_472),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_525),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_434),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_455),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_503),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_470),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_470),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_456),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_482),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_463),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_479),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_424),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_467),
.B(n_238),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_471),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_471),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_484),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_424),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_488),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_489),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_526),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_494),
.B(n_276),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_425),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_510),
.B(n_204),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_425),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_491),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_503),
.B(n_245),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_517),
.B(n_204),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_426),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_495),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_426),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_526),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_485),
.B(n_514),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_502),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_533),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_509),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_511),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_533),
.Y(n_621)
);

CKINVDCx16_ASAP7_75t_R g622 ( 
.A(n_517),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_515),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_518),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_522),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_523),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_524),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_436),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_527),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_605),
.A2(n_505),
.B1(n_516),
.B2(n_501),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_581),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_574),
.Y(n_632)
);

BUFx10_ASAP7_75t_L g633 ( 
.A(n_616),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_540),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_583),
.B(n_508),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_606),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_581),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_575),
.Y(n_638)
);

BUFx6f_ASAP7_75t_SL g639 ( 
.A(n_581),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_581),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_581),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_597),
.B(n_453),
.Y(n_642)
);

BUFx8_ASAP7_75t_SL g643 ( 
.A(n_544),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_606),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_541),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_549),
.B(n_529),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_608),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_597),
.B(n_480),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_575),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_549),
.B(n_530),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_545),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_550),
.B(n_487),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_584),
.B(n_508),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_628),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_552),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_583),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_547),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_549),
.B(n_565),
.Y(n_658)
);

AND2x6_ASAP7_75t_L g659 ( 
.A(n_546),
.B(n_297),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_628),
.Y(n_660)
);

AND2x2_ASAP7_75t_SL g661 ( 
.A(n_622),
.B(n_448),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_574),
.B(n_444),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_589),
.B(n_497),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_628),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_553),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_554),
.B(n_512),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_628),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_582),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_608),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_558),
.Y(n_670)
);

INVx6_ASAP7_75t_L g671 ( 
.A(n_628),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_560),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_614),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_546),
.B(n_535),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_562),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_562),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_563),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_546),
.B(n_537),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_576),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_565),
.B(n_252),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_579),
.B(n_255),
.Y(n_681)
);

INVx5_ASAP7_75t_L g682 ( 
.A(n_581),
.Y(n_682)
);

OA22x2_ASAP7_75t_L g683 ( 
.A1(n_546),
.A2(n_433),
.B1(n_427),
.B2(n_413),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_579),
.B(n_262),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_563),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_577),
.Y(n_686)
);

INVx5_ASAP7_75t_L g687 ( 
.A(n_581),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_579),
.B(n_265),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_568),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_601),
.B(n_267),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_568),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_589),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_587),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_580),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_586),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_610),
.B(n_534),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_601),
.B(n_269),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_571),
.B(n_473),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_604),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_543),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_571),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_615),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_572),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_610),
.B(n_538),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_610),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_582),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_618),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_596),
.B(n_474),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_596),
.B(n_270),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_612),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_587),
.B(n_483),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_621),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_612),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_607),
.B(n_442),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_543),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_592),
.B(n_278),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_557),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_611),
.B(n_498),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_543),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_588),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_548),
.B(n_468),
.C(n_439),
.Y(n_721)
);

AO22x2_ASAP7_75t_L g722 ( 
.A1(n_539),
.A2(n_249),
.B1(n_344),
.B2(n_306),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_559),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_555),
.B(n_513),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_569),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_569),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_570),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_592),
.B(n_279),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_570),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_542),
.B(n_415),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_578),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_561),
.B(n_520),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_543),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_594),
.A2(n_481),
.B1(n_528),
.B2(n_536),
.Y(n_734)
);

AND2x6_ASAP7_75t_L g735 ( 
.A(n_610),
.B(n_297),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_594),
.B(n_287),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_543),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_567),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_588),
.B(n_538),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_578),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_590),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_590),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_591),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_551),
.B(n_531),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_595),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_595),
.B(n_396),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_591),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_598),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_598),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_600),
.B(n_238),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_598),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_620),
.B(n_532),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_551),
.B(n_475),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_585),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_L g755 ( 
.A(n_600),
.B(n_420),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_598),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_599),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_599),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_599),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_599),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_599),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_602),
.B(n_291),
.Y(n_762)
);

CKINVDCx11_ASAP7_75t_R g763 ( 
.A(n_593),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_602),
.B(n_475),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_603),
.Y(n_765)
);

NOR2x1p5_ASAP7_75t_L g766 ( 
.A(n_603),
.B(n_347),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_609),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_609),
.B(n_476),
.Y(n_768)
);

NOR2x1p5_ASAP7_75t_L g769 ( 
.A(n_613),
.B(n_347),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_613),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_617),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_617),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_619),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_556),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_619),
.B(n_476),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_623),
.B(n_478),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_623),
.Y(n_777)
);

INVx4_ASAP7_75t_SL g778 ( 
.A(n_624),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_653),
.B(n_624),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_701),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_722),
.A2(n_486),
.B1(n_490),
.B2(n_478),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_776),
.B(n_625),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_675),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_755),
.A2(n_477),
.B(n_443),
.C(n_449),
.Y(n_784)
);

NAND2x1_ASAP7_75t_L g785 ( 
.A(n_631),
.B(n_464),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_722),
.A2(n_490),
.B1(n_492),
.B2(n_486),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_755),
.A2(n_443),
.B(n_449),
.C(n_436),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_765),
.B(n_626),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_739),
.B(n_626),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_674),
.B(n_627),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_765),
.B(n_627),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_678),
.B(n_629),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_768),
.B(n_629),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_739),
.B(n_492),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_720),
.Y(n_795)
);

AND2x6_ASAP7_75t_SL g796 ( 
.A(n_752),
.B(n_416),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_722),
.A2(n_496),
.B1(n_493),
.B2(n_435),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_639),
.B(n_297),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_676),
.Y(n_799)
);

O2A1O1Ixp5_ASAP7_75t_L g800 ( 
.A1(n_680),
.A2(n_452),
.B(n_459),
.C(n_451),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_676),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_716),
.B(n_374),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_648),
.B(n_705),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_648),
.B(n_642),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_677),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_764),
.B(n_493),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_770),
.B(n_206),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_677),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_775),
.B(n_496),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_775),
.B(n_273),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_696),
.B(n_323),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_716),
.B(n_376),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_728),
.B(n_378),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_720),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_728),
.B(n_379),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_736),
.B(n_383),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_696),
.B(n_704),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_685),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_736),
.B(n_762),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_696),
.B(n_324),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_698),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_642),
.B(n_573),
.Y(n_822)
);

INVxp67_ASAP7_75t_SL g823 ( 
.A(n_704),
.Y(n_823)
);

AO22x1_ASAP7_75t_L g824 ( 
.A1(n_714),
.A2(n_573),
.B1(n_556),
.B2(n_566),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_762),
.B(n_389),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_704),
.B(n_336),
.Y(n_826)
);

AND3x1_ASAP7_75t_L g827 ( 
.A(n_721),
.B(n_772),
.C(n_771),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_732),
.B(n_342),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_693),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_772),
.B(n_208),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_663),
.B(n_215),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_658),
.A2(n_689),
.B(n_685),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_662),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_778),
.B(n_430),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_722),
.A2(n_441),
.B1(n_460),
.B2(n_355),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_663),
.B(n_222),
.Y(n_836)
);

OAI22xp33_ASAP7_75t_L g837 ( 
.A1(n_734),
.A2(n_405),
.B1(n_349),
.B2(n_371),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_643),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_730),
.B(n_564),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_652),
.B(n_225),
.Y(n_840)
);

INVx8_ASAP7_75t_L g841 ( 
.A(n_639),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_691),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_773),
.B(n_225),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_750),
.B(n_564),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_773),
.B(n_228),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_652),
.B(n_228),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_708),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_745),
.B(n_229),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_631),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_703),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_666),
.B(n_229),
.Y(n_851)
);

NOR2xp67_ASAP7_75t_L g852 ( 
.A(n_632),
.B(n_566),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_666),
.B(n_230),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_631),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_651),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_646),
.B(n_650),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_710),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_713),
.Y(n_858)
);

O2A1O1Ixp5_ASAP7_75t_L g859 ( 
.A1(n_680),
.A2(n_459),
.B(n_461),
.C(n_301),
.Y(n_859)
);

O2A1O1Ixp5_ASAP7_75t_L g860 ( 
.A1(n_681),
.A2(n_688),
.B(n_690),
.C(n_684),
.Y(n_860)
);

OR2x2_ASAP7_75t_SL g861 ( 
.A(n_746),
.B(n_605),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_641),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_713),
.A2(n_349),
.B1(n_350),
.B2(n_362),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_662),
.B(n_350),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_646),
.B(n_390),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_746),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_634),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_650),
.B(n_392),
.Y(n_868)
);

BUFx8_ASAP7_75t_L g869 ( 
.A(n_706),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_641),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_777),
.B(n_303),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_645),
.B(n_232),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_718),
.B(n_394),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_655),
.B(n_232),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_744),
.B(n_355),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_638),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_665),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_711),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_636),
.Y(n_879)
);

NAND2x1p5_ASAP7_75t_L g880 ( 
.A(n_637),
.B(n_312),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_670),
.B(n_236),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_656),
.B(n_395),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_656),
.B(n_399),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_672),
.B(n_236),
.Y(n_884)
);

AND2x6_ASAP7_75t_SL g885 ( 
.A(n_724),
.B(n_359),
.Y(n_885)
);

NOR2xp67_ASAP7_75t_L g886 ( 
.A(n_638),
.B(n_411),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_644),
.Y(n_887)
);

INVx8_ASAP7_75t_L g888 ( 
.A(n_639),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_679),
.B(n_239),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_753),
.A2(n_411),
.B1(n_410),
.B2(n_404),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_692),
.B(n_370),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_647),
.A2(n_370),
.B1(n_409),
.B2(n_408),
.Y(n_892)
);

AOI21x1_ASAP7_75t_L g893 ( 
.A1(n_681),
.A2(n_328),
.B(n_319),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_686),
.B(n_242),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_647),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_694),
.A2(n_330),
.B(n_335),
.C(n_341),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_643),
.Y(n_897)
);

INVx5_ASAP7_75t_L g898 ( 
.A(n_637),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_711),
.B(n_371),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_695),
.Y(n_900)
);

OAI22xp33_ASAP7_75t_L g901 ( 
.A1(n_777),
.A2(n_408),
.B1(n_407),
.B2(n_405),
.Y(n_901)
);

OR2x6_ASAP7_75t_L g902 ( 
.A(n_767),
.B(n_348),
.Y(n_902)
);

BUFx5_ASAP7_75t_L g903 ( 
.A(n_659),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_657),
.Y(n_904)
);

AND2x2_ASAP7_75t_SL g905 ( 
.A(n_661),
.B(n_353),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_753),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_L g907 ( 
.A(n_649),
.B(n_402),
.C(n_407),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_635),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_684),
.A2(n_410),
.B1(n_404),
.B2(n_246),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_633),
.B(n_403),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_669),
.Y(n_911)
);

INVx8_ASAP7_75t_L g912 ( 
.A(n_659),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_699),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_702),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_707),
.B(n_244),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_669),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_692),
.B(n_403),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_823),
.B(n_633),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_823),
.B(n_633),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_841),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_783),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_793),
.B(n_712),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_782),
.B(n_774),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_841),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_867),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_793),
.B(n_778),
.Y(n_926)
);

OAI21xp33_ASAP7_75t_L g927 ( 
.A1(n_873),
.A2(n_649),
.B(n_661),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_833),
.B(n_738),
.Y(n_928)
);

CKINVDCx16_ASAP7_75t_R g929 ( 
.A(n_838),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_833),
.B(n_668),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_862),
.A2(n_654),
.B(n_697),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_862),
.A2(n_654),
.B(n_697),
.Y(n_932)
);

AOI21x1_ASAP7_75t_L g933 ( 
.A1(n_832),
.A2(n_893),
.B(n_857),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_841),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_837),
.A2(n_709),
.B(n_769),
.C(n_766),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_873),
.B(n_778),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_828),
.B(n_635),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_819),
.B(n_790),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_875),
.B(n_878),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_877),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_855),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_860),
.A2(n_709),
.B(n_673),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_819),
.A2(n_733),
.B(n_751),
.C(n_719),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_800),
.A2(n_756),
.B(n_749),
.Y(n_944)
);

BUFx4f_ASAP7_75t_L g945 ( 
.A(n_795),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_849),
.A2(n_664),
.B(n_660),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_888),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_799),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_905),
.A2(n_668),
.B1(n_635),
.B2(n_659),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_876),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_821),
.B(n_668),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_790),
.B(n_754),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_888),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_SL g954 ( 
.A1(n_905),
.A2(n_630),
.B1(n_683),
.B2(n_651),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_866),
.B(n_683),
.Y(n_955)
);

NOR2x1_ASAP7_75t_L g956 ( 
.A(n_852),
.B(n_737),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_800),
.A2(n_759),
.B(n_758),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_856),
.A2(n_802),
.B(n_813),
.C(n_812),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_817),
.A2(n_671),
.B1(n_719),
.B2(n_733),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_888),
.Y(n_960)
);

BUFx12f_ASAP7_75t_L g961 ( 
.A(n_869),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_847),
.B(n_659),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_912),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_870),
.A2(n_667),
.B(n_733),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_854),
.A2(n_667),
.B(n_751),
.Y(n_965)
);

O2A1O1Ixp5_ASAP7_75t_L g966 ( 
.A1(n_856),
.A2(n_760),
.B(n_737),
.C(n_748),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_792),
.B(n_659),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_863),
.A2(n_827),
.B1(n_789),
.B2(n_892),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_837),
.A2(n_725),
.B(n_747),
.C(n_742),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_839),
.B(n_763),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_779),
.B(n_763),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_854),
.A2(n_667),
.B(n_737),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_869),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_802),
.A2(n_812),
.B1(n_815),
.B2(n_813),
.Y(n_974)
);

OR2x6_ASAP7_75t_SL g975 ( 
.A(n_899),
.B(n_246),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_804),
.B(n_717),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_787),
.A2(n_726),
.B(n_723),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_863),
.A2(n_671),
.B1(n_727),
.B2(n_743),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_844),
.B(n_671),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_814),
.B(n_906),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_829),
.B(n_671),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_850),
.A2(n_640),
.B(n_637),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_858),
.A2(n_640),
.B(n_637),
.Y(n_983)
);

INVx5_ASAP7_75t_L g984 ( 
.A(n_798),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_904),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_892),
.A2(n_717),
.B1(n_729),
.B2(n_743),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_806),
.A2(n_741),
.B1(n_740),
.B2(n_731),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_801),
.A2(n_808),
.B(n_805),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_809),
.A2(n_741),
.B1(n_740),
.B2(n_731),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_829),
.B(n_700),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_912),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_803),
.B(n_735),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_818),
.A2(n_682),
.B(n_687),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_810),
.B(n_735),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_912),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_891),
.B(n_735),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_891),
.B(n_735),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_917),
.B(n_700),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_794),
.B(n_700),
.Y(n_999)
);

NOR2x1_ASAP7_75t_R g1000 ( 
.A(n_897),
.B(n_345),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_901),
.A2(n_384),
.B(n_397),
.C(n_398),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_842),
.A2(n_687),
.B(n_682),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_910),
.B(n_904),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_780),
.A2(n_687),
.B1(n_757),
.B2(n_715),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_882),
.B(n_715),
.Y(n_1005)
);

BUFx8_ASAP7_75t_SL g1006 ( 
.A(n_871),
.Y(n_1006)
);

XOR2x2_ASAP7_75t_R g1007 ( 
.A(n_796),
.B(n_18),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_859),
.A2(n_345),
.B(n_352),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_784),
.A2(n_761),
.B(n_757),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_883),
.B(n_715),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_883),
.B(n_757),
.Y(n_1011)
);

CKINVDCx8_ASAP7_75t_R g1012 ( 
.A(n_885),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_SL g1013 ( 
.A(n_798),
.B(n_352),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_816),
.B(n_357),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_898),
.Y(n_1015)
);

NAND2x1p5_ASAP7_75t_L g1016 ( 
.A(n_898),
.B(n_785),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_825),
.B(n_357),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_886),
.B(n_358),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_807),
.A2(n_360),
.B(n_364),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_908),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_822),
.B(n_360),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_898),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_898),
.Y(n_1023)
);

AND2x4_ASAP7_75t_SL g1024 ( 
.A(n_871),
.B(n_297),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_900),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_825),
.B(n_364),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_798),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_SL g1028 ( 
.A1(n_788),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_879),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_840),
.B(n_368),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_830),
.A2(n_368),
.B(n_372),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_843),
.A2(n_372),
.B(n_388),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_887),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_845),
.A2(n_393),
.B(n_385),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_872),
.A2(n_380),
.B(n_377),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_798),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_835),
.A2(n_333),
.B1(n_332),
.B2(n_331),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_859),
.A2(n_327),
.B(n_326),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_846),
.B(n_251),
.Y(n_1039)
);

AO21x1_ASAP7_75t_L g1040 ( 
.A1(n_865),
.A2(n_316),
.B(n_309),
.Y(n_1040)
);

OAI22x1_ASAP7_75t_L g1041 ( 
.A1(n_868),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_874),
.A2(n_296),
.B(n_318),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_798),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_881),
.A2(n_286),
.B(n_260),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_868),
.A2(n_811),
.B1(n_826),
.B2(n_820),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_884),
.A2(n_298),
.B(n_261),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_851),
.B(n_259),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_853),
.B(n_263),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_834),
.B(n_309),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_913),
.B(n_271),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_L g1051 ( 
.A(n_791),
.B(n_834),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_914),
.B(n_831),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_895),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_889),
.A2(n_307),
.B(n_280),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_911),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_916),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_864),
.B(n_39),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_894),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_903),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_915),
.A2(n_325),
.B(n_316),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_902),
.B(n_44),
.Y(n_1061)
);

OR2x6_ASAP7_75t_L g1062 ( 
.A(n_824),
.B(n_325),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_848),
.A2(n_325),
.B(n_309),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_836),
.A2(n_325),
.B(n_112),
.Y(n_1064)
);

OAI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_890),
.A2(n_50),
.B(n_51),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_781),
.B(n_50),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_958),
.A2(n_896),
.B(n_909),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_974),
.B(n_781),
.Y(n_1068)
);

AND3x4_ASAP7_75t_L g1069 ( 
.A(n_1061),
.B(n_907),
.C(n_861),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_938),
.A2(n_902),
.B(n_880),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_941),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_923),
.B(n_786),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_921),
.Y(n_1073)
);

AO21x1_ASAP7_75t_L g1074 ( 
.A1(n_936),
.A2(n_880),
.B(n_786),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_L g1075 ( 
.A(n_1003),
.B(n_797),
.C(n_57),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_966),
.A2(n_903),
.B(n_57),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_927),
.B(n_918),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_922),
.B(n_903),
.Y(n_1078)
);

AO21x2_ASAP7_75t_L g1079 ( 
.A1(n_1040),
.A2(n_903),
.B(n_125),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_925),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_950),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_963),
.B(n_106),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_976),
.B(n_56),
.Y(n_1083)
);

O2A1O1Ixp5_ASAP7_75t_L g1084 ( 
.A1(n_926),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1005),
.A2(n_62),
.B(n_63),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_930),
.B(n_66),
.Y(n_1086)
);

AOI21x1_ASAP7_75t_L g1087 ( 
.A1(n_1010),
.A2(n_133),
.B(n_190),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_985),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1011),
.A2(n_66),
.B(n_67),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_942),
.A2(n_135),
.B(n_184),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_928),
.B(n_952),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1045),
.B(n_68),
.Y(n_1092)
);

OAI22x1_ASAP7_75t_L g1093 ( 
.A1(n_1061),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_998),
.A2(n_81),
.B(n_88),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_919),
.B(n_94),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_924),
.B(n_953),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1058),
.B(n_97),
.Y(n_1097)
);

OR2x6_ASAP7_75t_L g1098 ( 
.A(n_961),
.B(n_199),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_924),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_924),
.B(n_953),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_967),
.A2(n_141),
.B(n_146),
.Y(n_1101)
);

NOR2xp67_ASAP7_75t_L g1102 ( 
.A(n_951),
.B(n_147),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_940),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_953),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1025),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_937),
.B(n_151),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1052),
.B(n_176),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1001),
.A2(n_179),
.B(n_1017),
.C(n_1014),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_999),
.A2(n_997),
.B(n_996),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_945),
.B(n_949),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1006),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_945),
.B(n_979),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1026),
.A2(n_1065),
.B(n_935),
.C(n_968),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_929),
.Y(n_1114)
);

BUFx12f_ASAP7_75t_L g1115 ( 
.A(n_973),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_931),
.A2(n_932),
.B(n_977),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_SL g1117 ( 
.A(n_1062),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_970),
.B(n_971),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_946),
.A2(n_988),
.B(n_944),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1021),
.B(n_1030),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_977),
.A2(n_992),
.B(n_962),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_948),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1055),
.Y(n_1123)
);

NAND2x1p5_ASAP7_75t_L g1124 ( 
.A(n_963),
.B(n_991),
.Y(n_1124)
);

AO22x1_ASAP7_75t_L g1125 ( 
.A1(n_1007),
.A2(n_955),
.B1(n_1066),
.B2(n_1057),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1029),
.B(n_1033),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1053),
.B(n_1056),
.Y(n_1127)
);

AOI221x1_ASAP7_75t_L g1128 ( 
.A1(n_1038),
.A2(n_959),
.B1(n_1008),
.B2(n_1041),
.C(n_1064),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_957),
.A2(n_1059),
.B(n_965),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_987),
.A2(n_989),
.A3(n_986),
.B(n_1060),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_980),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_969),
.Y(n_1132)
);

AND3x1_ASAP7_75t_SL g1133 ( 
.A(n_975),
.B(n_1012),
.C(n_954),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_1020),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1013),
.A2(n_964),
.B(n_972),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_986),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1008),
.A2(n_994),
.B(n_987),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_990),
.B(n_991),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_978),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_981),
.B(n_1048),
.Y(n_1140)
);

OAI22x1_ASAP7_75t_L g1141 ( 
.A1(n_1051),
.A2(n_1049),
.B1(n_1037),
.B2(n_1018),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1039),
.B(n_1047),
.Y(n_1142)
);

AND3x4_ASAP7_75t_L g1143 ( 
.A(n_956),
.B(n_1000),
.C(n_1028),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1020),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1050),
.A2(n_934),
.B1(n_995),
.B2(n_1062),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_934),
.B(n_995),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1020),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1059),
.A2(n_1016),
.B(n_993),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1035),
.A2(n_1046),
.B(n_1054),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_L g1150 ( 
.A(n_920),
.B(n_947),
.Y(n_1150)
);

INVxp67_ASAP7_75t_SL g1151 ( 
.A(n_995),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_920),
.B(n_947),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1027),
.A2(n_984),
.B(n_1044),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_960),
.B(n_1015),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1049),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1024),
.B(n_960),
.Y(n_1156)
);

NAND2x1p5_ASAP7_75t_L g1157 ( 
.A(n_1022),
.B(n_1027),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1002),
.A2(n_1004),
.B(n_983),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1063),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1160)
);

NAND3xp33_ASAP7_75t_L g1161 ( 
.A(n_1042),
.B(n_1031),
.C(n_1019),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1023),
.B(n_1036),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_984),
.B(n_1023),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_982),
.A2(n_1032),
.B(n_1034),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1043),
.A2(n_958),
.B(n_860),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_958),
.B(n_974),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_958),
.B(n_974),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_928),
.B(n_657),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_933),
.A2(n_966),
.B(n_1009),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_1040),
.A2(n_958),
.A3(n_943),
.B(n_987),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_938),
.A2(n_922),
.B(n_958),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_958),
.A2(n_860),
.B(n_938),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_974),
.A2(n_958),
.B(n_873),
.C(n_819),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_921),
.Y(n_1174)
);

AOI21xp33_ASAP7_75t_L g1175 ( 
.A1(n_974),
.A2(n_958),
.B(n_938),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_958),
.B(n_974),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_938),
.A2(n_922),
.B(n_958),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_928),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_938),
.A2(n_922),
.B(n_958),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_974),
.B(n_782),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_958),
.B(n_974),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_941),
.Y(n_1182)
);

OA21x2_ASAP7_75t_L g1183 ( 
.A1(n_1040),
.A2(n_942),
.B(n_943),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_938),
.A2(n_922),
.B(n_958),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_939),
.B(n_833),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_933),
.A2(n_966),
.B(n_1009),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_974),
.B(n_782),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_958),
.B(n_974),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_933),
.A2(n_966),
.B(n_1009),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1040),
.A2(n_958),
.A3(n_943),
.B(n_987),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_958),
.B(n_974),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_939),
.B(n_833),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1146),
.B(n_1096),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1104),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1072),
.A2(n_1068),
.B1(n_1069),
.B2(n_1181),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1185),
.B(n_1192),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1118),
.B(n_1071),
.Y(n_1198)
);

AOI21xp33_ASAP7_75t_SL g1199 ( 
.A1(n_1175),
.A2(n_1167),
.B(n_1166),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1176),
.A2(n_1188),
.B(n_1181),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1176),
.A2(n_1191),
.B(n_1188),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1191),
.A2(n_1175),
.B(n_1113),
.C(n_1108),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1080),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1124),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1068),
.A2(n_1092),
.B1(n_1171),
.B2(n_1177),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_1114),
.Y(n_1206)
);

NAND3xp33_ASAP7_75t_SL g1207 ( 
.A(n_1092),
.B(n_1067),
.C(n_1143),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_SL g1208 ( 
.A(n_1117),
.B(n_1075),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1146),
.B(n_1096),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1178),
.B(n_1142),
.Y(n_1210)
);

INVx5_ASAP7_75t_L g1211 ( 
.A(n_1115),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1182),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1142),
.B(n_1088),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1100),
.B(n_1099),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1100),
.B(n_1099),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1091),
.B(n_1168),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1081),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1104),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1086),
.B(n_1125),
.Y(n_1219)
);

INVx5_ASAP7_75t_L g1220 ( 
.A(n_1104),
.Y(n_1220)
);

NOR3xp33_ASAP7_75t_L g1221 ( 
.A(n_1112),
.B(n_1120),
.C(n_1140),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1103),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1134),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1077),
.A2(n_1132),
.B1(n_1133),
.B2(n_1093),
.Y(n_1224)
);

NOR2xp67_ASAP7_75t_L g1225 ( 
.A(n_1095),
.B(n_1179),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1078),
.A2(n_1184),
.B(n_1116),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1083),
.B(n_1105),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1123),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1144),
.B(n_1098),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1083),
.B(n_1147),
.Y(n_1230)
);

OAI21xp33_ASAP7_75t_SL g1231 ( 
.A1(n_1172),
.A2(n_1078),
.B(n_1139),
.Y(n_1231)
);

INVx4_ASAP7_75t_L g1232 ( 
.A(n_1111),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1150),
.B(n_1110),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1122),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1131),
.B(n_1174),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1117),
.A2(n_1126),
.B1(n_1127),
.B2(n_1141),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1152),
.B(n_1154),
.Y(n_1237)
);

CKINVDCx14_ASAP7_75t_R g1238 ( 
.A(n_1098),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1070),
.B(n_1127),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1085),
.A2(n_1089),
.B(n_1076),
.C(n_1137),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1152),
.B(n_1154),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1151),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1124),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1109),
.A2(n_1135),
.B(n_1106),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1156),
.B(n_1155),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1163),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1109),
.A2(n_1106),
.B(n_1165),
.Y(n_1247)
);

NOR2x1_ASAP7_75t_SL g1248 ( 
.A(n_1145),
.B(n_1138),
.Y(n_1248)
);

OAI21xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1136),
.A2(n_1107),
.B(n_1121),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1089),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1070),
.B(n_1138),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1082),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1107),
.A2(n_1102),
.B1(n_1097),
.B2(n_1074),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1084),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1162),
.B(n_1160),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1160),
.B(n_1162),
.Y(n_1256)
);

NOR2xp67_ASAP7_75t_L g1257 ( 
.A(n_1161),
.B(n_1153),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1163),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_SL g1259 ( 
.A1(n_1149),
.A2(n_1164),
.B(n_1101),
.C(n_1094),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1157),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1159),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1128),
.A2(n_1129),
.B(n_1119),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1157),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1170),
.Y(n_1264)
);

BUFx8_ASAP7_75t_L g1265 ( 
.A(n_1082),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1170),
.B(n_1190),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1148),
.Y(n_1267)
);

BUFx4f_ASAP7_75t_L g1268 ( 
.A(n_1183),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1190),
.B(n_1130),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1087),
.Y(n_1270)
);

BUFx12f_ASAP7_75t_L g1271 ( 
.A(n_1101),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1090),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1183),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1130),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1079),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1169),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1158),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1186),
.A2(n_1180),
.B1(n_1187),
.B2(n_974),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1189),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1173),
.A2(n_1167),
.B(n_1166),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1115),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1080),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1283)
);

INVxp67_ASAP7_75t_SL g1284 ( 
.A(n_1088),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1180),
.A2(n_1187),
.B1(n_974),
.B2(n_873),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1180),
.A2(n_1187),
.B1(n_974),
.B2(n_1173),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1071),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1173),
.A2(n_1167),
.B(n_1166),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1180),
.A2(n_1187),
.B1(n_974),
.B2(n_1173),
.Y(n_1291)
);

BUFx10_ASAP7_75t_L g1292 ( 
.A(n_1096),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1080),
.Y(n_1293)
);

AOI222xp33_ASAP7_75t_L g1294 ( 
.A1(n_1072),
.A2(n_905),
.B1(n_927),
.B2(n_1187),
.C1(n_1180),
.C2(n_1061),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1146),
.B(n_1096),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1080),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1180),
.A2(n_1187),
.B1(n_974),
.B2(n_1173),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1173),
.A2(n_958),
.B(n_1166),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1185),
.B(n_1192),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1180),
.A2(n_974),
.B(n_958),
.C(n_1187),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1180),
.A2(n_1187),
.B1(n_974),
.B2(n_873),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1088),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1080),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1185),
.B(n_1192),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1180),
.B(n_974),
.Y(n_1306)
);

OR2x6_ASAP7_75t_SL g1307 ( 
.A(n_1168),
.B(n_638),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1185),
.B(n_1192),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1178),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1173),
.A2(n_1167),
.B(n_1166),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1104),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1124),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1146),
.B(n_1096),
.Y(n_1315)
);

AO22x1_ASAP7_75t_L g1316 ( 
.A1(n_1069),
.A2(n_649),
.B1(n_638),
.B2(n_839),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1185),
.B(n_1192),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1319)
);

BUFx12f_ASAP7_75t_L g1320 ( 
.A(n_1115),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1080),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1080),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1173),
.A2(n_1167),
.B(n_1166),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1173),
.A2(n_1167),
.B(n_1166),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1114),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1080),
.Y(n_1326)
);

CKINVDCx11_ASAP7_75t_R g1327 ( 
.A(n_1114),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1185),
.B(n_1192),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1080),
.Y(n_1329)
);

O2A1O1Ixp5_ASAP7_75t_L g1330 ( 
.A1(n_1180),
.A2(n_1187),
.B(n_1173),
.C(n_1166),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1115),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1115),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1180),
.B(n_1187),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1180),
.A2(n_974),
.B(n_958),
.C(n_1187),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1104),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1073),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1180),
.A2(n_1187),
.B1(n_974),
.B2(n_1173),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1193),
.B(n_1209),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1302),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1196),
.B(n_1278),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1246),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1203),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1196),
.B(n_1278),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1300),
.B(n_1336),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1327),
.Y(n_1347)
);

AO21x1_ASAP7_75t_L g1348 ( 
.A1(n_1339),
.A2(n_1291),
.B(n_1287),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1246),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1284),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1219),
.A2(n_1297),
.B1(n_1208),
.B2(n_1339),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1208),
.A2(n_1238),
.B1(n_1194),
.B2(n_1319),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1288),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1271),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1267),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1281),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1198),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1294),
.A2(n_1207),
.B1(n_1301),
.B2(n_1286),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1286),
.A2(n_1301),
.B1(n_1335),
.B2(n_1303),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1294),
.A2(n_1306),
.B1(n_1224),
.B2(n_1309),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1224),
.A2(n_1317),
.B1(n_1289),
.B2(n_1285),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1283),
.A2(n_1334),
.B1(n_1333),
.B2(n_1310),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1246),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1222),
.Y(n_1364)
);

AO21x1_ASAP7_75t_SL g1365 ( 
.A1(n_1298),
.A2(n_1269),
.B(n_1250),
.Y(n_1365)
);

BUFx2_ASAP7_75t_SL g1366 ( 
.A(n_1220),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1298),
.B(n_1330),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1239),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1268),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1307),
.A2(n_1197),
.B1(n_1213),
.B2(n_1199),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1262),
.A2(n_1247),
.B(n_1226),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1251),
.B(n_1299),
.Y(n_1372)
);

CKINVDCx6p67_ASAP7_75t_R g1373 ( 
.A(n_1211),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1282),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1225),
.A2(n_1202),
.B(n_1324),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1293),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1296),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1258),
.Y(n_1378)
);

NOR2x1_ASAP7_75t_R g1379 ( 
.A(n_1211),
.B(n_1320),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1265),
.A2(n_1236),
.B1(n_1338),
.B2(n_1234),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1220),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1267),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1304),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1316),
.B(n_1212),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1210),
.B(n_1305),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1267),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1274),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1308),
.Y(n_1388)
);

INVx4_ASAP7_75t_L g1389 ( 
.A(n_1220),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1273),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1321),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1280),
.A2(n_1323),
.B1(n_1290),
.B2(n_1312),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1273),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1322),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1326),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1228),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1329),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1206),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1223),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1227),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1223),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1318),
.B(n_1328),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1216),
.B(n_1221),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1230),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1266),
.A2(n_1275),
.B(n_1257),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_1195),
.Y(n_1406)
);

BUFx2_ASAP7_75t_SL g1407 ( 
.A(n_1233),
.Y(n_1407)
);

INVx8_ASAP7_75t_L g1408 ( 
.A(n_1211),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1233),
.A2(n_1229),
.B1(n_1225),
.B2(n_1325),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1331),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1255),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1264),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1199),
.A2(n_1201),
.B1(n_1200),
.B2(n_1205),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_SL g1414 ( 
.A1(n_1240),
.A2(n_1248),
.B(n_1205),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1332),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1249),
.A2(n_1253),
.B(n_1231),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1258),
.Y(n_1417)
);

CKINVDCx11_ASAP7_75t_R g1418 ( 
.A(n_1232),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1231),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1292),
.Y(n_1420)
);

BUFx8_ASAP7_75t_L g1421 ( 
.A(n_1223),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1279),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1311),
.A2(n_1235),
.B1(n_1253),
.B2(n_1245),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1249),
.A2(n_1245),
.B1(n_1242),
.B2(n_1256),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1193),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1272),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1237),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1241),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1263),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1254),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1217),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1260),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1295),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1276),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1259),
.A2(n_1277),
.B(n_1313),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1195),
.Y(n_1436)
);

INVxp33_ASAP7_75t_L g1437 ( 
.A(n_1315),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_1232),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1195),
.B(n_1337),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1292),
.A2(n_1204),
.B1(n_1314),
.B2(n_1243),
.Y(n_1440)
);

BUFx8_ASAP7_75t_L g1441 ( 
.A(n_1214),
.Y(n_1441)
);

CKINVDCx6p67_ASAP7_75t_R g1442 ( 
.A(n_1337),
.Y(n_1442)
);

NAND2x1p5_ASAP7_75t_L g1443 ( 
.A(n_1260),
.B(n_1263),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1215),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1204),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1218),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1218),
.B(n_1337),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1203),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1219),
.A2(n_1072),
.B1(n_905),
.B2(n_722),
.Y(n_1449)
);

AO21x2_ASAP7_75t_L g1450 ( 
.A1(n_1244),
.A2(n_1270),
.B(n_1247),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1268),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1327),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1286),
.A2(n_1301),
.B1(n_974),
.B2(n_1196),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1203),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1219),
.A2(n_1072),
.B1(n_905),
.B2(n_722),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1196),
.B(n_1278),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1203),
.Y(n_1457)
);

AO21x1_ASAP7_75t_SL g1458 ( 
.A1(n_1278),
.A2(n_1167),
.B(n_1166),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1203),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1219),
.A2(n_1072),
.B1(n_905),
.B2(n_722),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1302),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1223),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1220),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1271),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1327),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1203),
.Y(n_1466)
);

INVxp67_ASAP7_75t_SL g1467 ( 
.A(n_1256),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1271),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1294),
.A2(n_905),
.B1(n_1072),
.B2(n_1207),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1203),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1203),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1196),
.B(n_1278),
.Y(n_1472)
);

NAND2x1p5_ASAP7_75t_L g1473 ( 
.A(n_1252),
.B(n_1268),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1302),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1294),
.A2(n_905),
.B1(n_1072),
.B2(n_1207),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1196),
.B(n_1278),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1203),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1203),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1194),
.B(n_1283),
.Y(n_1479)
);

AO21x1_ASAP7_75t_L g1480 ( 
.A1(n_1339),
.A2(n_1291),
.B(n_1287),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_1311),
.Y(n_1481)
);

BUFx4f_ASAP7_75t_SL g1482 ( 
.A(n_1281),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1268),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1286),
.A2(n_1301),
.B1(n_839),
.B2(n_974),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1203),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1219),
.A2(n_1072),
.B1(n_905),
.B2(n_722),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1302),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1203),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1203),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1193),
.B(n_1209),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1196),
.B(n_1278),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1203),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1302),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1271),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1261),
.Y(n_1495)
);

AOI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1413),
.A2(n_1480),
.B(n_1348),
.Y(n_1496)
);

NAND2x1_ASAP7_75t_L g1497 ( 
.A(n_1414),
.B(n_1419),
.Y(n_1497)
);

CKINVDCx14_ASAP7_75t_R g1498 ( 
.A(n_1398),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1479),
.B(n_1357),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1419),
.Y(n_1500)
);

AO21x2_ASAP7_75t_L g1501 ( 
.A1(n_1416),
.A2(n_1414),
.B(n_1375),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1368),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1430),
.Y(n_1503)
);

AO31x2_ASAP7_75t_L g1504 ( 
.A1(n_1392),
.A2(n_1348),
.A3(n_1480),
.B(n_1387),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1372),
.B(n_1342),
.Y(n_1505)
);

NAND2x1p5_ASAP7_75t_L g1506 ( 
.A(n_1354),
.B(n_1464),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1467),
.B(n_1427),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1495),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1484),
.A2(n_1453),
.B(n_1358),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1367),
.A2(n_1426),
.B(n_1434),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1421),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1367),
.A2(n_1426),
.B(n_1434),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1345),
.B(n_1456),
.Y(n_1513)
);

AOI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1359),
.A2(n_1435),
.B(n_1371),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1350),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1472),
.B(n_1476),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1435),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1421),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1341),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_1351),
.B(n_1362),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1398),
.B(n_1428),
.Y(n_1521)
);

AO21x2_ASAP7_75t_L g1522 ( 
.A1(n_1450),
.A2(n_1370),
.B(n_1412),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1422),
.A2(n_1393),
.B(n_1472),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1476),
.B(n_1491),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1491),
.A2(n_1346),
.B1(n_1460),
.B2(n_1455),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1388),
.B(n_1431),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1393),
.A2(n_1346),
.B(n_1423),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1396),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1435),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1405),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1355),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1438),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1405),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1344),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1355),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1364),
.Y(n_1536)
);

OR2x6_ASAP7_75t_L g1537 ( 
.A(n_1407),
.B(n_1369),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1374),
.Y(n_1538)
);

CKINVDCx6p67_ASAP7_75t_R g1539 ( 
.A(n_1373),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1376),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1377),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1383),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1391),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1390),
.A2(n_1371),
.B(n_1386),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1365),
.B(n_1458),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1361),
.A2(n_1360),
.B(n_1475),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1394),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1395),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1449),
.A2(n_1486),
.B1(n_1469),
.B2(n_1380),
.Y(n_1549)
);

AO21x2_ASAP7_75t_L g1550 ( 
.A1(n_1450),
.A2(n_1409),
.B(n_1454),
.Y(n_1550)
);

OA21x2_ASAP7_75t_L g1551 ( 
.A1(n_1397),
.A2(n_1477),
.B(n_1478),
.Y(n_1551)
);

NAND3xp33_ASAP7_75t_SL g1552 ( 
.A(n_1352),
.B(n_1347),
.C(n_1452),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1365),
.B(n_1458),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1448),
.Y(n_1554)
);

INVx5_ASAP7_75t_SL g1555 ( 
.A(n_1373),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1382),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1404),
.B(n_1411),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1402),
.B(n_1457),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1461),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1402),
.B(n_1459),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1385),
.B(n_1400),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1466),
.Y(n_1562)
);

AO21x2_ASAP7_75t_L g1563 ( 
.A1(n_1470),
.A2(n_1485),
.B(n_1471),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1488),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1489),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1492),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1390),
.A2(n_1371),
.B(n_1386),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1390),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1451),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1421),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1483),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1474),
.B(n_1487),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1473),
.A2(n_1494),
.B(n_1468),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1493),
.B(n_1424),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1354),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1356),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1445),
.Y(n_1577)
);

INVx2_ASAP7_75t_SL g1578 ( 
.A(n_1408),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1399),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1464),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1399),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1464),
.B(n_1494),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1468),
.Y(n_1583)
);

AO21x2_ASAP7_75t_L g1584 ( 
.A1(n_1403),
.A2(n_1436),
.B(n_1446),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1432),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1439),
.B(n_1447),
.Y(n_1586)
);

CKINVDCx14_ASAP7_75t_R g1587 ( 
.A(n_1347),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1432),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1432),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1447),
.B(n_1353),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1407),
.Y(n_1591)
);

AO21x2_ASAP7_75t_L g1592 ( 
.A1(n_1384),
.A2(n_1340),
.B(n_1490),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1429),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1429),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1343),
.Y(n_1595)
);

NAND2x1_ASAP7_75t_L g1596 ( 
.A(n_1389),
.B(n_1406),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1343),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1438),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1343),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1349),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1349),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1481),
.B(n_1401),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1462),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1442),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1408),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1497),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1500),
.B(n_1444),
.Y(n_1607)
);

NAND4xp25_ASAP7_75t_L g1608 ( 
.A(n_1509),
.B(n_1418),
.C(n_1440),
.D(n_1465),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1551),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1505),
.B(n_1558),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1497),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1576),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1560),
.B(n_1433),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1520),
.A2(n_1420),
.B1(n_1356),
.B2(n_1437),
.C(n_1408),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1511),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1523),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1551),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1545),
.B(n_1381),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1515),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1511),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1513),
.B(n_1516),
.Y(n_1621)
);

OAI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1546),
.A2(n_1437),
.B1(n_1425),
.B2(n_1420),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1507),
.B(n_1463),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1551),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1518),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1524),
.B(n_1586),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1513),
.B(n_1381),
.Y(n_1627)
);

OAI222xp33_ASAP7_75t_L g1628 ( 
.A1(n_1525),
.A2(n_1443),
.B1(n_1465),
.B2(n_1452),
.C1(n_1490),
.C2(n_1340),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1496),
.A2(n_1389),
.B(n_1443),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1519),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1586),
.B(n_1417),
.Y(n_1631)
);

INVx4_ASAP7_75t_L g1632 ( 
.A(n_1506),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1590),
.B(n_1417),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1590),
.B(n_1417),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_1518),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1559),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1602),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1499),
.B(n_1410),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1516),
.B(n_1366),
.Y(n_1639)
);

OAI221xp5_ASAP7_75t_L g1640 ( 
.A1(n_1549),
.A2(n_1410),
.B1(n_1415),
.B2(n_1366),
.C(n_1378),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1572),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1563),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1563),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1503),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1584),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1523),
.B(n_1363),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1570),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1523),
.B(n_1545),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1503),
.Y(n_1649)
);

OA332x1_ASAP7_75t_L g1650 ( 
.A1(n_1498),
.A2(n_1415),
.A3(n_1482),
.B1(n_1379),
.B2(n_1441),
.B3(n_1340),
.C1(n_1490),
.C2(n_1363),
.Y(n_1650)
);

INVxp67_ASAP7_75t_SL g1651 ( 
.A(n_1523),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1535),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1603),
.Y(n_1653)
);

OAI211xp5_ASAP7_75t_SL g1654 ( 
.A1(n_1521),
.A2(n_1363),
.B(n_1441),
.C(n_1532),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1508),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1553),
.B(n_1441),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1557),
.B(n_1577),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1501),
.B(n_1537),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1501),
.B(n_1534),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1517),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_1510),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1501),
.B(n_1534),
.Y(n_1662)
);

INVxp67_ASAP7_75t_SL g1663 ( 
.A(n_1510),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1508),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1496),
.A2(n_1574),
.B1(n_1598),
.B2(n_1526),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1584),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1584),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1541),
.B(n_1543),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1541),
.B(n_1543),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1554),
.B(n_1562),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1576),
.B(n_1587),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1610),
.B(n_1550),
.Y(n_1672)
);

OAI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1665),
.A2(n_1552),
.B1(n_1574),
.B2(n_1506),
.C(n_1536),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1651),
.A2(n_1530),
.B(n_1533),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1626),
.B(n_1569),
.Y(n_1675)
);

OAI221xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1616),
.A2(n_1591),
.B1(n_1571),
.B2(n_1569),
.C(n_1537),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1641),
.B(n_1504),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1626),
.B(n_1571),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1640),
.A2(n_1506),
.B1(n_1555),
.B2(n_1539),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1619),
.B(n_1504),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1630),
.B(n_1504),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1608),
.A2(n_1592),
.B1(n_1527),
.B2(n_1582),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1636),
.B(n_1504),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1621),
.B(n_1554),
.Y(n_1684)
);

AOI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1616),
.A2(n_1562),
.B1(n_1565),
.B2(n_1547),
.C(n_1542),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1659),
.B(n_1585),
.C(n_1588),
.Y(n_1686)
);

NAND3xp33_ASAP7_75t_L g1687 ( 
.A(n_1659),
.B(n_1585),
.C(n_1588),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1629),
.A2(n_1537),
.B(n_1596),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1662),
.B(n_1589),
.C(n_1565),
.Y(n_1689)
);

OAI221xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1608),
.A2(n_1614),
.B1(n_1648),
.B2(n_1639),
.C(n_1621),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1668),
.B(n_1538),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1668),
.B(n_1540),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1669),
.B(n_1540),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1662),
.B(n_1589),
.C(n_1591),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1658),
.A2(n_1596),
.B(n_1522),
.Y(n_1695)
);

NAND3xp33_ASAP7_75t_L g1696 ( 
.A(n_1653),
.B(n_1527),
.C(n_1547),
.Y(n_1696)
);

OA21x2_ASAP7_75t_L g1697 ( 
.A1(n_1642),
.A2(n_1530),
.B(n_1533),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1669),
.B(n_1542),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1670),
.B(n_1548),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1670),
.B(n_1548),
.Y(n_1700)
);

NOR3xp33_ASAP7_75t_L g1701 ( 
.A(n_1654),
.B(n_1514),
.C(n_1583),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1633),
.B(n_1556),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1634),
.B(n_1568),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1634),
.B(n_1568),
.Y(n_1704)
);

NOR3xp33_ASAP7_75t_L g1705 ( 
.A(n_1623),
.B(n_1514),
.C(n_1575),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1657),
.B(n_1564),
.Y(n_1706)
);

NAND3xp33_ASAP7_75t_L g1707 ( 
.A(n_1645),
.B(n_1527),
.C(n_1566),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1631),
.B(n_1527),
.Y(n_1708)
);

OA21x2_ASAP7_75t_L g1709 ( 
.A1(n_1642),
.A2(n_1544),
.B(n_1567),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1631),
.B(n_1522),
.Y(n_1710)
);

AND2x2_ASAP7_75t_SL g1711 ( 
.A(n_1656),
.B(n_1510),
.Y(n_1711)
);

OAI21xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1628),
.A2(n_1604),
.B(n_1580),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1637),
.B(n_1564),
.Y(n_1713)
);

NAND3xp33_ASAP7_75t_L g1714 ( 
.A(n_1666),
.B(n_1566),
.C(n_1597),
.Y(n_1714)
);

NAND3xp33_ASAP7_75t_L g1715 ( 
.A(n_1667),
.B(n_1599),
.C(n_1594),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1644),
.Y(n_1716)
);

OAI221xp5_ASAP7_75t_SL g1717 ( 
.A1(n_1661),
.A2(n_1561),
.B1(n_1529),
.B2(n_1600),
.C(n_1593),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1607),
.B(n_1529),
.Y(n_1718)
);

NAND3xp33_ASAP7_75t_L g1719 ( 
.A(n_1643),
.B(n_1593),
.C(n_1601),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1607),
.B(n_1512),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1663),
.A2(n_1561),
.B1(n_1582),
.B2(n_1528),
.C(n_1502),
.Y(n_1721)
);

NAND3xp33_ASAP7_75t_L g1722 ( 
.A(n_1643),
.B(n_1595),
.C(n_1597),
.Y(n_1722)
);

OAI221xp5_ASAP7_75t_SL g1723 ( 
.A1(n_1622),
.A2(n_1600),
.B1(n_1601),
.B2(n_1595),
.C(n_1570),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1613),
.B(n_1512),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1644),
.B(n_1579),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_SL g1726 ( 
.A1(n_1656),
.A2(n_1605),
.B(n_1578),
.Y(n_1726)
);

OAI21xp5_ASAP7_75t_SL g1727 ( 
.A1(n_1656),
.A2(n_1605),
.B(n_1578),
.Y(n_1727)
);

NOR3xp33_ASAP7_75t_L g1728 ( 
.A(n_1660),
.B(n_1573),
.C(n_1531),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1649),
.B(n_1581),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1649),
.B(n_1581),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1716),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1697),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1674),
.Y(n_1733)
);

BUFx3_ASAP7_75t_L g1734 ( 
.A(n_1674),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1720),
.B(n_1672),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1697),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1706),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1684),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1691),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1674),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1672),
.B(n_1652),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1677),
.B(n_1627),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1728),
.B(n_1606),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1711),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1682),
.A2(n_1696),
.B1(n_1673),
.B2(n_1592),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1692),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1693),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1711),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1698),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1699),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1709),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1708),
.B(n_1606),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1680),
.B(n_1609),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1708),
.B(n_1606),
.Y(n_1754)
);

INVxp67_ASAP7_75t_SL g1755 ( 
.A(n_1681),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1700),
.Y(n_1756)
);

NOR2xp67_ASAP7_75t_L g1757 ( 
.A(n_1695),
.B(n_1611),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1683),
.B(n_1609),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1709),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1709),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1724),
.B(n_1618),
.Y(n_1761)
);

BUFx2_ASAP7_75t_L g1762 ( 
.A(n_1718),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1685),
.B(n_1689),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1714),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1705),
.B(n_1710),
.Y(n_1765)
);

NAND2x1p5_ASAP7_75t_L g1766 ( 
.A(n_1688),
.B(n_1632),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1713),
.Y(n_1767)
);

NOR2xp67_ASAP7_75t_L g1768 ( 
.A(n_1719),
.B(n_1617),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1686),
.B(n_1617),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1722),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1707),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1687),
.B(n_1624),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1701),
.B(n_1646),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1731),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1744),
.B(n_1675),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1744),
.B(n_1761),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1735),
.B(n_1678),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1764),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1731),
.Y(n_1779)
);

INVx2_ASAP7_75t_SL g1780 ( 
.A(n_1733),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1767),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1735),
.B(n_1703),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1763),
.B(n_1717),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1770),
.B(n_1721),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1767),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1770),
.B(n_1612),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1763),
.B(n_1725),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1764),
.B(n_1655),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1762),
.B(n_1703),
.Y(n_1789)
);

AND3x2_ASAP7_75t_L g1790 ( 
.A(n_1771),
.B(n_1671),
.C(n_1638),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1737),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1733),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1737),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1762),
.B(n_1704),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1733),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1768),
.B(n_1694),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1734),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1739),
.Y(n_1798)
);

NOR2x1_ASAP7_75t_L g1799 ( 
.A(n_1734),
.B(n_1615),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1734),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1740),
.Y(n_1801)
);

INVx2_ASAP7_75t_SL g1802 ( 
.A(n_1743),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1769),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1739),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1740),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1766),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1746),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1742),
.B(n_1729),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1746),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1747),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1742),
.B(n_1730),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1747),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1771),
.B(n_1655),
.Y(n_1813)
);

OAI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1745),
.A2(n_1690),
.B1(n_1723),
.B2(n_1712),
.C(n_1676),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1759),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1741),
.B(n_1702),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1771),
.B(n_1664),
.Y(n_1817)
);

NOR2x1_ASAP7_75t_L g1818 ( 
.A(n_1768),
.B(n_1615),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1765),
.B(n_1715),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1777),
.B(n_1782),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1774),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1778),
.B(n_1738),
.Y(n_1822)
);

OAI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1814),
.A2(n_1745),
.B1(n_1765),
.B2(n_1748),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1787),
.B(n_1769),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1778),
.B(n_1738),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1777),
.B(n_1773),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1774),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1787),
.B(n_1772),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1788),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1779),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1777),
.B(n_1773),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1782),
.B(n_1773),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1783),
.B(n_1749),
.Y(n_1833)
);

OA21x2_ASAP7_75t_L g1834 ( 
.A1(n_1784),
.A2(n_1736),
.B(n_1732),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1783),
.B(n_1749),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1784),
.B(n_1772),
.Y(n_1836)
);

NAND3xp33_ASAP7_75t_SL g1837 ( 
.A(n_1814),
.B(n_1748),
.C(n_1766),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1779),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1796),
.A2(n_1748),
.B1(n_1773),
.B2(n_1592),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1819),
.B(n_1753),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1788),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1782),
.B(n_1752),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1801),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1801),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1803),
.B(n_1750),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1803),
.Y(n_1846)
);

OAI21xp33_ASAP7_75t_L g1847 ( 
.A1(n_1819),
.A2(n_1796),
.B(n_1813),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1790),
.B(n_1750),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1781),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1781),
.Y(n_1850)
);

INVx4_ASAP7_75t_L g1851 ( 
.A(n_1790),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1785),
.B(n_1756),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1789),
.B(n_1752),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1798),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1789),
.B(n_1794),
.Y(n_1855)
);

INVx1_ASAP7_75t_SL g1856 ( 
.A(n_1786),
.Y(n_1856)
);

INVx1_ASAP7_75t_SL g1857 ( 
.A(n_1806),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1785),
.B(n_1756),
.Y(n_1858)
);

NOR2x1_ASAP7_75t_L g1859 ( 
.A(n_1818),
.B(n_1620),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1789),
.B(n_1794),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1813),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1817),
.B(n_1755),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1794),
.B(n_1752),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1801),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1817),
.B(n_1753),
.Y(n_1865)
);

BUFx2_ASAP7_75t_L g1866 ( 
.A(n_1818),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1798),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1791),
.Y(n_1868)
);

NOR2x1_ASAP7_75t_L g1869 ( 
.A(n_1799),
.B(n_1620),
.Y(n_1869)
);

INVxp33_ASAP7_75t_L g1870 ( 
.A(n_1799),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1804),
.B(n_1758),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1816),
.B(n_1752),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1827),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1836),
.B(n_1796),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1834),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1834),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1836),
.B(n_1796),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1827),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1830),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1830),
.Y(n_1880)
);

INVx1_ASAP7_75t_SL g1881 ( 
.A(n_1856),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1833),
.B(n_1804),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1838),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1820),
.B(n_1776),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1838),
.Y(n_1885)
);

AOI22x1_ASAP7_75t_L g1886 ( 
.A1(n_1851),
.A2(n_1612),
.B1(n_1780),
.B2(n_1802),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1823),
.A2(n_1792),
.B1(n_1797),
.B2(n_1795),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_1851),
.B(n_1806),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1820),
.B(n_1776),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1824),
.B(n_1791),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1834),
.Y(n_1891)
);

OAI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1851),
.A2(n_1766),
.B1(n_1806),
.B2(n_1802),
.Y(n_1892)
);

INVx1_ASAP7_75t_SL g1893 ( 
.A(n_1857),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1835),
.B(n_1807),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1824),
.B(n_1807),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_1866),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1821),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1855),
.B(n_1860),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_1866),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1854),
.Y(n_1900)
);

INVx1_ASAP7_75t_SL g1901 ( 
.A(n_1848),
.Y(n_1901)
);

BUFx3_ASAP7_75t_L g1902 ( 
.A(n_1846),
.Y(n_1902)
);

BUFx3_ASAP7_75t_L g1903 ( 
.A(n_1849),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1854),
.Y(n_1904)
);

NAND2xp33_ASAP7_75t_L g1905 ( 
.A(n_1859),
.B(n_1802),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1828),
.B(n_1840),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1828),
.B(n_1793),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1847),
.A2(n_1811),
.B1(n_1808),
.B2(n_1754),
.Y(n_1908)
);

INVx1_ASAP7_75t_SL g1909 ( 
.A(n_1840),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1855),
.B(n_1816),
.Y(n_1910)
);

INVx1_ASAP7_75t_SL g1911 ( 
.A(n_1822),
.Y(n_1911)
);

NOR2x1_ASAP7_75t_L g1912 ( 
.A(n_1837),
.B(n_1792),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1843),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1843),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1909),
.B(n_1829),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1881),
.Y(n_1916)
);

NAND2x1p5_ASAP7_75t_L g1917 ( 
.A(n_1912),
.B(n_1869),
.Y(n_1917)
);

AOI21xp33_ASAP7_75t_SL g1918 ( 
.A1(n_1886),
.A2(n_1870),
.B(n_1780),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1902),
.Y(n_1919)
);

OAI211xp5_ASAP7_75t_SL g1920 ( 
.A1(n_1912),
.A2(n_1815),
.B(n_1780),
.C(n_1841),
.Y(n_1920)
);

O2A1O1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1901),
.A2(n_1870),
.B(n_1825),
.C(n_1792),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1884),
.Y(n_1922)
);

INVxp67_ASAP7_75t_SL g1923 ( 
.A(n_1875),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_SL g1924 ( 
.A1(n_1875),
.A2(n_1759),
.B1(n_1797),
.B2(n_1795),
.Y(n_1924)
);

AOI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1876),
.A2(n_1839),
.B1(n_1797),
.B2(n_1800),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1893),
.B(n_1860),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1906),
.B(n_1845),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_R g1928 ( 
.A(n_1902),
.B(n_1625),
.Y(n_1928)
);

OAI21xp33_ASAP7_75t_L g1929 ( 
.A1(n_1887),
.A2(n_1861),
.B(n_1831),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1873),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1902),
.B(n_1826),
.Y(n_1931)
);

AOI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1876),
.A2(n_1800),
.B1(n_1795),
.B2(n_1844),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1911),
.B(n_1898),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1898),
.B(n_1826),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1873),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1878),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1906),
.B(n_1865),
.Y(n_1937)
);

AOI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1891),
.A2(n_1800),
.B1(n_1864),
.B2(n_1844),
.Y(n_1938)
);

OAI21xp5_ASAP7_75t_SL g1939 ( 
.A1(n_1888),
.A2(n_1832),
.B(n_1831),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1878),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1910),
.B(n_1872),
.Y(n_1941)
);

INVxp67_ASAP7_75t_L g1942 ( 
.A(n_1896),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1874),
.B(n_1832),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1923),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1919),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1916),
.B(n_1899),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1917),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1916),
.B(n_1899),
.Y(n_1948)
);

NOR2xp67_ASAP7_75t_L g1949 ( 
.A(n_1918),
.B(n_1877),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1937),
.Y(n_1950)
);

AOI21xp33_ASAP7_75t_SL g1951 ( 
.A1(n_1917),
.A2(n_1886),
.B(n_1892),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1941),
.B(n_1910),
.Y(n_1952)
);

NOR2x1_ASAP7_75t_L g1953 ( 
.A(n_1920),
.B(n_1899),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1930),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1928),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1935),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1922),
.B(n_1884),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1933),
.B(n_1926),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1936),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1940),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1915),
.Y(n_1961)
);

NAND2x1_ASAP7_75t_SL g1962 ( 
.A(n_1932),
.B(n_1891),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1942),
.B(n_1896),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1934),
.B(n_1889),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1931),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1927),
.B(n_1889),
.Y(n_1966)
);

NAND4xp25_ASAP7_75t_L g1967 ( 
.A(n_1946),
.B(n_1915),
.C(n_1921),
.D(n_1943),
.Y(n_1967)
);

AOI21xp33_ASAP7_75t_L g1968 ( 
.A1(n_1944),
.A2(n_1938),
.B(n_1914),
.Y(n_1968)
);

AOI211xp5_ASAP7_75t_L g1969 ( 
.A1(n_1951),
.A2(n_1929),
.B(n_1939),
.C(n_1905),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1961),
.A2(n_1925),
.B1(n_1924),
.B2(n_1882),
.C(n_1894),
.Y(n_1970)
);

AOI211xp5_ASAP7_75t_L g1971 ( 
.A1(n_1949),
.A2(n_1946),
.B(n_1948),
.C(n_1955),
.Y(n_1971)
);

AOI222xp33_ASAP7_75t_L g1972 ( 
.A1(n_1962),
.A2(n_1903),
.B1(n_1913),
.B2(n_1914),
.C1(n_1864),
.C2(n_1895),
.Y(n_1972)
);

OAI211xp5_ASAP7_75t_SL g1973 ( 
.A1(n_1953),
.A2(n_1908),
.B(n_1880),
.C(n_1883),
.Y(n_1973)
);

NAND4xp25_ASAP7_75t_L g1974 ( 
.A(n_1948),
.B(n_1903),
.C(n_1880),
.D(n_1883),
.Y(n_1974)
);

AOI211xp5_ASAP7_75t_L g1975 ( 
.A1(n_1965),
.A2(n_1950),
.B(n_1958),
.C(n_1947),
.Y(n_1975)
);

NAND3xp33_ASAP7_75t_L g1976 ( 
.A(n_1963),
.B(n_1903),
.C(n_1897),
.Y(n_1976)
);

NOR2x1_ASAP7_75t_L g1977 ( 
.A(n_1945),
.B(n_1897),
.Y(n_1977)
);

AOI221x1_ASAP7_75t_L g1978 ( 
.A1(n_1963),
.A2(n_1885),
.B1(n_1879),
.B2(n_1900),
.C(n_1904),
.Y(n_1978)
);

AOI211xp5_ASAP7_75t_L g1979 ( 
.A1(n_1947),
.A2(n_1885),
.B(n_1900),
.C(n_1879),
.Y(n_1979)
);

NAND3xp33_ASAP7_75t_L g1980 ( 
.A(n_1954),
.B(n_1904),
.C(n_1890),
.Y(n_1980)
);

AOI221xp5_ASAP7_75t_L g1981 ( 
.A1(n_1956),
.A2(n_1914),
.B1(n_1913),
.B2(n_1759),
.C(n_1760),
.Y(n_1981)
);

AO22x2_ASAP7_75t_L g1982 ( 
.A1(n_1976),
.A2(n_1960),
.B1(n_1959),
.B2(n_1966),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1977),
.Y(n_1983)
);

NOR2x1_ASAP7_75t_L g1984 ( 
.A(n_1973),
.B(n_1957),
.Y(n_1984)
);

NOR3xp33_ASAP7_75t_L g1985 ( 
.A(n_1971),
.B(n_1964),
.C(n_1913),
.Y(n_1985)
);

NAND3xp33_ASAP7_75t_SL g1986 ( 
.A(n_1972),
.B(n_1952),
.C(n_1964),
.Y(n_1986)
);

OA21x2_ASAP7_75t_L g1987 ( 
.A1(n_1978),
.A2(n_1952),
.B(n_1867),
.Y(n_1987)
);

NOR2xp67_ASAP7_75t_L g1988 ( 
.A(n_1974),
.B(n_1890),
.Y(n_1988)
);

NAND5xp2_ASAP7_75t_L g1989 ( 
.A(n_1969),
.B(n_1726),
.C(n_1727),
.D(n_1853),
.E(n_1863),
.Y(n_1989)
);

NOR3xp33_ASAP7_75t_L g1990 ( 
.A(n_1975),
.B(n_1907),
.C(n_1815),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1980),
.Y(n_1991)
);

NAND3xp33_ASAP7_75t_L g1992 ( 
.A(n_1968),
.B(n_1907),
.C(n_1867),
.Y(n_1992)
);

XNOR2x1_ASAP7_75t_L g1993 ( 
.A(n_1967),
.B(n_1679),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1979),
.B(n_1865),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1989),
.B(n_1970),
.Y(n_1995)
);

NAND3xp33_ASAP7_75t_L g1996 ( 
.A(n_1983),
.B(n_1981),
.C(n_1759),
.Y(n_1996)
);

NOR4xp25_ASAP7_75t_SL g1997 ( 
.A(n_1991),
.B(n_1868),
.C(n_1850),
.D(n_1793),
.Y(n_1997)
);

NOR3x1_ASAP7_75t_L g1998 ( 
.A(n_1986),
.B(n_1862),
.C(n_1858),
.Y(n_1998)
);

BUFx2_ASAP7_75t_L g1999 ( 
.A(n_1982),
.Y(n_1999)
);

AOI221xp5_ASAP7_75t_L g2000 ( 
.A1(n_1982),
.A2(n_1759),
.B1(n_1760),
.B2(n_1751),
.C(n_1805),
.Y(n_2000)
);

NOR4xp25_ASAP7_75t_L g2001 ( 
.A(n_1992),
.B(n_1815),
.C(n_1852),
.D(n_1805),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1999),
.A2(n_1984),
.B1(n_1985),
.B2(n_1988),
.Y(n_2002)
);

AOI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1995),
.A2(n_1987),
.B1(n_1990),
.B2(n_1993),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1998),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1996),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_2001),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_2000),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1997),
.Y(n_2008)
);

AOI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1999),
.A2(n_1994),
.B1(n_1805),
.B2(n_1815),
.Y(n_2009)
);

AND3x4_ASAP7_75t_L g2010 ( 
.A(n_2002),
.B(n_1635),
.C(n_1625),
.Y(n_2010)
);

AND3x4_ASAP7_75t_L g2011 ( 
.A(n_2003),
.B(n_1647),
.C(n_1635),
.Y(n_2011)
);

NOR3xp33_ASAP7_75t_L g2012 ( 
.A(n_2008),
.B(n_1871),
.C(n_1760),
.Y(n_2012)
);

AOI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_2007),
.A2(n_1759),
.B1(n_1751),
.B2(n_1740),
.Y(n_2013)
);

NOR2x1_ASAP7_75t_L g2014 ( 
.A(n_2006),
.B(n_1853),
.Y(n_2014)
);

BUFx2_ASAP7_75t_L g2015 ( 
.A(n_2005),
.Y(n_2015)
);

NAND3x1_ASAP7_75t_L g2016 ( 
.A(n_2014),
.B(n_2004),
.C(n_2009),
.Y(n_2016)
);

NAND4xp75_ASAP7_75t_L g2017 ( 
.A(n_2015),
.B(n_1650),
.C(n_1757),
.D(n_1863),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_2012),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_2011),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_2016),
.Y(n_2020)
);

INVxp67_ASAP7_75t_L g2021 ( 
.A(n_2018),
.Y(n_2021)
);

AOI321xp33_ASAP7_75t_L g2022 ( 
.A1(n_2020),
.A2(n_2019),
.A3(n_2010),
.B1(n_2013),
.B2(n_2017),
.C(n_1755),
.Y(n_2022)
);

AOI21xp33_ASAP7_75t_SL g2023 ( 
.A1(n_2022),
.A2(n_2021),
.B(n_1871),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_2022),
.B(n_1809),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_2023),
.B(n_1842),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2024),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_2025),
.B(n_2026),
.Y(n_2027)
);

AOI22xp5_ASAP7_75t_SL g2028 ( 
.A1(n_2025),
.A2(n_1842),
.B1(n_1872),
.B2(n_1647),
.Y(n_2028)
);

AOI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_2027),
.A2(n_1812),
.B1(n_1809),
.B2(n_1810),
.Y(n_2029)
);

AOI22xp5_ASAP7_75t_SL g2030 ( 
.A1(n_2029),
.A2(n_2028),
.B1(n_1743),
.B2(n_1775),
.Y(n_2030)
);

AOI221xp5_ASAP7_75t_L g2031 ( 
.A1(n_2030),
.A2(n_1751),
.B1(n_1812),
.B2(n_1810),
.C(n_1732),
.Y(n_2031)
);

AOI211xp5_ASAP7_75t_L g2032 ( 
.A1(n_2031),
.A2(n_1743),
.B(n_1757),
.C(n_1736),
.Y(n_2032)
);


endmodule