module fake_jpeg_13153_n_511 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_511);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_511;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_SL g41 ( 
.A(n_15),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_13),
.B(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_57),
.B(n_63),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g165 ( 
.A(n_58),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_60),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_61),
.Y(n_191)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_62),
.Y(n_178)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_64),
.B(n_66),
.Y(n_141)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_65),
.Y(n_174)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_67),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_69),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_17),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_70),
.B(n_83),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_71),
.B(n_74),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_75),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_18),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_76),
.B(n_77),
.Y(n_173)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_80),
.B(n_88),
.Y(n_179)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_82),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_15),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_84),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_86),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_29),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_90),
.B(n_91),
.Y(n_187)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

BUFx24_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

BUFx12f_ASAP7_75t_SL g145 ( 
.A(n_93),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_22),
.B(n_0),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_94),
.B(n_95),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_22),
.A2(n_1),
.B(n_2),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_97),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_40),
.B(n_2),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_98),
.B(n_99),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_24),
.B(n_2),
.Y(n_99)
);

BUFx16f_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_101),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_34),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_103),
.B(n_105),
.Y(n_201)
);

INVx11_ASAP7_75t_SL g104 ( 
.A(n_43),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_104),
.Y(n_131)
);

BUFx4f_ASAP7_75t_SL g105 ( 
.A(n_34),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

CKINVDCx9p33_ASAP7_75t_R g107 ( 
.A(n_34),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_34),
.Y(n_108)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_31),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_112),
.Y(n_160)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_54),
.Y(n_126)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_116),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_24),
.B(n_4),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_31),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_28),
.B(n_4),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_120),
.B(n_121),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_34),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_122),
.B(n_54),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_72),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_123),
.A2(n_127),
.B1(n_130),
.B2(n_133),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_126),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_75),
.A2(n_47),
.B1(n_56),
.B2(n_38),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_78),
.A2(n_53),
.B1(n_56),
.B2(n_49),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_79),
.A2(n_38),
.B1(n_51),
.B2(n_49),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_54),
.B1(n_53),
.B2(n_50),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_140),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_68),
.A2(n_54),
.B1(n_50),
.B2(n_51),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_61),
.A2(n_50),
.B1(n_51),
.B2(n_56),
.Y(n_137)
);

OA22x2_ASAP7_75t_SL g139 ( 
.A1(n_93),
.A2(n_50),
.B1(n_42),
.B2(n_45),
.Y(n_139)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_139),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_45),
.B1(n_38),
.B2(n_50),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_89),
.A2(n_45),
.B1(n_32),
.B2(n_28),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_142),
.A2(n_146),
.B1(n_151),
.B2(n_156),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_93),
.A2(n_42),
.B1(n_48),
.B2(n_44),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_96),
.A2(n_52),
.B1(n_32),
.B2(n_48),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_150),
.B(n_153),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_98),
.A2(n_52),
.B1(n_42),
.B2(n_6),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_84),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_92),
.A2(n_15),
.B1(n_7),
.B2(n_9),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_157),
.B(n_184),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_113),
.A2(n_5),
.B1(n_10),
.B2(n_13),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_158),
.A2(n_168),
.B1(n_169),
.B2(n_171),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_73),
.A2(n_5),
.B1(n_13),
.B2(n_14),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_163),
.B(n_175),
.Y(n_260)
);

HAxp5_ASAP7_75t_SL g167 ( 
.A(n_65),
.B(n_13),
.CON(n_167),
.SN(n_167)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_167),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_114),
.A2(n_14),
.B1(n_15),
.B2(n_112),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_62),
.A2(n_106),
.B1(n_117),
.B2(n_101),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_86),
.A2(n_97),
.B1(n_102),
.B2(n_65),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_102),
.A2(n_85),
.B1(n_108),
.B2(n_69),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_172),
.A2(n_177),
.B1(n_185),
.B2(n_195),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_60),
.A2(n_58),
.B1(n_105),
.B2(n_59),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_85),
.A2(n_108),
.B1(n_59),
.B2(n_69),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_104),
.A2(n_58),
.B1(n_105),
.B2(n_100),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_180),
.A2(n_148),
.B(n_155),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_100),
.A2(n_55),
.B1(n_82),
.B2(n_81),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_67),
.A2(n_81),
.B1(n_82),
.B2(n_111),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_192),
.B(n_140),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_70),
.A2(n_83),
.B1(n_90),
.B2(n_55),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_148),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_107),
.A2(n_54),
.B1(n_53),
.B2(n_21),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_107),
.A2(n_54),
.B1(n_53),
.B2(n_21),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_203),
.Y(n_226)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_205),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_187),
.B(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_206),
.B(n_216),
.Y(n_299)
);

BUFx4f_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_207),
.Y(n_280)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_128),
.Y(n_209)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_212),
.Y(n_275)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_141),
.Y(n_214)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_214),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_129),
.C(n_183),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_215),
.B(n_238),
.C(n_249),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_183),
.B(n_197),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_217),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_218),
.B(n_219),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_186),
.B(n_188),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_220),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g222 ( 
.A(n_129),
.B(n_192),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_224),
.Y(n_273)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_144),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_225),
.B(n_246),
.Y(n_289)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_159),
.Y(n_228)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_228),
.Y(n_298)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_159),
.Y(n_230)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_230),
.Y(n_301)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_152),
.Y(n_231)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_231),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_201),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_232),
.B(n_234),
.Y(n_276)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_233),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_160),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_235),
.B(n_242),
.Y(n_284)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

INVx6_ASAP7_75t_SL g302 ( 
.A(n_236),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_237),
.A2(n_262),
.B1(n_268),
.B2(n_270),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_138),
.B(n_149),
.C(n_202),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_138),
.B(n_149),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_241),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_142),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_160),
.B(n_165),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_243),
.B(n_251),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_165),
.B(n_131),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_244),
.B(n_245),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_165),
.B(n_131),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_185),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_143),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_145),
.B(n_166),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_248),
.B(n_250),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_170),
.B(n_178),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_165),
.B(n_178),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_170),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_145),
.B(n_204),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_252),
.B(n_253),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_200),
.B(n_204),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_161),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_254),
.B(n_258),
.Y(n_305)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_132),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_174),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_143),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_256),
.Y(n_300)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_161),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_162),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_259),
.B(n_263),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_162),
.B(n_164),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_125),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_164),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_200),
.B(n_134),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_264),
.B(n_266),
.Y(n_319)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_132),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_267),
.Y(n_306)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_181),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_213),
.A2(n_133),
.B1(n_127),
.B2(n_123),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_274),
.A2(n_241),
.B1(n_269),
.B2(n_265),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_SL g277 ( 
.A1(n_229),
.A2(n_167),
.B(n_139),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_277),
.A2(n_285),
.B(n_256),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_282),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_224),
.A2(n_180),
.B(n_139),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_287),
.B(n_294),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_213),
.A2(n_125),
.B1(n_189),
.B2(n_174),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_288),
.A2(n_303),
.B1(n_226),
.B2(n_271),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_222),
.B(n_176),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_291),
.B(n_297),
.C(n_309),
.Y(n_341)
);

AO22x1_ASAP7_75t_SL g294 ( 
.A1(n_243),
.A2(n_189),
.B1(n_191),
.B2(n_154),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_222),
.B(n_154),
.C(n_176),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_221),
.A2(n_191),
.B1(n_147),
.B2(n_134),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_234),
.B(n_147),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_304),
.B(n_307),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_239),
.B(n_181),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_215),
.B(n_238),
.C(n_243),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_255),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_240),
.A2(n_271),
.B(n_229),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_249),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_260),
.B(n_208),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_249),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_276),
.B(n_260),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_320),
.B(n_325),
.Y(n_387)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_305),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_330),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_286),
.A2(n_221),
.B1(n_208),
.B2(n_227),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_324),
.A2(n_331),
.B1(n_332),
.B2(n_273),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_251),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_276),
.B(n_257),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_326),
.B(n_328),
.Y(n_386)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_327),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_205),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_314),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_286),
.A2(n_261),
.B1(n_256),
.B2(n_231),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_289),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_333),
.B(n_335),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_334),
.B(n_339),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_302),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_302),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_336),
.B(n_347),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_337),
.A2(n_343),
.B(n_282),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_309),
.B(n_296),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_296),
.C(n_291),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_273),
.B(n_207),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_299),
.B(n_212),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_342),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_247),
.Y(n_342)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_345),
.Y(n_377)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_301),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_350),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_319),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_283),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_348),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_217),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_313),
.A2(n_220),
.B1(n_223),
.B2(n_258),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_351),
.A2(n_356),
.B1(n_300),
.B2(n_280),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_303),
.A2(n_259),
.B1(n_262),
.B2(n_211),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_352),
.Y(n_371)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_287),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_357),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_282),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_358),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_273),
.A2(n_237),
.B1(n_210),
.B2(n_236),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_307),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_312),
.B(n_207),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_363),
.B(n_367),
.C(n_373),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_364),
.A2(n_374),
.B1(n_344),
.B2(n_322),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_316),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_342),
.C(n_329),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_328),
.Y(n_366)
);

INVx13_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_297),
.C(n_304),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_341),
.B(n_290),
.C(n_292),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_324),
.A2(n_290),
.B1(n_288),
.B2(n_294),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_334),
.B(n_290),
.C(n_293),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_378),
.C(n_380),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_294),
.C(n_285),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_357),
.C(n_349),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_326),
.A2(n_306),
.B1(n_280),
.B2(n_281),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_384),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_278),
.C(n_272),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_337),
.C(n_325),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_306),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_390),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_333),
.Y(n_389)
);

NAND3xp33_ASAP7_75t_L g403 ( 
.A(n_389),
.B(n_379),
.C(n_320),
.Y(n_403)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_369),
.Y(n_391)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_391),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_370),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_392),
.B(n_403),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_393),
.A2(n_331),
.B1(n_378),
.B2(n_390),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_347),
.Y(n_394)
);

INVxp33_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_323),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_396),
.B(n_400),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_375),
.Y(n_397)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_399),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_362),
.B(n_340),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_359),
.A2(n_336),
.B1(n_335),
.B2(n_330),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_402),
.A2(n_381),
.B(n_351),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_368),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_404),
.B(n_410),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_365),
.B(n_337),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_409),
.C(n_411),
.Y(n_422)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_361),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_406),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_375),
.B(n_332),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_363),
.B(n_343),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_383),
.B(n_355),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_412),
.B(n_413),
.Y(n_438)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_372),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_367),
.B(n_344),
.C(n_350),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_414),
.B(n_417),
.C(n_388),
.Y(n_425)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_372),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_415),
.A2(n_416),
.B1(n_300),
.B2(n_377),
.Y(n_434)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_377),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_410),
.A2(n_364),
.B1(n_374),
.B2(n_359),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_418),
.A2(n_439),
.B1(n_408),
.B2(n_397),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_405),
.B(n_388),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_419),
.B(n_414),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_420),
.A2(n_423),
.B1(n_429),
.B2(n_409),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_393),
.A2(n_408),
.B1(n_395),
.B2(n_404),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_425),
.B(n_426),
.C(n_435),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_373),
.C(n_380),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_408),
.A2(n_385),
.B1(n_366),
.B2(n_371),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_346),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_376),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_436),
.A2(n_318),
.B(n_348),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_382),
.C(n_386),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_407),
.C(n_399),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_395),
.A2(n_371),
.B1(n_368),
.B2(n_360),
.Y(n_439)
);

AOI322xp5_ASAP7_75t_L g440 ( 
.A1(n_401),
.A2(n_360),
.A3(n_361),
.B1(n_348),
.B2(n_354),
.C1(n_356),
.C2(n_327),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_295),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_441),
.A2(n_443),
.B1(n_451),
.B2(n_434),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_442),
.B(n_435),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_418),
.A2(n_392),
.B1(n_417),
.B2(n_401),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_420),
.A2(n_412),
.B1(n_391),
.B2(n_413),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_444),
.A2(n_445),
.B1(n_447),
.B2(n_430),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_423),
.A2(n_429),
.B1(n_430),
.B2(n_424),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_448),
.B(n_450),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_438),
.B(n_400),
.Y(n_449)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_449),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_407),
.C(n_416),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_439),
.A2(n_415),
.B1(n_406),
.B2(n_345),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_438),
.Y(n_452)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_452),
.Y(n_464)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_424),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_453),
.A2(n_455),
.B1(n_458),
.B2(n_433),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_454),
.A2(n_456),
.B(n_457),
.Y(n_462)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_428),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_436),
.A2(n_321),
.B(n_281),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_446),
.B(n_437),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_461),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_425),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_443),
.B(n_419),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_463),
.B(n_466),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_448),
.B(n_421),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_465),
.B(n_468),
.Y(n_473)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_449),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_470),
.B(n_444),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_447),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_422),
.C(n_442),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_472),
.B(n_441),
.Y(n_476)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_474),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_475),
.A2(n_477),
.B(n_478),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_476),
.A2(n_467),
.B1(n_462),
.B2(n_463),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_421),
.C(n_422),
.Y(n_477)
);

A2O1A1O1Ixp25_ASAP7_75t_L g478 ( 
.A1(n_469),
.A2(n_445),
.B(n_453),
.C(n_452),
.D(n_457),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_431),
.C(n_458),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g485 ( 
.A(n_480),
.B(n_471),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_460),
.B(n_427),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_483),
.A2(n_427),
.B1(n_464),
.B2(n_472),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_484),
.B(n_489),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_SL g497 ( 
.A(n_485),
.B(n_492),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_482),
.B(n_464),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_488),
.Y(n_493)
);

BUFx4f_ASAP7_75t_SL g490 ( 
.A(n_478),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_490),
.B(n_476),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_473),
.B(n_451),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_456),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_466),
.Y(n_492)
);

A2O1A1Ixp33_ASAP7_75t_SL g495 ( 
.A1(n_490),
.A2(n_488),
.B(n_491),
.C(n_462),
.Y(n_495)
);

NAND3xp33_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_496),
.C(n_498),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_487),
.B(n_479),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_499),
.B(n_490),
.Y(n_502)
);

BUFx24_ASAP7_75t_SL g501 ( 
.A(n_494),
.Y(n_501)
);

AOI322xp5_ASAP7_75t_L g505 ( 
.A1(n_501),
.A2(n_502),
.A3(n_495),
.B1(n_455),
.B2(n_433),
.C1(n_428),
.C2(n_432),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_486),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_503),
.B(n_504),
.C(n_278),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_497),
.A2(n_475),
.B(n_432),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_505),
.B(n_506),
.Y(n_508)
);

AOI322xp5_ASAP7_75t_L g506 ( 
.A1(n_500),
.A2(n_454),
.A3(n_492),
.B1(n_481),
.B2(n_283),
.C1(n_279),
.C2(n_311),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_507),
.A2(n_272),
.B(n_295),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_509),
.A2(n_275),
.B1(n_317),
.B2(n_315),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_510),
.B(n_508),
.Y(n_511)
);


endmodule