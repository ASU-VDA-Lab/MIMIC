module real_jpeg_3697_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_286;
wire n_288;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_290;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_244;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_2),
.A2(n_21),
.B1(n_22),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_2),
.A2(n_48),
.B1(n_59),
.B2(n_60),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_48),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_2),
.A2(n_48),
.B1(n_69),
.B2(n_70),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_50),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_3),
.A2(n_50),
.B1(n_59),
.B2(n_60),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_3),
.A2(n_50),
.B1(n_69),
.B2(n_70),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_3),
.B(n_29),
.C(n_33),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_3),
.B(n_31),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_3),
.B(n_56),
.C(n_60),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_3),
.B(n_90),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_3),
.B(n_67),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_3),
.B(n_68),
.C(n_70),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_3),
.B(n_62),
.Y(n_232)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_6),
.A2(n_21),
.B1(n_22),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_39),
.B1(n_69),
.B2(n_70),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_6),
.A2(n_39),
.B1(n_59),
.B2(n_60),
.Y(n_112)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_10),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_15),
.B(n_291),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_11),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_12),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_12),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_12),
.A2(n_25),
.B1(n_59),
.B2(n_60),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_12),
.A2(n_25),
.B1(n_69),
.B2(n_70),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_41),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_40),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_26),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_20),
.A2(n_27),
.B1(n_36),
.B2(n_38),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_29),
.Y(n_30)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_22),
.B(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_26),
.B(n_49),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_36),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_28),
.A2(n_31),
.B1(n_46),
.B2(n_49),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_28),
.B(n_49),
.Y(n_78)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_32),
.A2(n_33),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_33),
.B(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_36),
.A2(n_38),
.B(n_78),
.Y(n_77)
);

OA21x2_ASAP7_75t_L g127 ( 
.A1(n_36),
.A2(n_47),
.B(n_78),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_37),
.B(n_43),
.Y(n_290)
);

AO21x1_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_79),
.B(n_290),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_75),
.C(n_77),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_44),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.C(n_64),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_45),
.A2(n_100),
.B1(n_104),
.B2(n_105),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_45),
.A2(n_105),
.B1(n_142),
.B2(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_45),
.B(n_142),
.C(n_152),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_45),
.A2(n_105),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_51),
.A2(n_64),
.B1(n_262),
.B2(n_279),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_51),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_63),
.Y(n_51)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_52),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_53),
.A2(n_62),
.B1(n_101),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_54),
.B(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_54),
.A2(n_58),
.B(n_103),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

AOI22x1_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_58),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_60),
.B1(n_68),
.B2(n_71),
.Y(n_73)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_60),
.B(n_225),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AO21x1_ASAP7_75t_L g100 ( 
.A1(n_62),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_64),
.A2(n_262),
.B1(n_263),
.B2(n_266),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_64),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_64),
.B(n_127),
.C(n_263),
.Y(n_280)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_74),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_72),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_66),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_66),
.A2(n_72),
.B1(n_96),
.B2(n_97),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_66),
.A2(n_72),
.B(n_97),
.Y(n_168)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_67),
.A2(n_74),
.B1(n_115),
.B2(n_141),
.Y(n_140)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_67)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_70),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_75),
.B(n_77),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_285),
.B(n_289),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_256),
.B(n_282),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_146),
.B(n_255),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_128),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_83),
.B(n_128),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_106),
.C(n_117),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_84),
.B(n_106),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_98),
.B2(n_99),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_100),
.C(n_105),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_94),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_87),
.A2(n_94),
.B1(n_95),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_87),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_89),
.A2(n_90),
.B1(n_122),
.B2(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_92),
.B(n_121),
.Y(n_120)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_92),
.A2(n_121),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_94),
.A2(n_95),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_94),
.A2(n_95),
.B1(n_205),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_95),
.B(n_200),
.C(n_205),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_95),
.B(n_157),
.C(n_232),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_100),
.B(n_126),
.C(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_100),
.A2(n_104),
.B1(n_168),
.B2(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_100),
.A2(n_104),
.B1(n_123),
.B2(n_124),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_100),
.B(n_123),
.C(n_239),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_102),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B1(n_111),
.B2(n_116),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_111),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_116),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_109),
.B(n_122),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_116),
.A2(n_132),
.B(n_137),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_117),
.B(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.C(n_126),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_118),
.A2(n_119),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_120),
.A2(n_123),
.B1(n_124),
.B2(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_120),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_123),
.A2(n_124),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_123),
.B(n_226),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_126),
.A2(n_127),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_126),
.A2(n_127),
.B1(n_261),
.B2(n_267),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_126),
.A2(n_127),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_127),
.B(n_276),
.C(n_280),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_145),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_138),
.B2(n_139),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_131),
.B(n_138),
.C(n_145),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_136),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_142),
.B(n_144),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_142),
.Y(n_144)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_176),
.C(n_177),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_142),
.A2(n_160),
.B1(n_201),
.B2(n_204),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_144),
.A2(n_260),
.B1(n_268),
.B2(n_269),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_144),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_250),
.B(n_254),
.Y(n_146)
);

OAI211xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_179),
.B(n_193),
.C(n_249),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_169),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_169),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_161),
.B2(n_162),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_164),
.C(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_159),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_156),
.A2(n_157),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_157),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_157),
.B(n_220),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.C(n_175),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_175),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_177),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_SL g193 ( 
.A(n_180),
.B(n_194),
.C(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_181),
.B(n_182),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_183),
.B(n_185),
.C(n_191),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_190),
.B2(n_191),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_211),
.B(n_248),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_199),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_223),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_242),
.B(n_247),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_236),
.B(n_241),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_228),
.B(n_235),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_222),
.B(n_227),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_219),
.B(n_221),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_224),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_234),
.Y(n_235)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_246),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_252),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_272),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_271),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_271),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_270),
.Y(n_258)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_260),
.Y(n_269)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_263),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_269),
.C(n_270),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_281),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_281),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_288),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);


endmodule