module fake_jpeg_22413_n_87 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_87);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_87;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_2),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_27),
.Y(n_43)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_14),
.Y(n_41)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

OR2x2_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_19),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_29),
.B(n_18),
.Y(n_42)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_39),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_19),
.B1(n_21),
.B2(n_15),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.C(n_44),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_18),
.C(n_23),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_12),
.B1(n_20),
.B2(n_17),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_0),
.Y(n_47)
);

A2O1A1O1Ixp25_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_26),
.B(n_0),
.C(n_5),
.D(n_6),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_23),
.B1(n_20),
.B2(n_17),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_56),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_59),
.B(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_3),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_8),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_8),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_11),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_37),
.B1(n_34),
.B2(n_44),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_63),
.B1(n_69),
.B2(n_61),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_35),
.B1(n_46),
.B2(n_49),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_46),
.C(n_51),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_68),
.C(n_67),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_74),
.Y(n_76)
);

MAJx2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_65),
.C(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_73),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_79),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_76),
.B1(n_82),
.B2(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_83),
.B(n_81),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);


endmodule