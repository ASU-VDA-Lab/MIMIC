module fake_jpeg_4742_n_109 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx11_ASAP7_75t_SL g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx2_ASAP7_75t_SL g33 ( 
.A(n_22),
.Y(n_33)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_20),
.Y(n_24)
);

CKINVDCx6p67_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_13),
.B1(n_12),
.B2(n_14),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_13),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_18),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_23),
.A2(n_27),
.B1(n_12),
.B2(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_11),
.Y(n_42)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_19),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

NOR3xp33_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_37),
.C(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_54),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_34),
.C(n_37),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_26),
.B(n_24),
.Y(n_68)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_45),
.B1(n_52),
.B2(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_31),
.B1(n_29),
.B2(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_65),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_29),
.B(n_50),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_37),
.B(n_24),
.C(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_69),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_24),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_24),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_10),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_74),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_75),
.B1(n_65),
.B2(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI322xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_56),
.A3(n_19),
.B1(n_10),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_71),
.B(n_63),
.C(n_77),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_86),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_68),
.C(n_80),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_25),
.C(n_28),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_82),
.B1(n_67),
.B2(n_31),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_90),
.B1(n_87),
.B2(n_28),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_0),
.B(n_1),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_7),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_97),
.B1(n_96),
.B2(n_3),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_101),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_25),
.C(n_2),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_101),
.B(n_1),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_106),
.B(n_103),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_103),
.Y(n_109)
);


endmodule