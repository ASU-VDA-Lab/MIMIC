module fake_netlist_1_12442_n_673 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_673);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_673;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g83 ( .A(n_33), .Y(n_83) );
CKINVDCx14_ASAP7_75t_R g84 ( .A(n_79), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_78), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_23), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_53), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_32), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_43), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_51), .Y(n_90) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_66), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_28), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_67), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_80), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_3), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_41), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_63), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_82), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_49), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_44), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_52), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_4), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_69), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_58), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_56), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_48), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_74), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_54), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_3), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_9), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_60), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_36), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_6), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_73), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_42), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_61), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_27), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_26), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_55), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_13), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_34), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_85), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_109), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_106), .B(n_0), .Y(n_124) );
NOR2x1_ASAP7_75t_L g125 ( .A(n_87), .B(n_0), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_102), .B(n_1), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_94), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_96), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_120), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_109), .A2(n_2), .B1(n_5), .B2(n_6), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_91), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
INVx4_ASAP7_75t_L g134 ( .A(n_91), .Y(n_134) );
NOR2x1_ASAP7_75t_L g135 ( .A(n_97), .B(n_5), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_101), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_115), .Y(n_137) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_89), .A2(n_35), .B(n_81), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_91), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_113), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_89), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_134), .Y(n_143) );
INVx4_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_132), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_132), .Y(n_146) );
INVx2_ASAP7_75t_SL g147 ( .A(n_122), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_133), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_133), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_134), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_133), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_137), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_133), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_123), .B(n_86), .Y(n_154) );
AO22x2_ASAP7_75t_L g155 ( .A1(n_122), .A2(n_95), .B1(n_90), .B2(n_112), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_123), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_127), .B(n_103), .Y(n_157) );
INVx2_ASAP7_75t_SL g158 ( .A(n_127), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_130), .A2(n_113), .B1(n_95), .B2(n_110), .Y(n_159) );
AOI21x1_ASAP7_75t_L g160 ( .A1(n_128), .A2(n_99), .B(n_90), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_128), .B(n_84), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_134), .Y(n_162) );
AND3x2_ASAP7_75t_L g163 ( .A(n_126), .B(n_107), .C(n_111), .Y(n_163) );
INVx5_ASAP7_75t_L g164 ( .A(n_134), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_132), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_132), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_138), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_132), .Y(n_168) );
OAI22xp33_ASAP7_75t_L g169 ( .A1(n_130), .A2(n_121), .B1(n_119), .B2(n_86), .Y(n_169) );
AND2x6_ASAP7_75t_L g170 ( .A(n_125), .B(n_105), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_136), .A2(n_114), .B1(n_118), .B2(n_119), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_131), .A2(n_121), .B1(n_117), .B2(n_116), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_132), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_136), .B(n_88), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_129), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_124), .B(n_88), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_155), .A2(n_125), .B1(n_135), .B2(n_142), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_147), .B(n_92), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_161), .B(n_135), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_161), .B(n_92), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_159), .A2(n_141), .B1(n_142), .B2(n_129), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_155), .A2(n_138), .B1(n_93), .B2(n_108), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_155), .B(n_93), .Y(n_184) );
BUFx8_ASAP7_75t_L g185 ( .A(n_170), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_147), .B(n_158), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_147), .B(n_100), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_158), .B(n_100), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_144), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_155), .B(n_104), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
O2A1O1Ixp5_ASAP7_75t_L g193 ( .A1(n_144), .A2(n_112), .B(n_98), .C(n_99), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_163), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_144), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_158), .B(n_104), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_174), .B(n_108), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_175), .B(n_116), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_159), .A2(n_117), .B1(n_98), .B2(n_138), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_171), .B(n_91), .Y(n_200) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_152), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_176), .B(n_140), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_144), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_157), .B(n_140), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_163), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_175), .B(n_7), .Y(n_206) );
NOR2xp67_ASAP7_75t_L g207 ( .A(n_148), .B(n_38), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_148), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_169), .A2(n_140), .B1(n_139), .B2(n_11), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_154), .B(n_140), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_170), .B(n_140), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_149), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_170), .A2(n_140), .B1(n_139), .B2(n_11), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_172), .A2(n_139), .B1(n_10), .B2(n_12), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_167), .B(n_139), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_167), .A2(n_139), .B(n_37), .Y(n_216) );
NAND2x1_ASAP7_75t_L g217 ( .A(n_167), .B(n_139), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_167), .Y(n_218) );
AND3x1_ASAP7_75t_L g219 ( .A(n_172), .B(n_8), .C(n_10), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_177), .A2(n_149), .B1(n_151), .B2(n_153), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_180), .B(n_143), .Y(n_221) );
NOR2xp33_ASAP7_75t_SL g222 ( .A(n_201), .B(n_170), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_206), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_190), .Y(n_224) );
OR2x6_ASAP7_75t_L g225 ( .A(n_194), .B(n_151), .Y(n_225) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_216), .A2(n_160), .B(n_153), .Y(n_226) );
OAI21x1_ASAP7_75t_L g227 ( .A1(n_216), .A2(n_160), .B(n_146), .Y(n_227) );
AND2x6_ASAP7_75t_L g228 ( .A(n_177), .B(n_162), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_215), .A2(n_143), .B(n_150), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_193), .A2(n_143), .B(n_150), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_198), .B(n_170), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_189), .Y(n_232) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_199), .A2(n_173), .B(n_168), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_186), .A2(n_143), .B(n_150), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_214), .A2(n_150), .B(n_162), .C(n_170), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_185), .Y(n_236) );
NAND3xp33_ASAP7_75t_L g237 ( .A(n_183), .B(n_199), .C(n_178), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_198), .B(n_170), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_180), .B(n_170), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_192), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_181), .B(n_162), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_184), .B(n_162), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_206), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_208), .Y(n_244) );
AOI221xp5_ASAP7_75t_L g245 ( .A1(n_182), .A2(n_164), .B1(n_168), .B2(n_166), .C(n_165), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_208), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_185), .A2(n_164), .B1(n_168), .B2(n_166), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_184), .B(n_164), .Y(n_248) );
OR2x6_ASAP7_75t_L g249 ( .A(n_194), .B(n_12), .Y(n_249) );
OAI21xp33_ASAP7_75t_L g250 ( .A1(n_191), .A2(n_173), .B(n_166), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_191), .B(n_164), .Y(n_251) );
INVx4_ASAP7_75t_L g252 ( .A(n_192), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_196), .B(n_164), .Y(n_253) );
NOR2x1_ASAP7_75t_L g254 ( .A(n_225), .B(n_200), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_223), .B(n_212), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_232), .A2(n_203), .B(n_195), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_243), .B(n_182), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_244), .B(n_246), .Y(n_258) );
BUFx10_ASAP7_75t_L g259 ( .A(n_236), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_221), .B(n_205), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_221), .B(n_205), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_224), .B(n_197), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_239), .B(n_209), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_232), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_235), .A2(n_195), .B(n_189), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_252), .Y(n_266) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_249), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_234), .A2(n_217), .B(n_195), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_252), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_227), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_227), .A2(n_217), .B(n_189), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_SL g272 ( .A1(n_231), .A2(n_238), .B(n_245), .C(n_211), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_229), .A2(n_203), .B(n_218), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_230), .A2(n_203), .B(n_218), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_252), .B(n_219), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_237), .A2(n_214), .B1(n_213), .B2(n_219), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_257), .B(n_242), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_267), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_272), .A2(n_225), .B(n_226), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_258), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_267), .Y(n_281) );
AO31x2_ASAP7_75t_L g282 ( .A1(n_276), .A2(n_220), .A3(n_233), .B(n_204), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_258), .B(n_249), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_271), .A2(n_226), .B(n_247), .Y(n_284) );
INVx1_ASAP7_75t_SL g285 ( .A(n_262), .Y(n_285) );
A2O1A1Ixp33_ASAP7_75t_L g286 ( .A1(n_276), .A2(n_241), .B(n_250), .C(n_222), .Y(n_286) );
OR2x6_ASAP7_75t_L g287 ( .A(n_266), .B(n_225), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_271), .A2(n_226), .B(n_247), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_255), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_274), .A2(n_225), .B(n_253), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_264), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_268), .A2(n_218), .B(n_233), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_264), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_275), .A2(n_249), .B1(n_241), .B2(n_185), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_255), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_264), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_270), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_266), .Y(n_298) );
NOR2x1p5_ASAP7_75t_L g299 ( .A(n_275), .B(n_236), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_297), .Y(n_300) );
OR2x6_ASAP7_75t_L g301 ( .A(n_287), .B(n_254), .Y(n_301) );
OA21x2_ASAP7_75t_L g302 ( .A1(n_284), .A2(n_270), .B(n_265), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_291), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_291), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_297), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_297), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_291), .Y(n_307) );
INVx4_ASAP7_75t_SL g308 ( .A(n_287), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_293), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_293), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_293), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_296), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_296), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_289), .B(n_270), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_287), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_284), .Y(n_317) );
OA21x2_ASAP7_75t_L g318 ( .A1(n_288), .A2(n_265), .B(n_273), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_280), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_287), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_280), .Y(n_321) );
AOI33xp33_ASAP7_75t_L g322 ( .A1(n_285), .A2(n_213), .A3(n_269), .B1(n_15), .B2(n_16), .B3(n_17), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_298), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_298), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_295), .B(n_269), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_295), .B(n_256), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_282), .Y(n_327) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_292), .A2(n_263), .B(n_256), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_282), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_287), .Y(n_330) );
OR2x6_ASAP7_75t_L g331 ( .A(n_279), .B(n_254), .Y(n_331) );
OA21x2_ASAP7_75t_L g332 ( .A1(n_288), .A2(n_261), .B(n_260), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_282), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_308), .B(n_282), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_300), .B(n_282), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_300), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_304), .B(n_282), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_304), .B(n_283), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_313), .B(n_299), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_313), .B(n_277), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_300), .B(n_299), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_319), .B(n_294), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_314), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_315), .Y(n_344) );
OR2x6_ASAP7_75t_L g345 ( .A(n_330), .B(n_290), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_305), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_315), .B(n_286), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_305), .Y(n_348) );
OR2x6_ASAP7_75t_L g349 ( .A(n_330), .B(n_248), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_315), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_308), .B(n_316), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_305), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_306), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_306), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_306), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_308), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_303), .B(n_13), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_323), .B(n_278), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_319), .B(n_251), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_303), .B(n_14), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_323), .B(n_324), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_327), .B(n_14), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_321), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_330), .A2(n_281), .B1(n_262), .B2(n_259), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_321), .B(n_228), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_324), .B(n_15), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_307), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_307), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_309), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_309), .B(n_16), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_308), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_310), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_310), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_311), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_326), .B(n_228), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_311), .B(n_17), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_312), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_312), .B(n_18), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_314), .B(n_18), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_325), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_327), .B(n_19), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_314), .B(n_19), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_314), .B(n_20), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_317), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_329), .B(n_20), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_326), .B(n_228), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_326), .B(n_228), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_325), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_329), .B(n_21), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_317), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_308), .B(n_207), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_314), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_340), .B(n_338), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_362), .B(n_325), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_363), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_362), .B(n_316), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_340), .B(n_316), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_338), .B(n_316), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_346), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_346), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_361), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_368), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_358), .B(n_320), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_348), .Y(n_406) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_381), .B(n_301), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_368), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_339), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_389), .B(n_320), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_369), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_389), .B(n_320), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_369), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_373), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_389), .B(n_320), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_373), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_380), .B(n_388), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_356), .B(n_301), .Y(n_418) );
NOR2x1_ASAP7_75t_R g419 ( .A(n_356), .B(n_259), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_374), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_374), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_371), .B(n_301), .Y(n_422) );
INVx3_ASAP7_75t_L g423 ( .A(n_336), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_377), .Y(n_424) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_379), .B(n_382), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_336), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_336), .Y(n_427) );
AND2x4_ASAP7_75t_SL g428 ( .A(n_341), .B(n_259), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_367), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_367), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_344), .B(n_333), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_350), .B(n_333), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_350), .B(n_333), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_337), .B(n_328), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_337), .B(n_328), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_357), .B(n_301), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_360), .B(n_332), .Y(n_437) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_392), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_360), .B(n_332), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_367), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_372), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_371), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_372), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_381), .B(n_332), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_372), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_354), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_354), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_370), .B(n_332), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_385), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_354), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_352), .B(n_328), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_347), .B(n_328), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_366), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_352), .B(n_328), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_366), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_334), .B(n_322), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_353), .B(n_302), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_353), .B(n_302), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_342), .B(n_21), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_355), .B(n_302), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_347), .B(n_335), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_342), .B(n_331), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_379), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_383), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_395), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_446), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_442), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_393), .B(n_355), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_402), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_396), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_409), .B(n_334), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_446), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_394), .B(n_334), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_461), .B(n_335), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_437), .B(n_335), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_418), .B(n_351), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_404), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_461), .B(n_392), .Y(n_478) );
OAI33xp33_ASAP7_75t_L g479 ( .A1(n_456), .A2(n_359), .A3(n_365), .B1(n_375), .B2(n_387), .B3(n_386), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_408), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_411), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_456), .A2(n_364), .B1(n_349), .B2(n_376), .Y(n_482) );
AOI311xp33_ASAP7_75t_L g483 ( .A1(n_459), .A2(n_359), .A3(n_386), .B(n_387), .C(n_375), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_405), .B(n_343), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_459), .B(n_364), .Y(n_485) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_402), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_398), .B(n_403), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_413), .Y(n_488) );
NAND2xp33_ASAP7_75t_SL g489 ( .A(n_427), .B(n_376), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_414), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_416), .Y(n_491) );
OR2x6_ASAP7_75t_L g492 ( .A(n_425), .B(n_345), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_405), .B(n_343), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_426), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_400), .B(n_343), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_450), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_453), .B(n_378), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_455), .B(n_378), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_420), .Y(n_499) );
NOR2xp67_ASAP7_75t_L g500 ( .A(n_426), .B(n_383), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_418), .B(n_345), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_397), .B(n_410), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_421), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_423), .B(n_391), .Y(n_504) );
OR3x2_ASAP7_75t_L g505 ( .A(n_419), .B(n_322), .C(n_259), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_412), .B(n_349), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_422), .B(n_345), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_460), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_445), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_449), .B(n_349), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_424), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_464), .B(n_349), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_417), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_445), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_415), .B(n_345), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_431), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_431), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_430), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_447), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_433), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_436), .B(n_331), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_428), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_429), .Y(n_523) );
OR2x6_ASAP7_75t_L g524 ( .A(n_407), .B(n_331), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_433), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_423), .B(n_463), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_401), .Y(n_527) );
NOR3x1_ASAP7_75t_L g528 ( .A(n_452), .B(n_365), .C(n_210), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_440), .Y(n_529) );
INVx1_ASAP7_75t_SL g530 ( .A(n_399), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_441), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_443), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_462), .B(n_391), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_439), .B(n_331), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_432), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_406), .B(n_390), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_457), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_438), .Y(n_538) );
NAND5xp2_ASAP7_75t_L g539 ( .A(n_482), .B(n_462), .C(n_448), .D(n_435), .E(n_434), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_501), .B(n_422), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_468), .B(n_474), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_537), .B(n_434), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_473), .B(n_435), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_516), .B(n_451), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_502), .B(n_438), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_517), .B(n_454), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_465), .Y(n_547) );
NAND2x1_ASAP7_75t_L g548 ( .A(n_492), .B(n_438), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_520), .B(n_444), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_525), .B(n_458), .Y(n_550) );
OAI31xp33_ASAP7_75t_L g551 ( .A1(n_489), .A2(n_391), .A3(n_390), .B(n_384), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_470), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_467), .Y(n_553) );
O2A1O1Ixp33_ASAP7_75t_L g554 ( .A1(n_485), .A2(n_391), .B(n_202), .C(n_188), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_513), .B(n_390), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_475), .B(n_384), .Y(n_556) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_504), .A2(n_318), .B(n_302), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_475), .B(n_318), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_530), .B(n_318), .Y(n_559) );
INVxp67_ASAP7_75t_L g560 ( .A(n_527), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_535), .B(n_318), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_477), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_480), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_508), .B(n_318), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_471), .B(n_302), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_508), .B(n_207), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_487), .B(n_218), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_478), .B(n_22), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_481), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_488), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_490), .Y(n_571) );
OAI21xp33_ASAP7_75t_L g572 ( .A1(n_482), .A2(n_173), .B(n_146), .Y(n_572) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_485), .B(n_185), .C(n_145), .Y(n_573) );
BUFx2_ASAP7_75t_L g574 ( .A(n_494), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_469), .B(n_218), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_469), .B(n_218), .Y(n_576) );
INVxp67_ASAP7_75t_L g577 ( .A(n_527), .Y(n_577) );
NOR2x1p5_ASAP7_75t_L g578 ( .A(n_486), .B(n_240), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_522), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_509), .B(n_24), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_491), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g582 ( .A(n_483), .B(n_145), .C(n_187), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_514), .B(n_25), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_489), .A2(n_179), .B1(n_240), .B2(n_165), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_499), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_503), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g587 ( .A1(n_500), .A2(n_29), .B(n_30), .C(n_31), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_494), .B(n_514), .Y(n_588) );
OA21x2_ASAP7_75t_L g589 ( .A1(n_486), .A2(n_504), .B(n_472), .Y(n_589) );
NAND3xp33_ASAP7_75t_SL g590 ( .A(n_538), .B(n_39), .C(n_40), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_511), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_531), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_592), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_578), .A2(n_505), .B1(n_492), .B2(n_524), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_549), .B(n_526), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_556), .B(n_466), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_547), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_543), .B(n_472), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_552), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_562), .Y(n_600) );
OAI221xp5_ASAP7_75t_L g601 ( .A1(n_551), .A2(n_492), .B1(n_533), .B2(n_512), .C(n_510), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_572), .A2(n_533), .B1(n_479), .B2(n_515), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_544), .B(n_496), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_573), .A2(n_524), .B1(n_501), .B2(n_507), .Y(n_604) );
NAND2x1_ASAP7_75t_L g605 ( .A(n_589), .B(n_476), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_546), .B(n_532), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_572), .A2(n_479), .B1(n_507), .B2(n_501), .Y(n_607) );
NOR2x1p5_ASAP7_75t_L g608 ( .A(n_548), .B(n_590), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_546), .B(n_497), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_542), .B(n_498), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_563), .Y(n_611) );
OAI32xp33_ASAP7_75t_L g612 ( .A1(n_541), .A2(n_495), .A3(n_506), .B1(n_521), .B2(n_493), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_569), .Y(n_613) );
OAI22xp33_ASAP7_75t_L g614 ( .A1(n_579), .A2(n_524), .B1(n_529), .B2(n_523), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_574), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_570), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g617 ( .A1(n_573), .A2(n_523), .B1(n_529), .B2(n_534), .Y(n_617) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_554), .A2(n_536), .B(n_484), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_571), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_581), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_550), .B(n_518), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_558), .B(n_528), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_553), .A2(n_519), .B1(n_145), .B2(n_47), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_560), .B(n_577), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_540), .B(n_45), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_588), .A2(n_145), .B(n_50), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_612), .A2(n_539), .B1(n_591), .B2(n_586), .C(n_585), .Y(n_627) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_605), .A2(n_587), .B(n_539), .C(n_580), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_622), .A2(n_565), .B1(n_545), .B2(n_589), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_604), .A2(n_584), .B(n_582), .Y(n_630) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_604), .A2(n_568), .B(n_583), .Y(n_631) );
OAI221xp5_ASAP7_75t_L g632 ( .A1(n_601), .A2(n_559), .B1(n_555), .B2(n_561), .C(n_564), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_602), .B(n_564), .Y(n_633) );
AOI322xp5_ASAP7_75t_L g634 ( .A1(n_615), .A2(n_567), .A3(n_566), .B1(n_575), .B2(n_576), .C1(n_557), .C2(n_582), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_606), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_618), .A2(n_46), .B1(n_57), .B2(n_59), .C(n_62), .Y(n_636) );
OAI21xp33_ASAP7_75t_L g637 ( .A1(n_607), .A2(n_64), .B(n_65), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_617), .A2(n_68), .B(n_70), .Y(n_638) );
AOI22xp33_ASAP7_75t_SL g639 ( .A1(n_625), .A2(n_71), .B1(n_72), .B2(n_75), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_603), .Y(n_640) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_614), .A2(n_76), .B(n_77), .Y(n_641) );
AOI311xp33_ASAP7_75t_L g642 ( .A1(n_609), .A2(n_164), .A3(n_593), .B(n_620), .C(n_619), .Y(n_642) );
NAND3x1_ASAP7_75t_L g643 ( .A(n_624), .B(n_595), .C(n_611), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_621), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_625), .Y(n_645) );
AOI21xp33_ASAP7_75t_L g646 ( .A1(n_597), .A2(n_613), .B(n_616), .Y(n_646) );
AOI211xp5_ASAP7_75t_L g647 ( .A1(n_626), .A2(n_599), .B(n_600), .C(n_610), .Y(n_647) );
OA22x2_ASAP7_75t_L g648 ( .A1(n_598), .A2(n_623), .B1(n_608), .B2(n_596), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_612), .A2(n_618), .B1(n_622), .B2(n_601), .C(n_539), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_605), .A2(n_594), .B(n_604), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_605), .A2(n_594), .B(n_604), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_651), .B(n_650), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_642), .B(n_649), .C(n_634), .Y(n_653) );
NOR3xp33_ASAP7_75t_L g654 ( .A(n_630), .B(n_636), .C(n_637), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_627), .A2(n_632), .B1(n_633), .B2(n_646), .C(n_631), .Y(n_655) );
BUFx12f_ASAP7_75t_L g656 ( .A(n_639), .Y(n_656) );
AND3x2_ASAP7_75t_L g657 ( .A(n_647), .B(n_643), .C(n_640), .Y(n_657) );
NOR4xp25_ASAP7_75t_L g658 ( .A(n_653), .B(n_652), .C(n_655), .D(n_657), .Y(n_658) );
NOR3xp33_ASAP7_75t_L g659 ( .A(n_654), .B(n_628), .C(n_641), .Y(n_659) );
BUFx2_ASAP7_75t_L g660 ( .A(n_656), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_652), .B(n_635), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_660), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_658), .B(n_629), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_661), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_662), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_664), .B(n_659), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_665), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_666), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_667), .A2(n_663), .B(n_648), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_669), .B(n_668), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_670), .B(n_668), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_671), .B(n_645), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_672), .A2(n_638), .B(n_644), .Y(n_673) );
endmodule