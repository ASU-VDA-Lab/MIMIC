module real_aes_3726_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_635;
wire n_503;
wire n_357;
wire n_386;
wire n_673;
wire n_905;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_962;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_947;
wire n_142;
wire n_561;
wire n_970;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_954;
wire n_296;
wire n_702;
wire n_969;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_972;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_926;
wire n_922;
wire n_149;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_134;
wire n_946;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_646;
wire n_650;
wire n_105;
wire n_743;
wire n_710;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_823;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
INVx1_ASAP7_75t_L g676 ( .A(n_0), .Y(n_676) );
OAI22x1_ASAP7_75t_SL g112 ( .A1(n_1), .A2(n_53), .B1(n_113), .B2(n_114), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_1), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_2), .A2(n_22), .B1(n_126), .B2(n_129), .Y(n_125) );
INVx1_ASAP7_75t_L g270 ( .A(n_3), .Y(n_270) );
INVx2_ASAP7_75t_L g296 ( .A(n_4), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_5), .B(n_575), .Y(n_632) );
INVx1_ASAP7_75t_SL g246 ( .A(n_6), .Y(n_246) );
INVxp67_ASAP7_75t_L g542 ( .A(n_7), .Y(n_542) );
INVx1_ASAP7_75t_L g561 ( .A(n_7), .Y(n_561) );
INVx1_ASAP7_75t_L g944 ( .A(n_7), .Y(n_944) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_8), .B(n_203), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_9), .A2(n_43), .B1(n_574), .B2(n_619), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_10), .A2(n_49), .B1(n_190), .B2(n_593), .Y(n_699) );
XOR2xp5_ASAP7_75t_R g946 ( .A(n_11), .B(n_947), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_12), .A2(n_70), .B1(n_654), .B2(n_655), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_13), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_14), .B(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g671 ( .A(n_15), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_16), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_17), .A2(n_105), .B1(n_965), .B2(n_968), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_18), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g534 ( .A(n_18), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_19), .A2(n_58), .B1(n_202), .B2(n_203), .Y(n_201) );
INVx1_ASAP7_75t_L g674 ( .A(n_20), .Y(n_674) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_21), .A2(n_74), .B(n_142), .Y(n_141) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_21), .A2(n_74), .B(n_142), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_23), .A2(n_72), .B1(n_654), .B2(n_655), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_24), .B(n_127), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_25), .A2(n_84), .B1(n_291), .B2(n_292), .Y(n_290) );
INVx2_ASAP7_75t_L g195 ( .A(n_26), .Y(n_195) );
INVx1_ASAP7_75t_L g668 ( .A(n_27), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_28), .A2(n_32), .B1(n_133), .B2(n_135), .Y(n_132) );
BUFx3_ASAP7_75t_L g108 ( .A(n_29), .Y(n_108) );
O2A1O1Ixp5_ASAP7_75t_L g189 ( .A1(n_30), .A2(n_130), .B(n_190), .C(n_192), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_31), .A2(n_67), .B1(n_155), .B2(n_191), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_33), .Y(n_232) );
AO22x1_ASAP7_75t_L g629 ( .A1(n_34), .A2(n_82), .B1(n_250), .B2(n_630), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_35), .Y(n_578) );
AND2x2_ASAP7_75t_L g592 ( .A(n_36), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_37), .B(n_250), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_38), .A2(n_85), .B1(n_210), .B2(n_213), .Y(n_209) );
INVx1_ASAP7_75t_L g547 ( .A(n_39), .Y(n_547) );
INVx1_ASAP7_75t_L g183 ( .A(n_40), .Y(n_183) );
AOI22x1_ASAP7_75t_L g701 ( .A1(n_41), .A2(n_100), .B1(n_615), .B2(n_654), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_42), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g971 ( .A(n_44), .B(n_972), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_45), .B(n_179), .Y(n_265) );
INVx2_ASAP7_75t_L g193 ( .A(n_46), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_47), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_48), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g156 ( .A(n_50), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_51), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_SL g249 ( .A(n_52), .Y(n_249) );
INVx1_ASAP7_75t_L g113 ( .A(n_53), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_54), .B(n_135), .Y(n_644) );
INVx1_ASAP7_75t_L g227 ( .A(n_55), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_56), .B(n_185), .Y(n_581) );
INVx1_ASAP7_75t_L g142 ( .A(n_57), .Y(n_142) );
AND2x4_ASAP7_75t_L g144 ( .A(n_59), .B(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g187 ( .A(n_59), .B(n_145), .Y(n_187) );
INVx1_ASAP7_75t_L g253 ( .A(n_60), .Y(n_253) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_61), .Y(n_131) );
INVx2_ASAP7_75t_L g657 ( .A(n_62), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g947 ( .A1(n_63), .A2(n_101), .B1(n_948), .B2(n_949), .Y(n_947) );
INVx1_ASAP7_75t_L g949 ( .A(n_63), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_64), .A2(n_77), .B1(n_574), .B2(n_615), .Y(n_614) );
CKINVDCx14_ASAP7_75t_R g635 ( .A(n_65), .Y(n_635) );
AND2x2_ASAP7_75t_L g599 ( .A(n_66), .B(n_250), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_68), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_69), .B(n_263), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_71), .B(n_257), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g603 ( .A(n_73), .B(n_587), .Y(n_603) );
CKINVDCx14_ASAP7_75t_R g704 ( .A(n_75), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_76), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_78), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_79), .B(n_575), .Y(n_642) );
OR2x6_ASAP7_75t_L g544 ( .A(n_80), .B(n_545), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g970 ( .A(n_80), .B(n_542), .C(n_971), .Y(n_970) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_81), .B(n_136), .Y(n_251) );
INVx1_ASAP7_75t_L g546 ( .A(n_83), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_83), .B(n_547), .Y(n_969) );
INVx1_ASAP7_75t_L g972 ( .A(n_86), .Y(n_972) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_87), .Y(n_552) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_88), .Y(n_128) );
BUFx5_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
INVx1_ASAP7_75t_L g163 ( .A(n_88), .Y(n_163) );
INVx2_ASAP7_75t_L g678 ( .A(n_89), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_90), .B(n_165), .Y(n_247) );
OAI21x1_ASAP7_75t_L g109 ( .A1(n_91), .A2(n_110), .B(n_548), .Y(n_109) );
INVx1_ASAP7_75t_L g550 ( .A(n_91), .Y(n_550) );
INVx2_ASAP7_75t_L g160 ( .A(n_92), .Y(n_160) );
INVx1_ASAP7_75t_L g170 ( .A(n_93), .Y(n_170) );
NAND2xp33_ASAP7_75t_L g595 ( .A(n_94), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g236 ( .A(n_95), .Y(n_236) );
INVx2_ASAP7_75t_SL g145 ( .A(n_96), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_97), .B(n_225), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_98), .B(n_602), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_99), .B(n_257), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g948 ( .A(n_101), .Y(n_948) );
AO32x2_ASAP7_75t_L g123 ( .A1(n_102), .A2(n_124), .A3(n_139), .B1(n_143), .B2(n_146), .Y(n_123) );
AO22x2_ASAP7_75t_L g307 ( .A1(n_102), .A2(n_124), .B1(n_308), .B2(n_310), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_103), .B(n_585), .Y(n_584) );
OA21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_109), .B(n_553), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx6p67_ASAP7_75t_R g964 ( .A(n_108), .Y(n_964) );
OR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_538), .Y(n_110) );
AOI21xp5_ASAP7_75t_SL g548 ( .A1(n_111), .A2(n_549), .B(n_551), .Y(n_548) );
XNOR2x1_ASAP7_75t_L g111 ( .A(n_112), .B(n_115), .Y(n_111) );
NOR2xp67_ASAP7_75t_L g941 ( .A(n_115), .B(n_942), .Y(n_941) );
AO22x2_ASAP7_75t_L g951 ( .A1(n_115), .A2(n_952), .B1(n_953), .B2(n_954), .Y(n_951) );
OR2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_531), .Y(n_115) );
NOR3xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_405), .C(n_463), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_117), .A2(n_533), .B(n_534), .Y(n_532) );
NAND4xp75_ASAP7_75t_L g117 ( .A(n_118), .B(n_322), .C(n_353), .D(n_386), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_297), .Y(n_118) );
AOI22xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_196), .B1(n_272), .B2(n_278), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_149), .Y(n_121) );
BUFx3_ASAP7_75t_L g336 ( .A(n_122), .Y(n_336) );
AND2x4_ASAP7_75t_L g346 ( .A(n_122), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g369 ( .A(n_122), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_SL g383 ( .A(n_122), .B(n_150), .Y(n_383) );
AND2x2_ASAP7_75t_L g452 ( .A(n_122), .B(n_424), .Y(n_452) );
AND2x2_ASAP7_75t_L g491 ( .A(n_122), .B(n_399), .Y(n_491) );
BUFx8_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g280 ( .A(n_123), .Y(n_280) );
AND2x2_ASAP7_75t_L g481 ( .A(n_123), .B(n_482), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_130), .B1(n_132), .B2(n_137), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_126), .B(n_193), .Y(n_192) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
INVx2_ASAP7_75t_L g177 ( .A(n_127), .Y(n_177) );
INVx2_ASAP7_75t_L g233 ( .A(n_127), .Y(n_233) );
INVx1_ASAP7_75t_L g596 ( .A(n_127), .Y(n_596) );
INVx1_ASAP7_75t_L g602 ( .A(n_127), .Y(n_602) );
INVx6_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g129 ( .A(n_128), .Y(n_129) );
INVx3_ASAP7_75t_L g136 ( .A(n_128), .Y(n_136) );
INVx2_ASAP7_75t_L g212 ( .A(n_128), .Y(n_212) );
INVx2_ASAP7_75t_L g185 ( .A(n_129), .Y(n_185) );
INVxp67_ASAP7_75t_SL g213 ( .A(n_129), .Y(n_213) );
INVx4_ASAP7_75t_L g230 ( .A(n_130), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_130), .A2(n_260), .B(n_262), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_130), .A2(n_574), .B1(n_576), .B2(n_579), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_130), .B(n_613), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_130), .A2(n_641), .B(n_642), .Y(n_640) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_131), .Y(n_138) );
INVx3_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
INVx4_ASAP7_75t_L g180 ( .A(n_131), .Y(n_180) );
INVx1_ASAP7_75t_L g215 ( .A(n_131), .Y(n_215) );
INVxp67_ASAP7_75t_L g597 ( .A(n_131), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_131), .B(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_131), .B(n_671), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g231 ( .A1(n_133), .A2(n_232), .B1(n_233), .B2(n_234), .Y(n_231) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g202 ( .A(n_134), .Y(n_202) );
INVx2_ASAP7_75t_L g250 ( .A(n_134), .Y(n_250) );
INVx2_ASAP7_75t_L g263 ( .A(n_134), .Y(n_263) );
INVx1_ASAP7_75t_L g267 ( .A(n_134), .Y(n_267) );
INVx2_ASAP7_75t_L g575 ( .A(n_134), .Y(n_575) );
INVx1_ASAP7_75t_L g245 ( .A(n_135), .Y(n_245) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g203 ( .A(n_136), .Y(n_203) );
INVx1_ASAP7_75t_L g261 ( .A(n_136), .Y(n_261) );
INVx2_ASAP7_75t_L g292 ( .A(n_136), .Y(n_292) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g159 ( .A1(n_138), .A2(n_160), .B(n_161), .C(n_164), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_138), .B(n_205), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_138), .A2(n_245), .B(n_246), .C(n_247), .Y(n_244) );
INVx1_ASAP7_75t_L g293 ( .A(n_138), .Y(n_293) );
INVxp67_ASAP7_75t_L g583 ( .A(n_138), .Y(n_583) );
INVx2_ASAP7_75t_SL g605 ( .A(n_138), .Y(n_605) );
INVx1_ASAP7_75t_L g646 ( .A(n_138), .Y(n_646) );
AO31x2_ASAP7_75t_L g173 ( .A1(n_139), .A2(n_174), .A3(n_188), .B(n_194), .Y(n_173) );
INVx2_ASAP7_75t_L g310 ( .A(n_139), .Y(n_310) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_140), .B(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g257 ( .A(n_140), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_140), .B(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_140), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx4_ASAP7_75t_L g243 ( .A(n_141), .Y(n_243) );
BUFx3_ASAP7_75t_L g303 ( .A(n_141), .Y(n_303) );
OAI21x1_ASAP7_75t_L g572 ( .A1(n_143), .A2(n_573), .B(n_580), .Y(n_572) );
AO31x2_ASAP7_75t_L g697 ( .A1(n_143), .A2(n_698), .A3(n_702), .B(n_703), .Y(n_697) );
AO31x2_ASAP7_75t_L g717 ( .A1(n_143), .A2(n_698), .A3(n_702), .B(n_703), .Y(n_717) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
AND2x2_ASAP7_75t_L g287 ( .A(n_144), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g308 ( .A(n_144), .B(n_309), .Y(n_308) );
INVx3_ASAP7_75t_L g608 ( .A(n_144), .Y(n_608) );
INVx1_ASAP7_75t_L g627 ( .A(n_144), .Y(n_627) );
INVxp67_ASAP7_75t_L g217 ( .A(n_146), .Y(n_217) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_147), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_148), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
NOR2xp67_ASAP7_75t_L g205 ( .A(n_148), .B(n_168), .Y(n_205) );
BUFx3_ASAP7_75t_L g207 ( .A(n_148), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_148), .B(n_168), .Y(n_271) );
INVx1_ASAP7_75t_L g309 ( .A(n_148), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_148), .B(n_168), .Y(n_613) );
INVx2_ASAP7_75t_L g652 ( .A(n_148), .Y(n_652) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g483 ( .A(n_150), .Y(n_483) );
AND2x2_ASAP7_75t_L g513 ( .A(n_150), .B(n_313), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_150), .B(n_433), .Y(n_520) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_172), .Y(n_150) );
AND2x4_ASAP7_75t_L g279 ( .A(n_151), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g305 ( .A(n_151), .B(n_173), .Y(n_305) );
INVx2_ASAP7_75t_L g317 ( .A(n_151), .Y(n_317) );
INVx1_ASAP7_75t_L g359 ( .A(n_151), .Y(n_359) );
BUFx3_ASAP7_75t_L g394 ( .A(n_151), .Y(n_394) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AO31x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_159), .A3(n_167), .B(n_169), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_156), .B(n_157), .C(n_158), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g223 ( .A(n_158), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_158), .A2(n_249), .B(n_250), .C(n_251), .Y(n_248) );
NOR2xp67_ASAP7_75t_L g220 ( .A(n_161), .B(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g291 ( .A(n_162), .Y(n_291) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g166 ( .A(n_163), .Y(n_166) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g191 ( .A(n_166), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_168), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g252 ( .A(n_171), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g621 ( .A(n_171), .Y(n_621) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_173), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g348 ( .A(n_173), .Y(n_348) );
OR2x2_ASAP7_75t_L g362 ( .A(n_173), .B(n_330), .Y(n_362) );
AND2x2_ASAP7_75t_L g424 ( .A(n_173), .B(n_317), .Y(n_424) );
AOI221x1_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_178), .B1(n_182), .B2(n_184), .C(n_186), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_181), .Y(n_178) );
AND2x2_ASAP7_75t_L g182 ( .A(n_179), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_180), .B(n_270), .Y(n_269) );
NAND3xp33_ASAP7_75t_SL g651 ( .A(n_180), .B(n_607), .C(n_652), .Y(n_651) );
NOR2xp33_ASAP7_75t_SL g673 ( .A(n_180), .B(n_674), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_180), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_185), .B(n_670), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_185), .A2(n_250), .B1(n_673), .B2(n_675), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_186), .B(n_223), .Y(n_222) );
NOR3xp33_ASAP7_75t_L g226 ( .A(n_186), .B(n_223), .C(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_186), .B(n_230), .Y(n_229) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_237), .Y(n_196) );
AND2x2_ASAP7_75t_L g446 ( .A(n_197), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g510 ( .A(n_197), .B(n_390), .Y(n_510) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_216), .Y(n_197) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_198), .Y(n_340) );
AND2x2_ASAP7_75t_L g435 ( .A(n_198), .B(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g455 ( .A(n_198), .Y(n_455) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g277 ( .A(n_199), .Y(n_277) );
AND2x2_ASAP7_75t_L g299 ( .A(n_199), .B(n_255), .Y(n_299) );
INVx1_ASAP7_75t_L g366 ( .A(n_199), .Y(n_366) );
AND2x2_ASAP7_75t_L g373 ( .A(n_199), .B(n_343), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g199 ( .A(n_200), .B(n_208), .Y(n_199) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_200), .B(n_208), .Y(n_420) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_204), .B(n_206), .Y(n_200) );
INVx2_ASAP7_75t_L g654 ( .A(n_202), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_205), .B(n_215), .Y(n_214) );
OR2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_214), .Y(n_208) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g225 ( .A(n_212), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_215), .B(n_613), .Y(n_617) );
INVx1_ASAP7_75t_L g700 ( .A(n_215), .Y(n_700) );
AND2x2_ASAP7_75t_L g320 ( .A(n_216), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g342 ( .A(n_216), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g367 ( .A(n_216), .B(n_240), .Y(n_367) );
AND2x2_ASAP7_75t_L g512 ( .A(n_216), .B(n_419), .Y(n_512) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_235), .Y(n_216) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_218), .A2(n_235), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_228), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_222), .B1(n_224), .B2(n_226), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_223), .A2(n_290), .B1(n_293), .B2(n_294), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g659 ( .A(n_223), .B(n_607), .C(n_652), .Y(n_659) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_230), .B(n_577), .Y(n_576) );
OAI22x1_ASAP7_75t_L g698 ( .A1(n_230), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_233), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g593 ( .A(n_233), .Y(n_593) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_254), .Y(n_237) );
AND2x2_ASAP7_75t_L g319 ( .A(n_238), .B(n_277), .Y(n_319) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_238), .Y(n_325) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g283 ( .A(n_240), .Y(n_283) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_240), .Y(n_345) );
OR2x2_ASAP7_75t_L g379 ( .A(n_240), .B(n_301), .Y(n_379) );
INVx2_ASAP7_75t_L g391 ( .A(n_240), .Y(n_391) );
INVx1_ASAP7_75t_L g448 ( .A(n_240), .Y(n_448) );
AO31x2_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_244), .A3(n_248), .B(n_252), .Y(n_240) );
INVx2_ASAP7_75t_L g288 ( .A(n_242), .Y(n_288) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx3_ASAP7_75t_L g587 ( .A(n_243), .Y(n_587) );
INVx1_ASAP7_75t_L g461 ( .A(n_254), .Y(n_461) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g275 ( .A(n_255), .Y(n_275) );
INVx1_ASAP7_75t_L g321 ( .A(n_255), .Y(n_321) );
INVx2_ASAP7_75t_L g343 ( .A(n_255), .Y(n_343) );
AND2x2_ASAP7_75t_L g390 ( .A(n_255), .B(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
NOR2x1_ASAP7_75t_L g647 ( .A(n_257), .B(n_608), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_264), .B(n_271), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_266), .B(n_268), .Y(n_264) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVxp67_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx2_ASAP7_75t_L g326 ( .A(n_274), .Y(n_326) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g495 ( .A(n_275), .B(n_420), .Y(n_495) );
INVx1_ASAP7_75t_L g505 ( .A(n_276), .Y(n_505) );
BUFx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_279), .B(n_314), .Y(n_472) );
INVx2_ASAP7_75t_L g488 ( .A(n_279), .Y(n_488) );
AND2x2_ASAP7_75t_L g508 ( .A(n_279), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g398 ( .A(n_280), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_280), .B(n_348), .Y(n_459) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
AND2x2_ASAP7_75t_L g334 ( .A(n_283), .B(n_301), .Y(n_334) );
INVxp67_ASAP7_75t_SL g475 ( .A(n_283), .Y(n_475) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_283), .Y(n_523) );
AND2x2_ASAP7_75t_L g371 ( .A(n_284), .B(n_358), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_284), .B(n_399), .Y(n_427) );
BUFx3_ASAP7_75t_L g444 ( .A(n_284), .Y(n_444) );
AND2x2_ASAP7_75t_L g462 ( .A(n_284), .B(n_424), .Y(n_462) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_285), .Y(n_333) );
AND2x2_ASAP7_75t_L g347 ( .A(n_285), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g490 ( .A(n_285), .B(n_317), .Y(n_490) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g315 ( .A(n_286), .Y(n_315) );
INVx1_ASAP7_75t_L g330 ( .A(n_286), .Y(n_330) );
AOI21x1_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_289), .B(n_295), .Y(n_286) );
AOI21xp33_ASAP7_75t_SL g606 ( .A1(n_288), .A2(n_607), .B(n_609), .Y(n_606) );
INVx2_ASAP7_75t_L g630 ( .A(n_291), .Y(n_630) );
INVx1_ASAP7_75t_L g619 ( .A(n_292), .Y(n_619) );
INVx1_ASAP7_75t_L g655 ( .A(n_292), .Y(n_655) );
AOI21x1_ASAP7_75t_L g628 ( .A1(n_293), .A2(n_629), .B(n_631), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_304), .B1(n_311), .B2(n_318), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g350 ( .A(n_298), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g337 ( .A(n_299), .Y(n_337) );
AND2x2_ASAP7_75t_L g344 ( .A(n_299), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g425 ( .A(n_299), .B(n_367), .Y(n_425) );
AND2x2_ASAP7_75t_L g516 ( .A(n_299), .B(n_334), .Y(n_516) );
INVx2_ASAP7_75t_L g415 ( .A(n_300), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_300), .B(n_373), .Y(n_467) );
BUFx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g436 ( .A(n_301), .Y(n_436) );
OR2x2_ASAP7_75t_L g634 ( .A(n_302), .B(n_635), .Y(n_634) );
NOR2xp67_ASAP7_75t_SL g703 ( .A(n_302), .B(n_704), .Y(n_703) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OA21x2_ASAP7_75t_L g571 ( .A1(n_303), .A2(n_572), .B(n_584), .Y(n_571) );
OA21x2_ASAP7_75t_L g687 ( .A1(n_303), .A2(n_572), .B(n_584), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_304), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_305), .B(n_313), .Y(n_352) );
INVx2_ASAP7_75t_L g401 ( .A(n_305), .Y(n_401) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g316 ( .A(n_307), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g360 ( .A(n_307), .Y(n_360) );
AND2x4_ASAP7_75t_L g393 ( .A(n_307), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g433 ( .A(n_307), .B(n_330), .Y(n_433) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .Y(n_312) );
AND2x4_ASAP7_75t_L g397 ( .A(n_313), .B(n_398), .Y(n_397) );
INVx4_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g423 ( .A(n_314), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g509 ( .A(n_314), .Y(n_509) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g482 ( .A(n_315), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_316), .B(n_328), .Y(n_327) );
INVx4_ASAP7_75t_L g421 ( .A(n_316), .Y(n_421) );
AND2x4_ASAP7_75t_L g469 ( .A(n_316), .B(n_470), .Y(n_469) );
AND2x4_ASAP7_75t_L g501 ( .A(n_316), .B(n_361), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_318), .A2(n_423), .B1(n_425), .B2(n_426), .Y(n_422) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g411 ( .A(n_319), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g447 ( .A(n_321), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g504 ( .A(n_321), .Y(n_504) );
NOR3x1_ASAP7_75t_L g322 ( .A(n_323), .B(n_338), .C(n_349), .Y(n_322) );
OAI21xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .B(n_331), .Y(n_323) );
NOR3xp33_ASAP7_75t_L g413 ( .A(n_324), .B(n_414), .C(n_418), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g438 ( .A(n_328), .B(n_421), .Y(n_438) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g370 ( .A(n_329), .Y(n_370) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_330), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_335), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g440 ( .A(n_334), .B(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_337), .B(n_522), .Y(n_521) );
OA21x2_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_344), .B(n_346), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVxp67_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g412 ( .A(n_342), .Y(n_412) );
OR2x6_ASAP7_75t_L g474 ( .A(n_342), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g451 ( .A(n_347), .B(n_358), .Y(n_451) );
INVx2_ASAP7_75t_SL g399 ( .A(n_348), .Y(n_399) );
INVx1_ASAP7_75t_L g417 ( .A(n_348), .Y(n_417) );
BUFx3_ASAP7_75t_L g470 ( .A(n_348), .Y(n_470) );
INVxp67_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_351), .A2(n_503), .B1(n_526), .B2(n_528), .Y(n_525) );
INVx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NOR2x1_ASAP7_75t_L g353 ( .A(n_354), .B(n_374), .Y(n_353) );
OAI21xp5_ASAP7_75t_SL g354 ( .A1(n_355), .A2(n_363), .B(n_368), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_361), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_358), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g445 ( .A(n_358), .Y(n_445) );
AND2x4_ASAP7_75t_SL g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_362), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_471) );
OAI21xp5_ASAP7_75t_SL g487 ( .A1(n_362), .A2(n_488), .B(n_489), .Y(n_487) );
INVx2_ASAP7_75t_L g530 ( .A(n_362), .Y(n_530) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
OR2x2_ASAP7_75t_L g385 ( .A(n_365), .B(n_379), .Y(n_385) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g389 ( .A(n_366), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g372 ( .A(n_367), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g454 ( .A(n_367), .B(n_455), .Y(n_454) );
OAI21xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B(n_372), .Y(n_368) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_371), .Y(n_375) );
BUFx3_ASAP7_75t_L g381 ( .A(n_373), .Y(n_381) );
NAND2xp67_ASAP7_75t_L g403 ( .A(n_373), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_373), .B(n_415), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B(n_382), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_380), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g404 ( .A(n_379), .Y(n_404) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OA21x2_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_392), .B(n_396), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_388), .A2(n_457), .B1(n_460), .B2(n_462), .Y(n_456) );
BUFx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g468 ( .A(n_389), .Y(n_468) );
AND2x2_ASAP7_75t_L g434 ( .A(n_390), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g494 ( .A(n_391), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx2_ASAP7_75t_L g431 ( .A(n_393), .Y(n_431) );
OAI21xp33_ASAP7_75t_L g443 ( .A1(n_393), .A2(n_444), .B(n_445), .Y(n_443) );
NAND3xp33_ASAP7_75t_L g502 ( .A(n_393), .B(n_503), .C(n_505), .Y(n_502) );
AND2x2_ASAP7_75t_L g524 ( .A(n_393), .B(n_509), .Y(n_524) );
INVx2_ASAP7_75t_SL g529 ( .A(n_394), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_395), .B(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g458 ( .A(n_395), .B(n_459), .Y(n_458) );
OAI21xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .B(n_402), .Y(n_396) );
INVx1_ASAP7_75t_L g410 ( .A(n_399), .Y(n_410) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g536 ( .A(n_406), .Y(n_536) );
NOR3x1_ASAP7_75t_L g406 ( .A(n_407), .B(n_428), .C(n_449), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_422), .Y(n_407) );
A2O1A1Ixp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B(n_413), .C(n_421), .Y(n_408) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g527 ( .A(n_412), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g441 ( .A(n_420), .Y(n_441) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_426), .A2(n_515), .B(n_516), .Y(n_514) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_437), .C(n_442), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_434), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
AND2x4_ASAP7_75t_L g460 ( .A(n_435), .B(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g493 ( .A(n_436), .B(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_441), .B(n_493), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_446), .Y(n_442) );
INVx1_ASAP7_75t_L g478 ( .A(n_444), .Y(n_478) );
INVx1_ASAP7_75t_L g484 ( .A(n_447), .Y(n_484) );
AND2x4_ASAP7_75t_L g511 ( .A(n_447), .B(n_512), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_453), .B(n_456), .Y(n_449) );
NOR2x1_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_452), .A2(n_460), .B1(n_499), .B2(n_501), .Y(n_498) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_454), .A2(n_519), .B1(n_521), .B2(n_524), .Y(n_518) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_496), .Y(n_463) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_476), .C(n_485), .Y(n_464) );
OR3x1_ASAP7_75t_L g533 ( .A(n_465), .B(n_476), .C(n_485), .Y(n_533) );
AO21x1_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_469), .B(n_471), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_470), .B(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g515 ( .A(n_470), .B(n_490), .Y(n_515) );
AOI21xp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_479), .B(n_484), .Y(n_476) );
OR2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_483), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI21xp33_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_491), .B(n_492), .Y(n_486) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
AND2x4_ASAP7_75t_L g503 ( .A(n_493), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g537 ( .A(n_496), .Y(n_537) );
NOR3xp33_ASAP7_75t_SL g496 ( .A(n_497), .B(n_506), .C(n_517), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_498), .B(n_502), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_507), .B(n_514), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_510), .B1(n_511), .B2(n_513), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_525), .Y(n_517) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_535), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g535 ( .A1(n_534), .A2(n_536), .B(n_537), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_538), .B(n_550), .Y(n_549) );
INVx5_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_540), .B(n_552), .Y(n_551) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
OR2x6_ASAP7_75t_L g560 ( .A(n_543), .B(n_561), .Y(n_560) );
INVx8_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g943 ( .A(n_544), .B(n_944), .Y(n_943) );
OR2x6_ASAP7_75t_L g962 ( .A(n_544), .B(n_944), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g956 ( .A(n_551), .Y(n_956) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_554), .B(n_950), .Y(n_553) );
NAND2xp33_ASAP7_75t_SL g554 ( .A(n_555), .B(n_945), .Y(n_554) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_562), .B(n_941), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g952 ( .A(n_557), .Y(n_952) );
BUFx12f_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
CKINVDCx11_ASAP7_75t_R g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g953 ( .A(n_562), .Y(n_953) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND3x1_ASAP7_75t_L g563 ( .A(n_564), .B(n_804), .C(n_880), .Y(n_563) );
NOR2x1_ASAP7_75t_L g564 ( .A(n_565), .B(n_733), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_688), .C(n_713), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_622), .B1(n_679), .B2(n_683), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_588), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_569), .B(n_752), .Y(n_902) );
AND3x2_ASAP7_75t_L g908 ( .A(n_569), .B(n_685), .C(n_788), .Y(n_908) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g741 ( .A(n_570), .B(n_697), .Y(n_741) );
AND2x2_ASAP7_75t_L g778 ( .A(n_570), .B(n_610), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_570), .B(n_821), .Y(n_856) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g728 ( .A(n_571), .Y(n_728) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B(n_583), .Y(n_580) );
OR2x2_ASAP7_75t_L g626 ( .A(n_585), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g656 ( .A(n_586), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_610), .Y(n_588) );
INVx1_ASAP7_75t_L g939 ( .A(n_589), .Y(n_939) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVxp67_ASAP7_75t_L g685 ( .A(n_590), .Y(n_685) );
AND2x2_ASAP7_75t_L g695 ( .A(n_590), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g740 ( .A(n_590), .Y(n_740) );
AO21x2_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_598), .B(n_606), .Y(n_590) );
AO21x2_ASAP7_75t_L g720 ( .A1(n_591), .A2(n_598), .B(n_606), .Y(n_720) );
OAI21x1_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_594), .B(n_597), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_593), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g615 ( .A(n_596), .Y(n_615) );
OAI21x1_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_600), .B(n_604), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_603), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g609 ( .A(n_603), .Y(n_609) );
AOI21x1_ASAP7_75t_L g631 ( .A1(n_605), .A2(n_632), .B(n_633), .Y(n_631) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g686 ( .A(n_610), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g725 ( .A(n_610), .Y(n_725) );
INVx1_ASAP7_75t_L g765 ( .A(n_610), .Y(n_765) );
INVx2_ASAP7_75t_L g821 ( .A(n_610), .Y(n_821) );
NAND2x1p5_ASAP7_75t_L g610 ( .A(n_611), .B(n_616), .Y(n_610) );
AND2x2_ASAP7_75t_L g693 ( .A(n_611), .B(n_616), .Y(n_693) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
OA21x2_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B(n_620), .Y(n_616) );
INVx1_ASAP7_75t_L g702 ( .A(n_621), .Y(n_702) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_648), .Y(n_623) );
INVx2_ASAP7_75t_L g748 ( .A(n_624), .Y(n_748) );
AND2x4_ASAP7_75t_L g784 ( .A(n_624), .B(n_785), .Y(n_784) );
AND2x2_ASAP7_75t_L g870 ( .A(n_624), .B(n_769), .Y(n_870) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_636), .Y(n_624) );
AND2x2_ASAP7_75t_L g681 ( .A(n_625), .B(n_637), .Y(n_681) );
INVx2_ASAP7_75t_SL g712 ( .A(n_625), .Y(n_712) );
OAI21x1_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_628), .B(n_634), .Y(n_625) );
OAI21xp5_ASAP7_75t_L g827 ( .A1(n_626), .A2(n_628), .B(n_634), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_627), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g757 ( .A(n_636), .Y(n_757) );
AND2x2_ASAP7_75t_L g879 ( .A(n_636), .B(n_649), .Y(n_879) );
INVx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g708 ( .A(n_637), .Y(n_708) );
AND2x2_ASAP7_75t_L g800 ( .A(n_637), .B(n_712), .Y(n_800) );
AND2x4_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
OAI21x1_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_643), .B(n_647), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B(n_646), .Y(n_643) );
INVx2_ASAP7_75t_L g682 ( .A(n_648), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_648), .B(n_791), .Y(n_790) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_648), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_648), .B(n_934), .Y(n_933) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_661), .Y(n_648) );
INVx1_ASAP7_75t_L g709 ( .A(n_649), .Y(n_709) );
INVx1_ASAP7_75t_L g747 ( .A(n_649), .Y(n_747) );
INVx1_ASAP7_75t_L g755 ( .A(n_649), .Y(n_755) );
INVx2_ASAP7_75t_L g770 ( .A(n_649), .Y(n_770) );
NOR2x1_ASAP7_75t_L g785 ( .A(n_649), .B(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_L g796 ( .A(n_649), .B(n_662), .Y(n_796) );
OR2x6_ASAP7_75t_L g649 ( .A(n_650), .B(n_658), .Y(n_649) );
OAI21x1_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_653), .B(n_656), .Y(n_650) );
INVx1_ASAP7_75t_L g664 ( .A(n_652), .Y(n_664) );
NOR2xp67_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
AND2x2_ASAP7_75t_L g769 ( .A(n_661), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g711 ( .A(n_662), .B(n_712), .Y(n_711) );
INVxp67_ASAP7_75t_L g732 ( .A(n_662), .Y(n_732) );
INVx1_ASAP7_75t_L g781 ( .A(n_662), .Y(n_781) );
INVx1_ASAP7_75t_L g786 ( .A(n_662), .Y(n_786) );
OR2x2_ASAP7_75t_L g826 ( .A(n_662), .B(n_827), .Y(n_826) );
AO21x2_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_665), .B(n_677), .Y(n_662) );
NAND3xp33_ASAP7_75t_SL g665 ( .A(n_666), .B(n_669), .C(n_672), .Y(n_665) );
NAND2xp33_ASAP7_75t_SL g851 ( .A(n_679), .B(n_852), .Y(n_851) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g803 ( .A(n_681), .B(n_796), .Y(n_803) );
AND2x2_ASAP7_75t_L g818 ( .A(n_681), .B(n_746), .Y(n_818) );
AND2x2_ASAP7_75t_L g831 ( .A(n_681), .B(n_832), .Y(n_831) );
HB1xp67_ASAP7_75t_L g926 ( .A(n_682), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_683), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_686), .B(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_686), .B(n_876), .Y(n_875) );
AND2x2_ASAP7_75t_L g935 ( .A(n_686), .B(n_936), .Y(n_935) );
AND2x2_ASAP7_75t_L g692 ( .A(n_687), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g719 ( .A(n_687), .B(n_720), .Y(n_719) );
NAND2x1_ASAP7_75t_L g762 ( .A(n_687), .B(n_696), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_689), .B(n_705), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_694), .Y(n_690) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x4_ASAP7_75t_L g751 ( .A(n_692), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g844 ( .A(n_692), .Y(n_844) );
AND2x2_ASAP7_75t_L g864 ( .A(n_692), .B(n_743), .Y(n_864) );
INVx2_ASAP7_75t_SL g722 ( .A(n_693), .Y(n_722) );
BUFx3_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_695), .B(n_838), .Y(n_837) );
AND2x2_ASAP7_75t_L g894 ( .A(n_695), .B(n_788), .Y(n_894) );
AOI32xp33_ASAP7_75t_L g904 ( .A1(n_695), .A2(n_825), .A3(n_905), .B1(n_906), .B2(n_908), .Y(n_904) );
INVx2_ASAP7_75t_L g730 ( .A(n_696), .Y(n_730) );
INVx1_ASAP7_75t_L g936 ( .A(n_696), .Y(n_936) );
INVx3_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OAI321xp33_ASAP7_75t_L g923 ( .A1(n_706), .A2(n_924), .A3(n_926), .B1(n_927), .B2(n_929), .C(n_930), .Y(n_923) );
NAND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_710), .Y(n_706) );
AND2x2_ASAP7_75t_L g887 ( .A(n_707), .B(n_825), .Y(n_887) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_708), .B(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g768 ( .A(n_708), .Y(n_768) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_708), .Y(n_824) );
OR2x2_ASAP7_75t_L g843 ( .A(n_708), .B(n_826), .Y(n_843) );
OR2x2_ASAP7_75t_L g866 ( .A(n_709), .B(n_748), .Y(n_866) );
AND2x2_ASAP7_75t_L g914 ( .A(n_709), .B(n_800), .Y(n_914) );
BUFx3_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_711), .B(n_755), .Y(n_774) );
AND2x4_ASAP7_75t_L g878 ( .A(n_711), .B(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g758 ( .A(n_712), .Y(n_758) );
INVx1_ASAP7_75t_L g791 ( .A(n_712), .Y(n_791) );
OAI21xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_723), .B(n_731), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_716), .B(n_728), .Y(n_859) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g744 ( .A(n_717), .B(n_720), .Y(n_744) );
AND2x4_ASAP7_75t_L g752 ( .A(n_717), .B(n_740), .Y(n_752) );
AND2x2_ASAP7_75t_L g766 ( .A(n_717), .B(n_720), .Y(n_766) );
INVx2_ASAP7_75t_L g801 ( .A(n_718), .Y(n_801) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_721), .Y(n_718) );
INVx2_ASAP7_75t_L g849 ( .A(n_719), .Y(n_849) );
AND2x2_ASAP7_75t_L g867 ( .A(n_719), .B(n_729), .Y(n_867) );
AND2x4_ASAP7_75t_L g727 ( .A(n_720), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g761 ( .A(n_722), .B(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g788 ( .A(n_722), .Y(n_788) );
AND2x2_ASAP7_75t_L g850 ( .A(n_722), .B(n_730), .Y(n_850) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
AND2x2_ASAP7_75t_L g905 ( .A(n_724), .B(n_779), .Y(n_905) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g783 ( .A1(n_726), .A2(n_784), .B1(n_787), .B2(n_789), .C(n_792), .Y(n_783) );
AND2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
AND2x2_ASAP7_75t_L g820 ( .A(n_727), .B(n_821), .Y(n_820) );
BUFx3_ASAP7_75t_L g861 ( .A(n_727), .Y(n_861) );
INVxp67_ASAP7_75t_SL g884 ( .A(n_728), .Y(n_884) );
INVx1_ASAP7_75t_L g916 ( .A(n_729), .Y(n_916) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g809 ( .A(n_730), .Y(n_809) );
AND2x2_ASAP7_75t_L g912 ( .A(n_731), .B(n_891), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_783), .Y(n_733) );
NOR3xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_749), .C(n_771), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_745), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_742), .Y(n_736) );
OAI21xp33_ASAP7_75t_L g771 ( .A1(n_737), .A2(n_772), .B(n_775), .Y(n_771) );
NAND2x1p5_ASAP7_75t_L g737 ( .A(n_738), .B(n_741), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g929 ( .A(n_741), .Y(n_929) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g794 ( .A(n_744), .Y(n_794) );
INVx1_ASAP7_75t_L g846 ( .A(n_745), .Y(n_846) );
OR2x2_ASAP7_75t_SL g745 ( .A(n_746), .B(n_748), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_L g931 ( .A(n_747), .B(n_922), .Y(n_931) );
OR2x2_ASAP7_75t_L g812 ( .A(n_748), .B(n_813), .Y(n_812) );
OAI21xp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_753), .B(n_759), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
BUFx3_ASAP7_75t_L g782 ( .A(n_752), .Y(n_782) );
AND2x2_ASAP7_75t_L g787 ( .A(n_752), .B(n_788), .Y(n_787) );
NOR2xp67_ASAP7_75t_L g816 ( .A(n_752), .B(n_777), .Y(n_816) );
INVx3_ASAP7_75t_L g876 ( .A(n_752), .Y(n_876) );
OR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g891 ( .A(n_755), .B(n_892), .Y(n_891) );
OR2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g779 ( .A(n_757), .Y(n_779) );
INVxp67_ASAP7_75t_SL g841 ( .A(n_758), .Y(n_841) );
OAI21xp33_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_763), .B(n_767), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g832 ( .A(n_765), .Y(n_832) );
INVx1_ASAP7_75t_L g910 ( .A(n_765), .Y(n_910) );
NOR3xp33_ASAP7_75t_L g872 ( .A(n_766), .B(n_794), .C(n_850), .Y(n_872) );
INVx2_ASAP7_75t_L g911 ( .A(n_766), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g913 ( .A1(n_766), .A2(n_914), .B1(n_915), .B2(n_918), .Y(n_913) );
AND2x2_ASAP7_75t_L g928 ( .A(n_766), .B(n_788), .Y(n_928) );
INVx2_ASAP7_75t_L g897 ( .A(n_767), .Y(n_897) );
AND2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
AND2x2_ASAP7_75t_L g890 ( .A(n_768), .B(n_781), .Y(n_890) );
INVx1_ASAP7_75t_L g934 ( .A(n_768), .Y(n_934) );
AND2x2_ASAP7_75t_L g874 ( .A(n_769), .B(n_800), .Y(n_874) );
INVx1_ASAP7_75t_L g907 ( .A(n_769), .Y(n_907) );
OAI21xp33_ASAP7_75t_L g937 ( .A1(n_772), .A2(n_938), .B(n_940), .Y(n_937) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NAND4xp25_ASAP7_75t_L g775 ( .A(n_776), .B(n_779), .C(n_780), .D(n_782), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g810 ( .A(n_778), .Y(n_810) );
INVx1_ASAP7_75t_L g925 ( .A(n_779), .Y(n_925) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g852 ( .A(n_784), .Y(n_852) );
NAND2x1_ASAP7_75t_L g793 ( .A(n_788), .B(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_789), .B(n_820), .Y(n_940) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OAI32xp33_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_795), .A3(n_797), .B1(n_801), .B2(n_802), .Y(n_792) );
INVx1_ASAP7_75t_L g806 ( .A(n_793), .Y(n_806) );
A2O1A1Ixp33_ASAP7_75t_L g909 ( .A1(n_794), .A2(n_910), .B(n_911), .C(n_912), .Y(n_909) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g813 ( .A(n_796), .Y(n_813) );
AND2x2_ASAP7_75t_L g840 ( .A(n_796), .B(n_841), .Y(n_840) );
NAND2x1_ASAP7_75t_SL g862 ( .A(n_796), .B(n_800), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_796), .B(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AND4x1_ASAP7_75t_L g804 ( .A(n_805), .B(n_828), .C(n_845), .D(n_863), .Y(n_804) );
O2A1O1Ixp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_807), .B(n_811), .C(n_814), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
NAND2xp5_ASAP7_75t_SL g830 ( .A(n_809), .B(n_831), .Y(n_830) );
INVx2_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_817), .B1(n_819), .B2(n_822), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g838 ( .A(n_821), .Y(n_838) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g922 ( .A(n_826), .Y(n_922) );
BUFx2_ASAP7_75t_L g892 ( .A(n_827), .Y(n_892) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_833), .B(n_836), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
OR2x2_ASAP7_75t_L g858 ( .A(n_832), .B(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
OAI22xp5_ASAP7_75t_SL g836 ( .A1(n_837), .A2(n_839), .B1(n_842), .B2(n_844), .Y(n_836) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
AOI221xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_847), .B1(n_851), .B2(n_853), .C(n_857), .Y(n_845) );
AND2x4_ASAP7_75t_L g847 ( .A(n_848), .B(n_850), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g917 ( .A(n_849), .Y(n_917) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
OR2x2_ASAP7_75t_L g938 ( .A(n_856), .B(n_939), .Y(n_938) );
AOI21xp33_ASAP7_75t_SL g857 ( .A1(n_858), .A2(n_860), .B(n_862), .Y(n_857) );
INVx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
AOI221xp5_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_865), .B1(n_867), .B2(n_868), .C(n_871), .Y(n_863) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
OAI22xp33_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_873), .B1(n_875), .B2(n_877), .Y(n_871) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g885 ( .A(n_876), .Y(n_885) );
INVx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx2_ASAP7_75t_L g920 ( .A(n_879), .Y(n_920) );
NOR4xp25_ASAP7_75t_L g880 ( .A(n_881), .B(n_903), .C(n_923), .D(n_937), .Y(n_880) );
OAI322xp33_ASAP7_75t_L g881 ( .A1(n_882), .A2(n_885), .A3(n_886), .B1(n_888), .B2(n_893), .C1(n_895), .C2(n_901), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
INVx1_ASAP7_75t_L g900 ( .A(n_892), .Y(n_900) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
INVxp67_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
HB1xp67_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
NAND3xp33_ASAP7_75t_SL g903 ( .A(n_904), .B(n_909), .C(n_913), .Y(n_903) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
AND2x2_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .Y(n_915) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
OR2x2_ASAP7_75t_L g919 ( .A(n_920), .B(n_921), .Y(n_919) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
OAI21xp5_ASAP7_75t_L g930 ( .A1(n_931), .A2(n_932), .B(n_935), .Y(n_930) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_SL g942 ( .A(n_943), .Y(n_942) );
HB1xp67_ASAP7_75t_L g954 ( .A(n_943), .Y(n_954) );
INVxp67_ASAP7_75t_R g945 ( .A(n_946), .Y(n_945) );
AOI21xp33_ASAP7_75t_SL g950 ( .A1(n_946), .A2(n_951), .B(n_955), .Y(n_950) );
NAND3xp33_ASAP7_75t_L g955 ( .A(n_956), .B(n_957), .C(n_963), .Y(n_955) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_959), .B(n_960), .Y(n_958) );
BUFx3_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
HB1xp67_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVx1_ASAP7_75t_SL g963 ( .A(n_964), .Y(n_963) );
BUFx4_ASAP7_75t_SL g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
BUFx3_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
OR2x6_ASAP7_75t_SL g968 ( .A(n_969), .B(n_970), .Y(n_968) );
endmodule