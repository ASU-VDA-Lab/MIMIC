module fake_jpeg_30041_n_212 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_212);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_49),
.Y(n_58)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_22),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_65),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_17),
.B1(n_25),
.B2(n_19),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_79),
.B1(n_52),
.B2(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_31),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_34),
.CON(n_67),
.SN(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_72),
.B(n_80),
.C(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_41),
.B(n_31),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_30),
.B(n_29),
.C(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_3),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_32),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_81),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_36),
.A2(n_25),
.B1(n_23),
.B2(n_19),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_50),
.B(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_22),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_38),
.C(n_45),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_96),
.C(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_98),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_42),
.B1(n_37),
.B2(n_38),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_108),
.B1(n_57),
.B2(n_76),
.Y(n_123)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_67),
.A2(n_39),
.B1(n_23),
.B2(n_46),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_83),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_99),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_49),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_110),
.B1(n_60),
.B2(n_8),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_14),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_14),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_101),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_105),
.B(n_111),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_4),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_6),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_11),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_109),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_60),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_12),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_54),
.B1(n_69),
.B2(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_116),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_77),
.B1(n_57),
.B2(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_121),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_94),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_72),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_132),
.C(n_98),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_85),
.B(n_12),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_15),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_105),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_83),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_134),
.A2(n_92),
.B1(n_101),
.B2(n_86),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_95),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_139),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_113),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_143),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_147),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_103),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_148),
.A2(n_120),
.B1(n_92),
.B2(n_127),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_151),
.B(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_120),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_122),
.B1(n_116),
.B2(n_118),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_157),
.B1(n_160),
.B2(n_7),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_122),
.B1(n_149),
.B2(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_122),
.B(n_121),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_154),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_114),
.B(n_117),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_167),
.B(n_146),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_109),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_102),
.B(n_89),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_166),
.B(n_152),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_182),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_149),
.B1(n_144),
.B2(n_136),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_173),
.A2(n_164),
.B1(n_170),
.B2(n_156),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_137),
.B(n_141),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_174),
.A2(n_161),
.B(n_167),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_179),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_110),
.C(n_104),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_104),
.C(n_7),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_180),
.Y(n_186)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_181),
.Y(n_188)
);

XOR2x2_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_163),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_165),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_173),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_194),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_185),
.A2(n_186),
.B1(n_174),
.B2(n_189),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_193),
.A2(n_196),
.B1(n_189),
.B2(n_181),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_177),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_197),
.C(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_200),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_170),
.C(n_176),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_202),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_195),
.A2(n_176),
.B1(n_162),
.B2(n_160),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_198),
.B(n_168),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_180),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_201),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_204),
.C(n_205),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_208),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_8),
.B1(n_188),
.B2(n_210),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_8),
.Y(n_212)
);


endmodule