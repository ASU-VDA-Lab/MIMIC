module fake_ariane_2634_n_2271 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_34, n_404, n_172, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_636, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_630, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_641, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_2271);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_630;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_641;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2271;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_2248;
wire n_813;
wire n_1985;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_1107;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2233;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_2185;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_1139;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_2220;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_1029;
wire n_1247;
wire n_760;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2168;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_2059;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_2075;
wire n_1726;
wire n_1945;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_1783;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_876;
wire n_791;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_1757;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_2158;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_683;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_1739;
wire n_1814;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_2097;
wire n_1982;
wire n_662;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_462),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_188),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_562),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_452),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_201),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_603),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_627),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_380),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_208),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_166),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_87),
.Y(n_667)
);

CKINVDCx16_ASAP7_75t_R g668 ( 
.A(n_303),
.Y(n_668)
);

BUFx2_ASAP7_75t_SL g669 ( 
.A(n_595),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_655),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_597),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_626),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_539),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_610),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_625),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_53),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_227),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_37),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_266),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_237),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_465),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_148),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_556),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_619),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_492),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_135),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_153),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_107),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_528),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_50),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_618),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_378),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_608),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_604),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_445),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_501),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_384),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_602),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_314),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_116),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_52),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_196),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_496),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_87),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_383),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_198),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_223),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_137),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_535),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_645),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_311),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_596),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_158),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_514),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_472),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_534),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_580),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_469),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_327),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_191),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_50),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_238),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_568),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_549),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_409),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_577),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_498),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_241),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_632),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_102),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_213),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_162),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_616),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_278),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_279),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_302),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_431),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_224),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_599),
.Y(n_739)
);

BUFx5_ASAP7_75t_L g740 ( 
.A(n_620),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_605),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_335),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_600),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_27),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_601),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_436),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_398),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_624),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_594),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_614),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_270),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_628),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_127),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_19),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_68),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_441),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_306),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_67),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_83),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_370),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_641),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_656),
.Y(n_762)
);

BUFx10_ASAP7_75t_L g763 ( 
.A(n_142),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_629),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_612),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_215),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_613),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_88),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_527),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_132),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_622),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_543),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_76),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_161),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_640),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_68),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_606),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_264),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_591),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_448),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_74),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_154),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_165),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_576),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_163),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_95),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_337),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_78),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_459),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_582),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_647),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_37),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_405),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_185),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_529),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_328),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_544),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_607),
.Y(n_798)
);

CKINVDCx16_ASAP7_75t_R g799 ( 
.A(n_490),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_371),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_524),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_344),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_623),
.Y(n_803)
);

BUFx5_ASAP7_75t_L g804 ( 
.A(n_362),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_611),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_617),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_481),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_621),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_587),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_521),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_363),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_598),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_247),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_345),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_593),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_419),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_274),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_28),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_140),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_40),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_374),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_609),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_273),
.Y(n_823)
);

BUFx10_ASAP7_75t_L g824 ( 
.A(n_643),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_133),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_457),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_19),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_287),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_454),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_433),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_104),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_615),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_55),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_688),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_700),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_704),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_754),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_759),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_721),
.Y(n_839)
);

CKINVDCx16_ASAP7_75t_R g840 ( 
.A(n_668),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_768),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_781),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_788),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_820),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_690),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_657),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_827),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_678),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_721),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_721),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_772),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_823),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_718),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_789),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_821),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_763),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_786),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_763),
.Y(n_858)
);

INVxp33_ASAP7_75t_SL g859 ( 
.A(n_667),
.Y(n_859)
);

INVxp67_ASAP7_75t_SL g860 ( 
.A(n_673),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_824),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_666),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_677),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_824),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_658),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_676),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_660),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_675),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_680),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_705),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_681),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_683),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_674),
.Y(n_873)
);

CKINVDCx16_ASAP7_75t_R g874 ( 
.A(n_799),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_701),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_687),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_689),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_693),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_695),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_730),
.Y(n_880)
);

CKINVDCx14_ASAP7_75t_R g881 ( 
.A(n_715),
.Y(n_881)
);

INVxp67_ASAP7_75t_SL g882 ( 
.A(n_753),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_739),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_809),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_697),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_708),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_714),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_748),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_716),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_816),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_719),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_806),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_722),
.Y(n_893)
);

CKINVDCx16_ASAP7_75t_R g894 ( 
.A(n_774),
.Y(n_894)
);

CKINVDCx16_ASAP7_75t_R g895 ( 
.A(n_779),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_723),
.Y(n_896)
);

INVxp67_ASAP7_75t_SL g897 ( 
.A(n_703),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_725),
.Y(n_898)
);

INVx1_ASAP7_75t_SL g899 ( 
.A(n_831),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_744),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_732),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_733),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_787),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_795),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_830),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_736),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_755),
.Y(n_907)
);

BUFx2_ASAP7_75t_SL g908 ( 
.A(n_832),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_737),
.Y(n_909)
);

INVxp33_ASAP7_75t_SL g910 ( 
.A(n_758),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_773),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_776),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_742),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_792),
.Y(n_914)
);

INVxp33_ASAP7_75t_SL g915 ( 
.A(n_818),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_750),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_765),
.Y(n_917)
);

INVxp33_ASAP7_75t_SL g918 ( 
.A(n_669),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_766),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_769),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_771),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_778),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_833),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_780),
.Y(n_924)
);

NOR2xp67_ASAP7_75t_L g925 ( 
.A(n_785),
.B(n_0),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_794),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_797),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_800),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_805),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_703),
.Y(n_930)
);

INVxp67_ASAP7_75t_SL g931 ( 
.A(n_703),
.Y(n_931)
);

INVx1_ASAP7_75t_SL g932 ( 
.A(n_665),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_807),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_808),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_860),
.B(n_873),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_882),
.B(n_810),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_849),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_883),
.Y(n_938)
);

INVx4_ASAP7_75t_L g939 ( 
.A(n_880),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_850),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_848),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_932),
.A2(n_685),
.B1(n_815),
.B2(n_710),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_884),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_839),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_897),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_890),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_834),
.Y(n_947)
);

NAND2xp33_ASAP7_75t_L g948 ( 
.A(n_912),
.B(n_740),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_932),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_911),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_840),
.A2(n_672),
.B1(n_814),
.B2(n_812),
.Y(n_951)
);

OAI21x1_ASAP7_75t_L g952 ( 
.A1(n_865),
.A2(n_828),
.B(n_825),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_909),
.Y(n_953)
);

INVx4_ASAP7_75t_L g954 ( 
.A(n_917),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_903),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_835),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_930),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_857),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_836),
.Y(n_959)
);

CKINVDCx11_ASAP7_75t_R g960 ( 
.A(n_923),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_856),
.B(n_858),
.Y(n_961)
);

CKINVDCx8_ASAP7_75t_R g962 ( 
.A(n_908),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_918),
.B(n_829),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_931),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_837),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_892),
.B(n_661),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_838),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_841),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_842),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_861),
.B(n_679),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_843),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_844),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_934),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_867),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_868),
.Y(n_975)
);

OAI22x1_ASAP7_75t_SL g976 ( 
.A1(n_846),
.A2(n_662),
.B1(n_663),
.B2(n_659),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_869),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_871),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_874),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_928),
.B(n_709),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_933),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_872),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_845),
.A2(n_726),
.B1(n_770),
.B2(n_691),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_857),
.B(n_0),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_859),
.A2(n_707),
.B1(n_752),
.B2(n_698),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_864),
.B(n_921),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_904),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_876),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_877),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_878),
.Y(n_990)
);

OAI22x1_ASAP7_75t_R g991 ( 
.A1(n_862),
.A2(n_670),
.B1(n_671),
.B2(n_664),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_929),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_L g993 ( 
.A(n_853),
.B(n_740),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_927),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_899),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_879),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_885),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_886),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_887),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_889),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_854),
.A2(n_724),
.B1(n_756),
.B2(n_702),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_910),
.A2(n_684),
.B1(n_686),
.B2(n_682),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_891),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_893),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_899),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_866),
.B(n_692),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_896),
.Y(n_1007)
);

INVx6_ASAP7_75t_L g1008 ( 
.A(n_894),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_898),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_901),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_902),
.Y(n_1011)
);

NAND2xp33_ASAP7_75t_L g1012 ( 
.A(n_855),
.B(n_740),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_906),
.Y(n_1013)
);

INVx5_ASAP7_75t_L g1014 ( 
.A(n_895),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_913),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_916),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_875),
.B(n_709),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_919),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_920),
.B(n_709),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_922),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_943),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_SL g1022 ( 
.A(n_950),
.B(n_851),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_949),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_958),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_946),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_995),
.B(n_900),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_941),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_965),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_969),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_1005),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_972),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_974),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_974),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_977),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_941),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_947),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_938),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_980),
.B(n_852),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_1003),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_935),
.B(n_1006),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_980),
.B(n_847),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_977),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_989),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_963),
.B(n_924),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_989),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_945),
.B(n_926),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_996),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_957),
.B(n_907),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_996),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_937),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_947),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1000),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_950),
.B(n_900),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_955),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_940),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1000),
.Y(n_1056)
);

OA21x2_ASAP7_75t_L g1057 ( 
.A1(n_952),
.A2(n_907),
.B(n_925),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1009),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1009),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_953),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_939),
.B(n_881),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_984),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_956),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_964),
.B(n_915),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_956),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_973),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_942),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_981),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_1002),
.B(n_1017),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_944),
.B(n_914),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_992),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_994),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1019),
.B(n_694),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1016),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_959),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_959),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_979),
.B(n_905),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_960),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_1008),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_966),
.A2(n_804),
.B(n_740),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1020),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_975),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_967),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_979),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_967),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_968),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_968),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_983),
.Y(n_1088)
);

BUFx8_ASAP7_75t_L g1089 ( 
.A(n_961),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_982),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_988),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_990),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_997),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_998),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_999),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1004),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1007),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1010),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_954),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1011),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1001),
.B(n_696),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_978),
.B(n_863),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1013),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_1015),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1018),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_936),
.A2(n_804),
.B(n_740),
.Y(n_1106)
);

AND2x6_ASAP7_75t_L g1107 ( 
.A(n_1019),
.B(n_791),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_971),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_951),
.B(n_699),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_970),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_986),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_993),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_985),
.B(n_962),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1012),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1040),
.B(n_987),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1066),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_1037),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_1024),
.Y(n_1118)
);

AND2x2_ASAP7_75t_SL g1119 ( 
.A(n_1037),
.B(n_991),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_SL g1120 ( 
.A(n_1038),
.Y(n_1120)
);

INVx4_ASAP7_75t_SL g1121 ( 
.A(n_1107),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1111),
.B(n_948),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1079),
.B(n_1014),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1068),
.Y(n_1124)
);

BUFx8_ASAP7_75t_SL g1125 ( 
.A(n_1077),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1023),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1071),
.Y(n_1127)
);

NAND2xp33_ASAP7_75t_SL g1128 ( 
.A(n_1053),
.B(n_870),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1088),
.A2(n_976),
.B1(n_888),
.B2(n_711),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1050),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1072),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1074),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1030),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_1026),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_1041),
.B(n_1014),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1039),
.B(n_962),
.Y(n_1136)
);

NOR3xp33_ASAP7_75t_L g1137 ( 
.A(n_1054),
.B(n_712),
.C(n_706),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_1102),
.Y(n_1138)
);

CKINVDCx16_ASAP7_75t_R g1139 ( 
.A(n_1078),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1081),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1036),
.Y(n_1141)
);

BUFx4f_ASAP7_75t_L g1142 ( 
.A(n_1041),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1084),
.B(n_713),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_1036),
.Y(n_1144)
);

AND2x6_ASAP7_75t_L g1145 ( 
.A(n_1112),
.B(n_791),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1062),
.B(n_717),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1093),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1044),
.B(n_1070),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1100),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1028),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1114),
.B(n_720),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1089),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1110),
.B(n_727),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1029),
.Y(n_1154)
);

NAND2xp33_ASAP7_75t_L g1155 ( 
.A(n_1108),
.B(n_1048),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1089),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1031),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_1051),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1051),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1063),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1082),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1055),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1038),
.B(n_1),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_SL g1164 ( 
.A1(n_1067),
.A2(n_729),
.B1(n_731),
.B2(n_728),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1061),
.B(n_1064),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1086),
.B(n_1),
.Y(n_1166)
);

BUFx10_ASAP7_75t_L g1167 ( 
.A(n_1060),
.Y(n_1167)
);

AND2x6_ASAP7_75t_L g1168 ( 
.A(n_1091),
.B(n_791),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1092),
.B(n_734),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1063),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1069),
.B(n_735),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1063),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1090),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1094),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1095),
.A2(n_817),
.B1(n_804),
.B2(n_741),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1096),
.Y(n_1176)
);

AO22x2_ASAP7_75t_L g1177 ( 
.A1(n_1113),
.A2(n_10),
.B1(n_18),
.B2(n_2),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1090),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1090),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1097),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1098),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1103),
.B(n_738),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1105),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1104),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1021),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1022),
.B(n_743),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_1104),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1104),
.A2(n_817),
.B1(n_804),
.B2(n_746),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_SL g1189 ( 
.A(n_1107),
.Y(n_1189)
);

BUFx4f_ASAP7_75t_L g1190 ( 
.A(n_1032),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1099),
.B(n_745),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1025),
.A2(n_817),
.B1(n_804),
.B2(n_749),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1065),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1033),
.B(n_2),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1075),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1027),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1046),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1076),
.B(n_3),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1073),
.B(n_747),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1109),
.B(n_1101),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1035),
.Y(n_1201)
);

OAI21xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1106),
.A2(n_3),
.B(n_4),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1034),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1042),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1043),
.A2(n_783),
.B1(n_784),
.B2(n_760),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1045),
.B(n_751),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1047),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1083),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1085),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1049),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1052),
.B(n_4),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1087),
.Y(n_1212)
);

AND3x2_ASAP7_75t_L g1213 ( 
.A(n_1056),
.B(n_5),
.C(n_6),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1142),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1144),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1148),
.B(n_1058),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1115),
.B(n_1059),
.Y(n_1217)
);

OAI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1134),
.A2(n_1057),
.B1(n_761),
.B2(n_762),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1133),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1116),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1165),
.B(n_757),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1171),
.A2(n_1107),
.B1(n_1057),
.B2(n_767),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1197),
.B(n_764),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1144),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1124),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1127),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1117),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1123),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1131),
.B(n_775),
.Y(n_1229)
);

BUFx5_ASAP7_75t_L g1230 ( 
.A(n_1147),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1132),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1122),
.B(n_777),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1140),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1130),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1146),
.B(n_782),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1150),
.Y(n_1236)
);

INVxp67_ASAP7_75t_L g1237 ( 
.A(n_1118),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1162),
.Y(n_1238)
);

OAI221xp5_ASAP7_75t_L g1239 ( 
.A1(n_1128),
.A2(n_796),
.B1(n_798),
.B2(n_793),
.C(n_790),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1200),
.B(n_1154),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1157),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1149),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1161),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1174),
.B(n_801),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1119),
.B(n_802),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1138),
.B(n_803),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1176),
.B(n_811),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1180),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1181),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1183),
.B(n_813),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1185),
.B(n_819),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1152),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1203),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1204),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1178),
.B(n_822),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1207),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1178),
.B(n_826),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1179),
.B(n_5),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1179),
.B(n_1080),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1199),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1135),
.B(n_7),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1126),
.B(n_8),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1210),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1139),
.B(n_9),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1156),
.B(n_9),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1196),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1120),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1155),
.B(n_10),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1153),
.B(n_1143),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1198),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1170),
.B(n_11),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1190),
.B(n_11),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1201),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1136),
.B(n_12),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1164),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1275)
);

NAND3xp33_ASAP7_75t_L g1276 ( 
.A(n_1137),
.B(n_13),
.C(n_14),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1158),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1173),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1184),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1163),
.B(n_15),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1193),
.B(n_15),
.Y(n_1281)
);

CKINVDCx11_ASAP7_75t_R g1282 ( 
.A(n_1167),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1158),
.B(n_16),
.Y(n_1283)
);

NOR2xp67_ASAP7_75t_L g1284 ( 
.A(n_1160),
.B(n_138),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1177),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1159),
.B(n_17),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1159),
.B(n_20),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1151),
.B(n_20),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1141),
.B(n_21),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1195),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1209),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1187),
.B(n_22),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1172),
.B(n_23),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1214),
.B(n_1129),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1216),
.B(n_1212),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1240),
.B(n_1166),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1237),
.A2(n_1205),
.B1(n_1194),
.B2(n_1211),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1219),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1228),
.B(n_1121),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1220),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1225),
.Y(n_1301)
);

OR2x6_ASAP7_75t_L g1302 ( 
.A(n_1267),
.B(n_1195),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1227),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1215),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1226),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1215),
.B(n_1121),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1231),
.B(n_1208),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1252),
.B(n_1208),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1224),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1233),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1280),
.B(n_1169),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1236),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1241),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1277),
.B(n_1186),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1217),
.B(n_1182),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1243),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1256),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1224),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1261),
.B(n_1206),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1269),
.A2(n_1274),
.B1(n_1246),
.B2(n_1235),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1248),
.B(n_1191),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1242),
.Y(n_1322)
);

OR2x6_ASAP7_75t_L g1323 ( 
.A(n_1265),
.B(n_1189),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1288),
.A2(n_1202),
.B(n_1175),
.C(n_1192),
.Y(n_1324)
);

INVx5_ASAP7_75t_L g1325 ( 
.A(n_1264),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1249),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1282),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1253),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1270),
.B(n_1223),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1245),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1254),
.B(n_1263),
.Y(n_1331)
);

INVx5_ASAP7_75t_L g1332 ( 
.A(n_1291),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1289),
.B(n_1125),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1239),
.B(n_1213),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1234),
.B(n_1145),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1281),
.B(n_1145),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1238),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1262),
.B(n_1229),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1266),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1271),
.B(n_1145),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1244),
.B(n_1188),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1273),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1221),
.B(n_1278),
.Y(n_1343)
);

NAND2x1p5_ASAP7_75t_L g1344 ( 
.A(n_1272),
.B(n_1168),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1258),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1279),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1247),
.B(n_1168),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1285),
.A2(n_1230),
.B1(n_1275),
.B2(n_1251),
.Y(n_1348)
);

BUFx4f_ASAP7_75t_L g1349 ( 
.A(n_1276),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1230),
.A2(n_1168),
.B1(n_26),
.B2(n_24),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1230),
.B(n_24),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1292),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1250),
.B(n_25),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1255),
.Y(n_1354)
);

OR2x6_ASAP7_75t_L g1355 ( 
.A(n_1283),
.B(n_28),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1290),
.B(n_29),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1293),
.Y(n_1357)
);

INVx4_ASAP7_75t_L g1358 ( 
.A(n_1230),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1268),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1257),
.B(n_29),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1286),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1287),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1232),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1259),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1260),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1284),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1222),
.B(n_30),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1309),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1311),
.A2(n_1218),
.B1(n_32),
.B2(n_30),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1309),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1299),
.B(n_128),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1295),
.B(n_31),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1308),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_1323),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1300),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1327),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1303),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1298),
.B(n_31),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1306),
.B(n_129),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1304),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_1318),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1302),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1320),
.B(n_32),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1302),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1296),
.B(n_33),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1329),
.B(n_1354),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1294),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1332),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1338),
.B(n_33),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1315),
.B(n_34),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1317),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1301),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1332),
.B(n_130),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1331),
.B(n_34),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1330),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_L g1396 ( 
.A(n_1348),
.B(n_35),
.C(n_36),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1325),
.B(n_35),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1333),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1322),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1305),
.Y(n_1400)
);

OR2x6_ASAP7_75t_L g1401 ( 
.A(n_1323),
.B(n_36),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1310),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1364),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1314),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_1325),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1312),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1342),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1313),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1316),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1343),
.Y(n_1410)
);

AOI22x1_ASAP7_75t_L g1411 ( 
.A1(n_1365),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1326),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1339),
.Y(n_1413)
);

O2A1O1Ixp5_ASAP7_75t_L g1414 ( 
.A1(n_1319),
.A2(n_41),
.B(n_38),
.C(n_39),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1328),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1307),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1337),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1355),
.B(n_41),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1345),
.B(n_42),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1346),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1359),
.B(n_42),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1321),
.Y(n_1422)
);

NOR2xp67_ASAP7_75t_L g1423 ( 
.A(n_1353),
.B(n_131),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1362),
.Y(n_1424)
);

NOR4xp25_ASAP7_75t_SL g1425 ( 
.A(n_1351),
.B(n_1357),
.C(n_1324),
.D(n_1361),
.Y(n_1425)
);

NOR3xp33_ASAP7_75t_L g1426 ( 
.A(n_1334),
.B(n_43),
.C(n_44),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_1349),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1336),
.B(n_43),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1355),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1367),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1360),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1340),
.B(n_47),
.Y(n_1432)
);

BUFx12f_ASAP7_75t_L g1433 ( 
.A(n_1340),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1297),
.B(n_48),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1363),
.B(n_48),
.Y(n_1435)
);

NAND2x1p5_ASAP7_75t_L g1436 ( 
.A(n_1335),
.B(n_1358),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1356),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1364),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1352),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1366),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1341),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1344),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1347),
.B(n_49),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1350),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1300),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1309),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1298),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1295),
.B(n_49),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1295),
.B(n_51),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1387),
.B(n_51),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1391),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1386),
.B(n_52),
.Y(n_1452)
);

NAND3xp33_ASAP7_75t_SL g1453 ( 
.A(n_1426),
.B(n_53),
.C(n_54),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1443),
.A2(n_136),
.B(n_134),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1396),
.A2(n_54),
.B(n_55),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1432),
.A2(n_56),
.B(n_57),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1439),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1447),
.Y(n_1458)
);

BUFx4_ASAP7_75t_SL g1459 ( 
.A(n_1427),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1441),
.A2(n_141),
.B(n_139),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1422),
.B(n_58),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1425),
.A2(n_59),
.B(n_60),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1437),
.B(n_59),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_SL g1464 ( 
.A1(n_1434),
.A2(n_60),
.B(n_61),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1390),
.B(n_61),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1389),
.A2(n_62),
.B(n_63),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1378),
.B(n_62),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1377),
.B(n_63),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1407),
.B(n_64),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1418),
.B(n_64),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1383),
.A2(n_65),
.B(n_66),
.Y(n_1471)
);

AO31x2_ASAP7_75t_L g1472 ( 
.A1(n_1369),
.A2(n_144),
.A3(n_145),
.B(n_143),
.Y(n_1472)
);

OA21x2_ASAP7_75t_L g1473 ( 
.A1(n_1414),
.A2(n_65),
.B(n_66),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1375),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1392),
.B(n_67),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1416),
.B(n_69),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1400),
.B(n_69),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1402),
.B(n_70),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1398),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1376),
.Y(n_1480)
);

AND2x2_ASAP7_75t_SL g1481 ( 
.A(n_1374),
.B(n_70),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1373),
.B(n_71),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_1395),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1444),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1406),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1430),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_1486)
);

NAND2x1_ASAP7_75t_L g1487 ( 
.A(n_1408),
.B(n_146),
.Y(n_1487)
);

AOI211x1_ASAP7_75t_L g1488 ( 
.A1(n_1372),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_1488)
);

BUFx12f_ASAP7_75t_L g1489 ( 
.A(n_1401),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1409),
.A2(n_149),
.B(n_147),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1394),
.A2(n_75),
.B(n_77),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1412),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1415),
.A2(n_151),
.B(n_150),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1445),
.B(n_78),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1405),
.B(n_152),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1399),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1397),
.B(n_79),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1424),
.A2(n_1411),
.B(n_1436),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1385),
.A2(n_79),
.B(n_80),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1423),
.A2(n_80),
.B(n_81),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1416),
.B(n_81),
.Y(n_1501)
);

AOI221x1_ASAP7_75t_L g1502 ( 
.A1(n_1448),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.C(n_85),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1442),
.A2(n_156),
.B(n_155),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1421),
.A2(n_1428),
.B(n_1449),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1403),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1432),
.A2(n_1403),
.B(n_1435),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1410),
.B(n_82),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1419),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1431),
.B(n_86),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1429),
.A2(n_88),
.B(n_89),
.Y(n_1510)
);

INVx5_ASAP7_75t_L g1511 ( 
.A(n_1401),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1440),
.A2(n_159),
.B(n_157),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1404),
.B(n_89),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1381),
.B(n_90),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1382),
.B(n_90),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1368),
.B(n_91),
.Y(n_1516)
);

NAND3x1_ASAP7_75t_L g1517 ( 
.A(n_1370),
.B(n_91),
.C(n_92),
.Y(n_1517)
);

AO21x1_ASAP7_75t_L g1518 ( 
.A1(n_1379),
.A2(n_92),
.B(n_93),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1446),
.B(n_93),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1433),
.Y(n_1520)
);

NAND2x1_ASAP7_75t_L g1521 ( 
.A(n_1379),
.B(n_160),
.Y(n_1521)
);

AOI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1384),
.A2(n_167),
.B(n_164),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1388),
.B(n_94),
.Y(n_1523)
);

AND3x4_ASAP7_75t_L g1524 ( 
.A(n_1371),
.B(n_94),
.C(n_95),
.Y(n_1524)
);

NOR2x1_ASAP7_75t_SL g1525 ( 
.A(n_1417),
.B(n_96),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1380),
.B(n_96),
.Y(n_1526)
);

AO31x2_ASAP7_75t_L g1527 ( 
.A1(n_1420),
.A2(n_169),
.A3(n_170),
.B(n_168),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1413),
.B(n_97),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1438),
.B(n_97),
.Y(n_1529)
);

AO32x2_ASAP7_75t_L g1530 ( 
.A1(n_1393),
.A2(n_1371),
.A3(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1393),
.A2(n_98),
.B(n_99),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1425),
.A2(n_100),
.B(n_101),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1443),
.A2(n_172),
.B(n_171),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1391),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1386),
.B(n_101),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1407),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1443),
.A2(n_174),
.B(n_173),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1398),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1407),
.Y(n_1539)
);

INVx6_ASAP7_75t_SL g1540 ( 
.A(n_1401),
.Y(n_1540)
);

OAI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1396),
.A2(n_102),
.B(n_103),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1386),
.B(n_103),
.Y(n_1542)
);

AO21x1_ASAP7_75t_L g1543 ( 
.A1(n_1434),
.A2(n_104),
.B(n_105),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1386),
.B(n_105),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1391),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1425),
.A2(n_106),
.B(n_107),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1443),
.A2(n_176),
.B(n_175),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1443),
.A2(n_178),
.B(n_177),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1407),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1447),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1396),
.A2(n_106),
.B(n_108),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1407),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1407),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1398),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1386),
.B(n_108),
.Y(n_1555)
);

OAI21xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1430),
.A2(n_109),
.B(n_110),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1386),
.B(n_109),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1387),
.B(n_110),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1396),
.A2(n_111),
.B(n_112),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1458),
.Y(n_1560)
);

INVx4_ASAP7_75t_L g1561 ( 
.A(n_1511),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1474),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1518),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1485),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1550),
.B(n_113),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1536),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1492),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1505),
.B(n_114),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1539),
.B(n_114),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1549),
.B(n_115),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1497),
.B(n_115),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1470),
.B(n_116),
.Y(n_1572)
);

CKINVDCx8_ASAP7_75t_R g1573 ( 
.A(n_1511),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1504),
.A2(n_117),
.B(n_118),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1552),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_SL g1576 ( 
.A1(n_1453),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1538),
.B(n_1554),
.Y(n_1577)
);

AOI22x1_ASAP7_75t_L g1578 ( 
.A1(n_1466),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1467),
.B(n_120),
.Y(n_1579)
);

BUFx2_ASAP7_75t_SL g1580 ( 
.A(n_1480),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1553),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1479),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1483),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1475),
.B(n_121),
.Y(n_1584)
);

OR2x6_ASAP7_75t_L g1585 ( 
.A(n_1489),
.B(n_1506),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1452),
.B(n_122),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1535),
.B(n_122),
.Y(n_1587)
);

INVx5_ASAP7_75t_L g1588 ( 
.A(n_1479),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1530),
.B(n_123),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1451),
.Y(n_1590)
);

NAND2x1p5_ASAP7_75t_L g1591 ( 
.A(n_1520),
.B(n_179),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1496),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1542),
.B(n_123),
.Y(n_1593)
);

INVx4_ASAP7_75t_L g1594 ( 
.A(n_1482),
.Y(n_1594)
);

BUFx4f_ASAP7_75t_L g1595 ( 
.A(n_1520),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1534),
.B(n_180),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1519),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1544),
.B(n_124),
.Y(n_1598)
);

CKINVDCx16_ASAP7_75t_R g1599 ( 
.A(n_1513),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1545),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1510),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1540),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1555),
.B(n_125),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1528),
.B(n_181),
.Y(n_1604)
);

O2A1O1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1457),
.A2(n_126),
.B(n_183),
.C(n_182),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1516),
.B(n_184),
.Y(n_1606)
);

NOR2x1_ASAP7_75t_R g1607 ( 
.A(n_1459),
.B(n_186),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1501),
.B(n_187),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1507),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1469),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_R g1611 ( 
.A(n_1481),
.B(n_1522),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1476),
.B(n_1523),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1477),
.Y(n_1613)
);

NAND2x1p5_ASAP7_75t_L g1614 ( 
.A(n_1521),
.B(n_189),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1557),
.B(n_190),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_SL g1616 ( 
.A(n_1461),
.B(n_192),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1478),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1525),
.B(n_193),
.Y(n_1618)
);

O2A1O1Ixp5_ASAP7_75t_L g1619 ( 
.A1(n_1455),
.A2(n_197),
.B(n_194),
.C(n_195),
.Y(n_1619)
);

BUFx4f_ASAP7_75t_SL g1620 ( 
.A(n_1450),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1494),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1463),
.B(n_199),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1495),
.Y(n_1623)
);

OR2x6_ASAP7_75t_L g1624 ( 
.A(n_1456),
.B(n_1531),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1524),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1468),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1541),
.A2(n_200),
.B(n_202),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1526),
.B(n_203),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1529),
.Y(n_1629)
);

NOR2x1_ASAP7_75t_SL g1630 ( 
.A(n_1558),
.B(n_204),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1509),
.B(n_205),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1498),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1530),
.B(n_1515),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1488),
.B(n_206),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1465),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1514),
.B(n_207),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1508),
.Y(n_1637)
);

OR2x6_ASAP7_75t_L g1638 ( 
.A(n_1462),
.B(n_209),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1487),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1543),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1551),
.A2(n_210),
.B(n_211),
.Y(n_1641)
);

INVx3_ASAP7_75t_SL g1642 ( 
.A(n_1473),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1559),
.A2(n_212),
.B(n_214),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1464),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1471),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1517),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1502),
.B(n_219),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1527),
.B(n_220),
.Y(n_1648)
);

CKINVDCx8_ASAP7_75t_R g1649 ( 
.A(n_1556),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1527),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1491),
.B(n_1499),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1503),
.B(n_221),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1484),
.B(n_222),
.Y(n_1653)
);

NAND2xp33_ASAP7_75t_L g1654 ( 
.A(n_1486),
.B(n_1532),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1546),
.A2(n_225),
.B(n_226),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1472),
.B(n_228),
.Y(n_1656)
);

NAND2x1p5_ASAP7_75t_L g1657 ( 
.A(n_1454),
.B(n_229),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1472),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1500),
.B(n_230),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1577),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1566),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1560),
.B(n_1490),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1575),
.B(n_1548),
.Y(n_1663)
);

A2O1A1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1628),
.A2(n_1537),
.B(n_1547),
.C(n_1533),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1599),
.B(n_1493),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1581),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1562),
.Y(n_1667)
);

AO22x2_ASAP7_75t_L g1668 ( 
.A1(n_1633),
.A2(n_1512),
.B1(n_1460),
.B2(n_233),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1635),
.B(n_654),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1609),
.B(n_231),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1595),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1600),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1564),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1588),
.B(n_232),
.Y(n_1674)
);

CKINVDCx11_ASAP7_75t_R g1675 ( 
.A(n_1583),
.Y(n_1675)
);

O2A1O1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1576),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1567),
.B(n_1617),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1609),
.B(n_653),
.Y(n_1678)
);

INVx8_ASAP7_75t_L g1679 ( 
.A(n_1588),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1585),
.B(n_239),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1571),
.B(n_652),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1627),
.A2(n_240),
.B(n_242),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1582),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1613),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1573),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1585),
.B(n_243),
.Y(n_1686)
);

A2O1A1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1605),
.A2(n_246),
.B(n_244),
.C(n_245),
.Y(n_1687)
);

NAND2x1p5_ASAP7_75t_L g1688 ( 
.A(n_1623),
.B(n_248),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1572),
.B(n_651),
.Y(n_1689)
);

NOR2xp67_ASAP7_75t_L g1690 ( 
.A(n_1561),
.B(n_249),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1579),
.B(n_650),
.Y(n_1691)
);

O2A1O1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1651),
.A2(n_252),
.B(n_250),
.C(n_251),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1654),
.A2(n_253),
.B(n_254),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1621),
.B(n_649),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1641),
.A2(n_255),
.B(n_256),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1610),
.B(n_257),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1590),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1592),
.Y(n_1698)
);

OR2x6_ASAP7_75t_SL g1699 ( 
.A(n_1626),
.B(n_258),
.Y(n_1699)
);

A2O1A1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1643),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1658),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1569),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1589),
.B(n_648),
.Y(n_1703)
);

INVx3_ASAP7_75t_L g1704 ( 
.A(n_1597),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1594),
.B(n_262),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1629),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1565),
.B(n_646),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1602),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1570),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1629),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1597),
.B(n_263),
.Y(n_1711)
);

OA21x2_ASAP7_75t_L g1712 ( 
.A1(n_1632),
.A2(n_265),
.B(n_267),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1650),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1640),
.B(n_644),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1645),
.A2(n_1624),
.B(n_1619),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1642),
.Y(n_1716)
);

OA21x2_ASAP7_75t_L g1717 ( 
.A1(n_1644),
.A2(n_268),
.B(n_269),
.Y(n_1717)
);

NAND2x1p5_ASAP7_75t_L g1718 ( 
.A(n_1596),
.B(n_271),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1586),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1612),
.Y(n_1720)
);

NOR2xp67_ASAP7_75t_L g1721 ( 
.A(n_1598),
.B(n_272),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1648),
.Y(n_1722)
);

OR2x6_ASAP7_75t_SL g1723 ( 
.A(n_1637),
.B(n_275),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1568),
.B(n_642),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1634),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1584),
.B(n_276),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1624),
.A2(n_277),
.B(n_280),
.Y(n_1727)
);

OR2x6_ASAP7_75t_SL g1728 ( 
.A(n_1587),
.B(n_281),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1604),
.B(n_282),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1580),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1606),
.B(n_283),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1649),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1601),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1656),
.Y(n_1734)
);

A2O1A1Ixp33_ASAP7_75t_SL g1735 ( 
.A1(n_1639),
.A2(n_293),
.B(n_291),
.C(n_292),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1593),
.Y(n_1736)
);

A2O1A1Ixp33_ASAP7_75t_SL g1737 ( 
.A1(n_1574),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_1737)
);

O2A1O1Ixp5_ASAP7_75t_L g1738 ( 
.A1(n_1646),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1625),
.B(n_639),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1603),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1625),
.B(n_300),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1608),
.B(n_301),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1616),
.B(n_304),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1611),
.B(n_638),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1647),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1618),
.Y(n_1746)
);

NAND2x1p5_ASAP7_75t_L g1747 ( 
.A(n_1652),
.B(n_305),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1638),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1630),
.B(n_307),
.Y(n_1749)
);

A2O1A1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1563),
.A2(n_310),
.B(n_308),
.C(n_309),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1615),
.B(n_637),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1620),
.A2(n_315),
.B1(n_312),
.B2(n_313),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1578),
.Y(n_1753)
);

BUFx10_ASAP7_75t_L g1754 ( 
.A(n_1607),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1636),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1631),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1657),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1622),
.B(n_319),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1638),
.B(n_320),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1591),
.B(n_1659),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1614),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1653),
.B(n_321),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1655),
.A2(n_322),
.B(n_323),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1560),
.B(n_636),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1560),
.B(n_324),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1575),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1575),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1560),
.B(n_635),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1560),
.B(n_325),
.Y(n_1769)
);

AOI211xp5_ASAP7_75t_L g1770 ( 
.A1(n_1576),
.A2(n_330),
.B(n_326),
.C(n_329),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1575),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1560),
.B(n_331),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1583),
.Y(n_1773)
);

OA21x2_ASAP7_75t_L g1774 ( 
.A1(n_1658),
.A2(n_332),
.B(n_333),
.Y(n_1774)
);

INVxp67_ASAP7_75t_L g1775 ( 
.A(n_1635),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1575),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1625),
.B(n_334),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1560),
.B(n_336),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1560),
.B(n_634),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1575),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1560),
.B(n_338),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1651),
.A2(n_339),
.B(n_340),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1560),
.B(n_633),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1560),
.B(n_341),
.Y(n_1784)
);

NAND2x1p5_ASAP7_75t_L g1785 ( 
.A(n_1588),
.B(n_342),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1560),
.B(n_343),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1575),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1775),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1677),
.Y(n_1789)
);

AO31x2_ASAP7_75t_L g1790 ( 
.A1(n_1701),
.A2(n_348),
.A3(n_346),
.B(n_347),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1660),
.B(n_349),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1716),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1661),
.Y(n_1793)
);

OAI21x1_ASAP7_75t_L g1794 ( 
.A1(n_1715),
.A2(n_350),
.B(n_351),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1684),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1666),
.Y(n_1796)
);

INVx4_ASAP7_75t_L g1797 ( 
.A(n_1679),
.Y(n_1797)
);

BUFx3_ASAP7_75t_L g1798 ( 
.A(n_1675),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_1773),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1671),
.Y(n_1800)
);

AO22x1_ASAP7_75t_L g1801 ( 
.A1(n_1748),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1766),
.B(n_355),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1767),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1697),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1771),
.B(n_356),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1776),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1672),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1723),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1734),
.A2(n_364),
.B1(n_360),
.B2(n_361),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1698),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1780),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1787),
.B(n_1662),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1665),
.B(n_365),
.Y(n_1813)
);

CKINVDCx14_ASAP7_75t_R g1814 ( 
.A(n_1699),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1667),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1730),
.B(n_1708),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1679),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1673),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1663),
.Y(n_1819)
);

OA21x2_ASAP7_75t_L g1820 ( 
.A1(n_1745),
.A2(n_366),
.B(n_367),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1719),
.B(n_368),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1725),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1702),
.Y(n_1823)
);

AO31x2_ASAP7_75t_L g1824 ( 
.A1(n_1713),
.A2(n_373),
.A3(n_369),
.B(n_372),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1710),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1709),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1736),
.Y(n_1827)
);

BUFx3_ASAP7_75t_L g1828 ( 
.A(n_1685),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1720),
.B(n_375),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1740),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1722),
.Y(n_1831)
);

AO21x2_ASAP7_75t_L g1832 ( 
.A1(n_1744),
.A2(n_376),
.B(n_377),
.Y(n_1832)
);

AOI21x1_ASAP7_75t_L g1833 ( 
.A1(n_1714),
.A2(n_1668),
.B(n_1717),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1756),
.B(n_379),
.Y(n_1834)
);

BUFx3_ASAP7_75t_L g1835 ( 
.A(n_1704),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1682),
.A2(n_381),
.B(n_382),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1706),
.Y(n_1837)
);

INVx2_ASAP7_75t_SL g1838 ( 
.A(n_1683),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1765),
.B(n_385),
.Y(n_1839)
);

INVx1_ASAP7_75t_SL g1840 ( 
.A(n_1670),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1668),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1746),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1757),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1774),
.Y(n_1844)
);

INVx1_ASAP7_75t_SL g1845 ( 
.A(n_1678),
.Y(n_1845)
);

CKINVDCx6p67_ASAP7_75t_R g1846 ( 
.A(n_1754),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1669),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1694),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1774),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1769),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1712),
.Y(n_1851)
);

AO31x2_ASAP7_75t_L g1852 ( 
.A1(n_1664),
.A2(n_388),
.A3(n_386),
.B(n_387),
.Y(n_1852)
);

INVxp33_ASAP7_75t_L g1853 ( 
.A(n_1681),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1778),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1712),
.Y(n_1855)
);

AO21x2_ASAP7_75t_L g1856 ( 
.A1(n_1696),
.A2(n_389),
.B(n_390),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1728),
.B(n_391),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1717),
.Y(n_1858)
);

AO21x2_ASAP7_75t_L g1859 ( 
.A1(n_1721),
.A2(n_1703),
.B(n_1707),
.Y(n_1859)
);

BUFx3_ASAP7_75t_L g1860 ( 
.A(n_1711),
.Y(n_1860)
);

INVx3_ASAP7_75t_L g1861 ( 
.A(n_1772),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1753),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1761),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1764),
.Y(n_1864)
);

OAI21x1_ASAP7_75t_L g1865 ( 
.A1(n_1738),
.A2(n_392),
.B(n_393),
.Y(n_1865)
);

BUFx2_ASAP7_75t_L g1866 ( 
.A(n_1768),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1741),
.B(n_394),
.Y(n_1867)
);

AND2x4_ASAP7_75t_SL g1868 ( 
.A(n_1674),
.B(n_395),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1783),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1779),
.Y(n_1870)
);

BUFx4f_ASAP7_75t_L g1871 ( 
.A(n_1739),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1786),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1689),
.B(n_396),
.Y(n_1873)
);

INVx2_ASAP7_75t_SL g1874 ( 
.A(n_1781),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1828),
.Y(n_1875)
);

AOI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1841),
.A2(n_1733),
.B1(n_1762),
.B2(n_1759),
.Y(n_1876)
);

NAND3xp33_ASAP7_75t_L g1877 ( 
.A(n_1862),
.B(n_1770),
.C(n_1676),
.Y(n_1877)
);

AO31x2_ASAP7_75t_L g1878 ( 
.A1(n_1822),
.A2(n_1760),
.A3(n_1687),
.B(n_1784),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1808),
.A2(n_1686),
.B1(n_1680),
.B2(n_1691),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1818),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1866),
.B(n_1705),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1822),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1866),
.B(n_1724),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1859),
.A2(n_1820),
.B1(n_1870),
.B2(n_1864),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1827),
.B(n_1726),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1826),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1830),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1792),
.B(n_1743),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1823),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1815),
.Y(n_1890)
);

OAI21xp5_ASAP7_75t_SL g1891 ( 
.A1(n_1814),
.A2(n_1777),
.B(n_1693),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1838),
.B(n_1729),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1795),
.B(n_1751),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1810),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1796),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1803),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1788),
.B(n_1747),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1798),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1819),
.B(n_1758),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1804),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1848),
.B(n_1727),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1806),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1843),
.Y(n_1903)
);

AO31x2_ASAP7_75t_L g1904 ( 
.A1(n_1858),
.A2(n_1700),
.A3(n_1732),
.B(n_1750),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1792),
.B(n_1731),
.Y(n_1905)
);

BUFx2_ASAP7_75t_L g1906 ( 
.A(n_1812),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1850),
.B(n_1692),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1811),
.Y(n_1908)
);

OAI21xp5_ASAP7_75t_SL g1909 ( 
.A1(n_1857),
.A2(n_1752),
.B(n_1695),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1789),
.Y(n_1910)
);

INVx4_ASAP7_75t_L g1911 ( 
.A(n_1817),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1800),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1874),
.B(n_1782),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1793),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1846),
.B(n_1742),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1807),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1812),
.Y(n_1917)
);

OR2x6_ASAP7_75t_L g1918 ( 
.A(n_1797),
.B(n_1785),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1816),
.B(n_1853),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1831),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1842),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1854),
.B(n_1749),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1863),
.Y(n_1923)
);

AOI222xp33_ASAP7_75t_L g1924 ( 
.A1(n_1801),
.A2(n_1755),
.B1(n_1737),
.B2(n_1690),
.C1(n_1735),
.C2(n_1718),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1847),
.B(n_1688),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1869),
.B(n_1872),
.Y(n_1926)
);

AO31x2_ASAP7_75t_L g1927 ( 
.A1(n_1844),
.A2(n_1763),
.A3(n_400),
.B(n_397),
.Y(n_1927)
);

BUFx2_ASAP7_75t_L g1928 ( 
.A(n_1835),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1837),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1861),
.B(n_399),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1825),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1840),
.B(n_401),
.Y(n_1932)
);

AO31x2_ASAP7_75t_L g1933 ( 
.A1(n_1849),
.A2(n_404),
.A3(n_402),
.B(n_403),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1833),
.Y(n_1934)
);

BUFx2_ASAP7_75t_L g1935 ( 
.A(n_1799),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1805),
.B(n_406),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1845),
.B(n_407),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1851),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1860),
.B(n_408),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1855),
.Y(n_1940)
);

AND2x4_ASAP7_75t_L g1941 ( 
.A(n_1805),
.B(n_631),
.Y(n_1941)
);

INVxp67_ASAP7_75t_L g1942 ( 
.A(n_1813),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1802),
.B(n_410),
.Y(n_1943)
);

INVx3_ASAP7_75t_L g1944 ( 
.A(n_1871),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_SL g1945 ( 
.A1(n_1820),
.A2(n_413),
.B1(n_411),
.B2(n_412),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1833),
.B(n_414),
.Y(n_1946)
);

INVxp67_ASAP7_75t_SL g1947 ( 
.A(n_1834),
.Y(n_1947)
);

AND2x4_ASAP7_75t_L g1948 ( 
.A(n_1791),
.B(n_630),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1821),
.Y(n_1949)
);

NAND3xp33_ASAP7_75t_L g1950 ( 
.A(n_1934),
.B(n_1836),
.C(n_1839),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1882),
.B(n_1880),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1938),
.Y(n_1952)
);

OAI22xp33_ASAP7_75t_L g1953 ( 
.A1(n_1907),
.A2(n_1867),
.B1(n_1829),
.B2(n_1852),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1908),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1929),
.B(n_1883),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1906),
.B(n_1873),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1890),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1887),
.Y(n_1958)
);

AO21x2_ASAP7_75t_L g1959 ( 
.A1(n_1946),
.A2(n_1794),
.B(n_1832),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1940),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1900),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1889),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1917),
.B(n_1881),
.Y(n_1963)
);

AND2x2_ASAP7_75t_SL g1964 ( 
.A(n_1928),
.B(n_1868),
.Y(n_1964)
);

BUFx2_ASAP7_75t_L g1965 ( 
.A(n_1935),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1901),
.B(n_1852),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1895),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1916),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1903),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1888),
.B(n_1852),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1919),
.B(n_1865),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1896),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1921),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1905),
.B(n_1856),
.Y(n_1974)
);

NOR4xp25_ASAP7_75t_SL g1975 ( 
.A(n_1891),
.B(n_1801),
.C(n_1790),
.D(n_1809),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1902),
.B(n_1790),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1875),
.B(n_1790),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1942),
.B(n_1824),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1892),
.B(n_1824),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1885),
.B(n_1824),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1898),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1920),
.Y(n_1982)
);

NAND2x1_ASAP7_75t_L g1983 ( 
.A(n_1944),
.B(n_1893),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1894),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1914),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1899),
.B(n_415),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1886),
.Y(n_1987)
);

BUFx3_ASAP7_75t_L g1988 ( 
.A(n_1912),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1922),
.B(n_416),
.Y(n_1989)
);

AOI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1877),
.A2(n_420),
.B1(n_417),
.B2(n_418),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1931),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1923),
.Y(n_1992)
);

NOR2x1_ASAP7_75t_L g1993 ( 
.A(n_1911),
.B(n_421),
.Y(n_1993)
);

AOI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1949),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1897),
.B(n_425),
.Y(n_1995)
);

INVx3_ASAP7_75t_L g1996 ( 
.A(n_1878),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1963),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1954),
.B(n_1947),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1962),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1962),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1965),
.B(n_1878),
.Y(n_2001)
);

NOR2xp67_ASAP7_75t_L g2002 ( 
.A(n_1996),
.B(n_1884),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1996),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1967),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1971),
.B(n_1915),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1991),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1952),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1956),
.B(n_1918),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1981),
.B(n_1913),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1983),
.B(n_1918),
.Y(n_2010)
);

INVx1_ASAP7_75t_SL g2011 ( 
.A(n_1964),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1974),
.B(n_1970),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1967),
.Y(n_2013)
);

BUFx2_ASAP7_75t_L g2014 ( 
.A(n_1954),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1960),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1955),
.B(n_1925),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_1972),
.Y(n_2017)
);

AND2x2_ASAP7_75t_SL g2018 ( 
.A(n_1977),
.B(n_1876),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1973),
.Y(n_2019)
);

INVxp33_ASAP7_75t_L g2020 ( 
.A(n_1993),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1972),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1961),
.Y(n_2022)
);

BUFx2_ASAP7_75t_L g2023 ( 
.A(n_1988),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1951),
.B(n_1926),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1957),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1958),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1968),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1984),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1984),
.Y(n_2029)
);

INVxp67_ASAP7_75t_SL g2030 ( 
.A(n_1966),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1987),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_1992),
.B(n_1910),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1977),
.B(n_1879),
.Y(n_2033)
);

OR2x2_ASAP7_75t_L g2034 ( 
.A(n_1992),
.B(n_1932),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1987),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1953),
.B(n_1909),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1979),
.B(n_1930),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_2023),
.B(n_1950),
.Y(n_2038)
);

AO21x2_ASAP7_75t_L g2039 ( 
.A1(n_2002),
.A2(n_1976),
.B(n_1978),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2017),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_2025),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_2010),
.B(n_2011),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2005),
.B(n_1975),
.Y(n_2043)
);

INVxp67_ASAP7_75t_L g2044 ( 
.A(n_2036),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_2003),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_2008),
.B(n_1959),
.Y(n_2046)
);

INVxp67_ASAP7_75t_L g2047 ( 
.A(n_2009),
.Y(n_2047)
);

OAI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_2020),
.A2(n_1986),
.B1(n_1980),
.B2(n_1989),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_2024),
.B(n_1995),
.Y(n_2049)
);

INVx2_ASAP7_75t_SL g2050 ( 
.A(n_1997),
.Y(n_2050)
);

INVx5_ASAP7_75t_L g2051 ( 
.A(n_2001),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1999),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2030),
.B(n_1985),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2016),
.B(n_2012),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2014),
.B(n_1937),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1999),
.Y(n_2056)
);

BUFx2_ASAP7_75t_L g2057 ( 
.A(n_2001),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2025),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2026),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2026),
.Y(n_2060)
);

AOI31xp33_ASAP7_75t_L g2061 ( 
.A1(n_1998),
.A2(n_1924),
.A3(n_1990),
.B(n_1936),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_2034),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2000),
.Y(n_2063)
);

INVxp67_ASAP7_75t_SL g2064 ( 
.A(n_2033),
.Y(n_2064)
);

AOI211x1_ASAP7_75t_L g2065 ( 
.A1(n_2004),
.A2(n_1939),
.B(n_1904),
.C(n_1945),
.Y(n_2065)
);

NOR2x1p5_ASAP7_75t_L g2066 ( 
.A(n_2042),
.B(n_2033),
.Y(n_2066)
);

INVx2_ASAP7_75t_SL g2067 ( 
.A(n_2051),
.Y(n_2067)
);

INVx1_ASAP7_75t_SL g2068 ( 
.A(n_2055),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_2062),
.B(n_2013),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_2050),
.B(n_2021),
.Y(n_2070)
);

NOR2x1p5_ASAP7_75t_SL g2071 ( 
.A(n_2045),
.B(n_2029),
.Y(n_2071)
);

HB1xp67_ASAP7_75t_L g2072 ( 
.A(n_2057),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_2049),
.Y(n_2073)
);

BUFx2_ASAP7_75t_L g2074 ( 
.A(n_2047),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_2051),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2054),
.B(n_2028),
.Y(n_2076)
);

NOR2xp33_ASAP7_75t_L g2077 ( 
.A(n_2044),
.B(n_2037),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2038),
.B(n_2031),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_2041),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2052),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_2053),
.B(n_2040),
.Y(n_2081)
);

OR2x6_ASAP7_75t_L g2082 ( 
.A(n_2065),
.B(n_1941),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2052),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2076),
.B(n_2046),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2079),
.Y(n_2085)
);

NOR2x1_ASAP7_75t_L g2086 ( 
.A(n_2074),
.B(n_2061),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_2068),
.B(n_2064),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2072),
.B(n_2058),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_2066),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2073),
.B(n_2059),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2067),
.Y(n_2091)
);

AOI22xp5_ASAP7_75t_L g2092 ( 
.A1(n_2082),
.A2(n_2018),
.B1(n_2043),
.B2(n_2048),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2080),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2083),
.Y(n_2094)
);

OAI21xp33_ASAP7_75t_L g2095 ( 
.A1(n_2071),
.A2(n_2060),
.B(n_2063),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2069),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2078),
.B(n_2051),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2077),
.B(n_2039),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2081),
.Y(n_2099)
);

OR2x2_ASAP7_75t_L g2100 ( 
.A(n_2070),
.B(n_2056),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2087),
.B(n_2075),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2084),
.B(n_2082),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2097),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2085),
.Y(n_2104)
);

NAND2x1p5_ASAP7_75t_L g2105 ( 
.A(n_2086),
.B(n_1948),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2099),
.B(n_2056),
.Y(n_2106)
);

OAI31xp33_ASAP7_75t_L g2107 ( 
.A1(n_2095),
.A2(n_2029),
.A3(n_2000),
.B(n_2006),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2089),
.B(n_2035),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2099),
.B(n_2091),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2100),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_2092),
.B(n_2032),
.Y(n_2111)
);

HB1xp67_ASAP7_75t_L g2112 ( 
.A(n_2096),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2088),
.Y(n_2113)
);

CKINVDCx16_ASAP7_75t_R g2114 ( 
.A(n_2090),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2098),
.B(n_2019),
.Y(n_2115)
);

INVx1_ASAP7_75t_SL g2116 ( 
.A(n_2114),
.Y(n_2116)
);

HB1xp67_ASAP7_75t_L g2117 ( 
.A(n_2109),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2112),
.Y(n_2118)
);

OA21x2_ASAP7_75t_L g2119 ( 
.A1(n_2101),
.A2(n_2094),
.B(n_2093),
.Y(n_2119)
);

INVx3_ASAP7_75t_SL g2120 ( 
.A(n_2103),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2102),
.B(n_2027),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2110),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_2105),
.Y(n_2123)
);

INVxp67_ASAP7_75t_L g2124 ( 
.A(n_2108),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2113),
.B(n_2007),
.Y(n_2125)
);

INVxp67_ASAP7_75t_L g2126 ( 
.A(n_2104),
.Y(n_2126)
);

OR2x2_ASAP7_75t_L g2127 ( 
.A(n_2113),
.B(n_2022),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2117),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2116),
.B(n_2107),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2119),
.Y(n_2130)
);

AOI322xp5_ASAP7_75t_L g2131 ( 
.A1(n_2122),
.A2(n_2111),
.A3(n_2115),
.B1(n_2106),
.B2(n_2015),
.C1(n_1969),
.C2(n_1982),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2120),
.B(n_1904),
.Y(n_2132)
);

O2A1O1Ixp33_ASAP7_75t_L g2133 ( 
.A1(n_2119),
.A2(n_1943),
.B(n_1994),
.C(n_1927),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2121),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2124),
.B(n_1927),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2118),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2125),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2127),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2134),
.B(n_2126),
.Y(n_2139)
);

OAI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_2130),
.A2(n_2123),
.B1(n_1933),
.B2(n_428),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2128),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_SL g2142 ( 
.A(n_2137),
.B(n_1933),
.Y(n_2142)
);

INVx2_ASAP7_75t_SL g2143 ( 
.A(n_2138),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2136),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2135),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2129),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_2132),
.Y(n_2147)
);

INVx3_ASAP7_75t_L g2148 ( 
.A(n_2131),
.Y(n_2148)
);

NOR3xp33_ASAP7_75t_L g2149 ( 
.A(n_2133),
.B(n_426),
.C(n_427),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2130),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2134),
.B(n_429),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2134),
.Y(n_2152)
);

BUFx8_ASAP7_75t_SL g2153 ( 
.A(n_2152),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2150),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2143),
.B(n_430),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2139),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2146),
.B(n_432),
.Y(n_2157)
);

NOR2xp33_ASAP7_75t_L g2158 ( 
.A(n_2144),
.B(n_434),
.Y(n_2158)
);

BUFx2_ASAP7_75t_L g2159 ( 
.A(n_2141),
.Y(n_2159)
);

OAI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_2148),
.A2(n_438),
.B1(n_435),
.B2(n_437),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2151),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2147),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2149),
.B(n_439),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2145),
.Y(n_2164)
);

AOI22xp5_ASAP7_75t_L g2165 ( 
.A1(n_2161),
.A2(n_2140),
.B1(n_2142),
.B2(n_443),
.Y(n_2165)
);

AOI221xp5_ASAP7_75t_L g2166 ( 
.A1(n_2154),
.A2(n_440),
.B1(n_442),
.B2(n_444),
.C(n_446),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2159),
.B(n_447),
.Y(n_2167)
);

AOI211xp5_ASAP7_75t_L g2168 ( 
.A1(n_2156),
.A2(n_451),
.B(n_449),
.C(n_450),
.Y(n_2168)
);

NAND3xp33_ASAP7_75t_L g2169 ( 
.A(n_2158),
.B(n_453),
.C(n_455),
.Y(n_2169)
);

NOR2xp67_ASAP7_75t_L g2170 ( 
.A(n_2164),
.B(n_456),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2153),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_2162),
.B(n_2155),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2157),
.B(n_458),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_2167),
.B(n_2160),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2172),
.Y(n_2175)
);

NOR3xp33_ASAP7_75t_L g2176 ( 
.A(n_2173),
.B(n_2163),
.C(n_460),
.Y(n_2176)
);

OAI221xp5_ASAP7_75t_L g2177 ( 
.A1(n_2165),
.A2(n_461),
.B1(n_463),
.B2(n_464),
.C(n_466),
.Y(n_2177)
);

AOI221xp5_ASAP7_75t_L g2178 ( 
.A1(n_2171),
.A2(n_467),
.B1(n_468),
.B2(n_470),
.C(n_471),
.Y(n_2178)
);

OR2x2_ASAP7_75t_L g2179 ( 
.A(n_2169),
.B(n_473),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2170),
.B(n_474),
.Y(n_2180)
);

NAND4xp25_ASAP7_75t_L g2181 ( 
.A(n_2168),
.B(n_475),
.C(n_476),
.D(n_477),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2166),
.Y(n_2182)
);

OAI211xp5_ASAP7_75t_L g2183 ( 
.A1(n_2171),
.A2(n_478),
.B(n_479),
.C(n_480),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2171),
.B(n_482),
.Y(n_2184)
);

AOI222xp33_ASAP7_75t_L g2185 ( 
.A1(n_2172),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.C1(n_486),
.C2(n_487),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2175),
.B(n_488),
.Y(n_2186)
);

NOR2xp67_ASAP7_75t_L g2187 ( 
.A(n_2184),
.B(n_489),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2180),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2182),
.Y(n_2189)
);

AOI22xp33_ASAP7_75t_L g2190 ( 
.A1(n_2174),
.A2(n_491),
.B1(n_493),
.B2(n_494),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2176),
.Y(n_2191)
);

AOI211xp5_ASAP7_75t_L g2192 ( 
.A1(n_2177),
.A2(n_495),
.B(n_497),
.C(n_499),
.Y(n_2192)
);

NOR3xp33_ASAP7_75t_L g2193 ( 
.A(n_2183),
.B(n_2181),
.C(n_2179),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2185),
.Y(n_2194)
);

AOI21xp5_ASAP7_75t_L g2195 ( 
.A1(n_2178),
.A2(n_500),
.B(n_502),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2175),
.B(n_503),
.Y(n_2196)
);

XNOR2xp5_ASAP7_75t_L g2197 ( 
.A(n_2184),
.B(n_504),
.Y(n_2197)
);

AOI21xp5_ASAP7_75t_L g2198 ( 
.A1(n_2175),
.A2(n_505),
.B(n_506),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2175),
.Y(n_2199)
);

O2A1O1Ixp33_ASAP7_75t_L g2200 ( 
.A1(n_2175),
.A2(n_507),
.B(n_508),
.C(n_509),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2196),
.B(n_510),
.Y(n_2201)
);

NOR2xp67_ASAP7_75t_SL g2202 ( 
.A(n_2199),
.B(n_511),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2186),
.Y(n_2203)
);

NOR3x2_ASAP7_75t_L g2204 ( 
.A(n_2189),
.B(n_512),
.C(n_513),
.Y(n_2204)
);

NOR3x1_ASAP7_75t_L g2205 ( 
.A(n_2194),
.B(n_515),
.C(n_516),
.Y(n_2205)
);

NAND3xp33_ASAP7_75t_L g2206 ( 
.A(n_2191),
.B(n_517),
.C(n_518),
.Y(n_2206)
);

NOR2x1_ASAP7_75t_L g2207 ( 
.A(n_2188),
.B(n_519),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_2193),
.B(n_520),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2197),
.B(n_522),
.Y(n_2209)
);

INVx5_ASAP7_75t_L g2210 ( 
.A(n_2187),
.Y(n_2210)
);

AND2x4_ASAP7_75t_L g2211 ( 
.A(n_2195),
.B(n_523),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2198),
.B(n_525),
.Y(n_2212)
);

NOR2x1p5_ASAP7_75t_L g2213 ( 
.A(n_2192),
.B(n_526),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_2200),
.B(n_530),
.Y(n_2214)
);

NAND2x1p5_ASAP7_75t_SL g2215 ( 
.A(n_2190),
.B(n_531),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2199),
.B(n_532),
.Y(n_2216)
);

NOR3xp33_ASAP7_75t_L g2217 ( 
.A(n_2199),
.B(n_533),
.C(n_536),
.Y(n_2217)
);

NAND3xp33_ASAP7_75t_L g2218 ( 
.A(n_2199),
.B(n_537),
.C(n_538),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_2199),
.B(n_540),
.Y(n_2219)
);

BUFx2_ASAP7_75t_L g2220 ( 
.A(n_2199),
.Y(n_2220)
);

BUFx2_ASAP7_75t_L g2221 ( 
.A(n_2220),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_2203),
.B(n_541),
.Y(n_2222)
);

XNOR2xp5_ASAP7_75t_L g2223 ( 
.A(n_2213),
.B(n_542),
.Y(n_2223)
);

AOI221xp5_ASAP7_75t_L g2224 ( 
.A1(n_2214),
.A2(n_545),
.B1(n_546),
.B2(n_547),
.C(n_548),
.Y(n_2224)
);

AOI221xp5_ASAP7_75t_L g2225 ( 
.A1(n_2208),
.A2(n_550),
.B1(n_551),
.B2(n_552),
.C(n_553),
.Y(n_2225)
);

NOR2x2_ASAP7_75t_L g2226 ( 
.A(n_2205),
.B(n_554),
.Y(n_2226)
);

NOR2x1_ASAP7_75t_L g2227 ( 
.A(n_2219),
.B(n_555),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_2210),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2216),
.B(n_557),
.Y(n_2229)
);

NAND3xp33_ASAP7_75t_SL g2230 ( 
.A(n_2217),
.B(n_558),
.C(n_559),
.Y(n_2230)
);

OR2x2_ASAP7_75t_L g2231 ( 
.A(n_2215),
.B(n_560),
.Y(n_2231)
);

NOR2x1_ASAP7_75t_L g2232 ( 
.A(n_2207),
.B(n_561),
.Y(n_2232)
);

NOR2x1_ASAP7_75t_L g2233 ( 
.A(n_2218),
.B(n_563),
.Y(n_2233)
);

BUFx3_ASAP7_75t_L g2234 ( 
.A(n_2221),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2226),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2231),
.Y(n_2236)
);

NAND4xp75_ASAP7_75t_L g2237 ( 
.A(n_2232),
.B(n_2209),
.C(n_2212),
.D(n_2201),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2223),
.B(n_2210),
.Y(n_2238)
);

NAND4xp75_ASAP7_75t_L g2239 ( 
.A(n_2227),
.B(n_2202),
.C(n_2204),
.D(n_2206),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2228),
.Y(n_2240)
);

AO22x2_ASAP7_75t_L g2241 ( 
.A1(n_2229),
.A2(n_2211),
.B1(n_565),
.B2(n_566),
.Y(n_2241)
);

INVx3_ASAP7_75t_L g2242 ( 
.A(n_2225),
.Y(n_2242)
);

OAI221xp5_ASAP7_75t_L g2243 ( 
.A1(n_2234),
.A2(n_2224),
.B1(n_2233),
.B2(n_2222),
.C(n_2230),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2241),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2237),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2235),
.Y(n_2246)
);

OAI221xp5_ASAP7_75t_SL g2247 ( 
.A1(n_2245),
.A2(n_2240),
.B1(n_2238),
.B2(n_2236),
.C(n_2242),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2244),
.Y(n_2248)
);

XOR2xp5_ASAP7_75t_L g2249 ( 
.A(n_2248),
.B(n_2246),
.Y(n_2249)
);

NOR2x1p5_ASAP7_75t_L g2250 ( 
.A(n_2247),
.B(n_2239),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2249),
.B(n_2243),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2250),
.Y(n_2252)
);

NAND3xp33_ASAP7_75t_SL g2253 ( 
.A(n_2252),
.B(n_564),
.C(n_567),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2251),
.Y(n_2254)
);

OAI22xp5_ASAP7_75t_SL g2255 ( 
.A1(n_2254),
.A2(n_569),
.B1(n_570),
.B2(n_571),
.Y(n_2255)
);

OAI21xp5_ASAP7_75t_L g2256 ( 
.A1(n_2253),
.A2(n_572),
.B(n_573),
.Y(n_2256)
);

HB1xp67_ASAP7_75t_L g2257 ( 
.A(n_2256),
.Y(n_2257)
);

OR2x2_ASAP7_75t_L g2258 ( 
.A(n_2255),
.B(n_574),
.Y(n_2258)
);

OA21x2_ASAP7_75t_L g2259 ( 
.A1(n_2257),
.A2(n_575),
.B(n_578),
.Y(n_2259)
);

AO21x1_ASAP7_75t_L g2260 ( 
.A1(n_2258),
.A2(n_579),
.B(n_581),
.Y(n_2260)
);

AOI21xp5_ASAP7_75t_L g2261 ( 
.A1(n_2257),
.A2(n_583),
.B(n_584),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2257),
.B(n_585),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2260),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2262),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2259),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2261),
.Y(n_2266)
);

OR2x6_ASAP7_75t_L g2267 ( 
.A(n_2265),
.B(n_586),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2263),
.B(n_588),
.Y(n_2268)
);

OR2x6_ASAP7_75t_L g2269 ( 
.A(n_2264),
.B(n_589),
.Y(n_2269)
);

AOI21xp5_ASAP7_75t_L g2270 ( 
.A1(n_2267),
.A2(n_2266),
.B(n_590),
.Y(n_2270)
);

AOI211xp5_ASAP7_75t_L g2271 ( 
.A1(n_2270),
.A2(n_2268),
.B(n_2269),
.C(n_592),
.Y(n_2271)
);


endmodule