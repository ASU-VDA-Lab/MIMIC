module fake_jpeg_1553_n_208 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_208);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_14),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_SL g66 ( 
.A(n_0),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_33),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_7),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_79),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_2),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_92),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_66),
.B1(n_52),
.B2(n_67),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_56),
.B1(n_64),
.B2(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_83),
.B(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_104),
.Y(n_120)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_54),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_58),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_67),
.B(n_66),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_115),
.B(n_114),
.Y(n_127)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_60),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_61),
.B1(n_68),
.B2(n_69),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_68),
.B1(n_74),
.B2(n_9),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_61),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_20),
.Y(n_136)
);

OA22x2_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_62),
.B1(n_74),
.B2(n_73),
.Y(n_115)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_115),
.A2(n_74),
.A3(n_62),
.B1(n_89),
.B2(n_73),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_70),
.C(n_65),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_62),
.Y(n_126)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_89),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_134),
.B1(n_117),
.B2(n_100),
.Y(n_142)
);

OR2x2_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_62),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_127),
.B(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_71),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_125),
.B(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_74),
.B(n_5),
.Y(n_129)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_107),
.B(n_105),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_34),
.B(n_32),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_4),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_132),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_116),
.B(n_4),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_101),
.B(n_5),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_137),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_22),
.B1(n_48),
.B2(n_47),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_7),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_21),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_178)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_147),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_8),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_156),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_25),
.C(n_44),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_157),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_19),
.Y(n_152)
);

A2O1A1O1Ixp25_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_155),
.B(n_16),
.C(n_17),
.D(n_18),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_49),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_10),
.C(n_11),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_41),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_39),
.C(n_38),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_8),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_159),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_9),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_28),
.B(n_26),
.Y(n_172)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_18),
.B(n_141),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_130),
.B1(n_118),
.B2(n_12),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_166),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_149),
.C(n_154),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_171),
.C(n_157),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_30),
.C(n_29),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_178),
.B(n_181),
.Y(n_190)
);

AO22x1_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_174)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

AO22x2_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_180),
.B(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_182),
.B(n_168),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_189),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_177),
.B(n_158),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_176),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_161),
.C(n_152),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_192),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_173),
.B(n_155),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_179),
.B1(n_144),
.B2(n_170),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_196),
.Y(n_197)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_189),
.C(n_182),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_200),
.A2(n_194),
.B(n_185),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_201),
.A2(n_202),
.B(n_199),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_174),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_200),
.C(n_197),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_203),
.A2(n_204),
.B1(n_190),
.B2(n_144),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_175),
.C(n_180),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g207 ( 
.A(n_206),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_172),
.Y(n_208)
);


endmodule