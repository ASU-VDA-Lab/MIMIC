module fake_jpeg_27205_n_250 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_SL g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_30),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_16),
.Y(n_50)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_35),
.B1(n_41),
.B2(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_51),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_18),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_21),
.B1(n_27),
.B2(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_21),
.B1(n_27),
.B2(n_31),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_60),
.C(n_43),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_31),
.B1(n_23),
.B2(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_63),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_19),
.C(n_24),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_34),
.A2(n_23),
.B1(n_32),
.B2(n_20),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_65),
.B(n_73),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_22),
.B(n_33),
.C(n_29),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_67),
.A2(n_29),
.B(n_52),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_70),
.B(n_76),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_25),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_25),
.Y(n_78)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_43),
.C(n_38),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_25),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_93),
.Y(n_128)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_56),
.B1(n_60),
.B2(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_94),
.B(n_104),
.Y(n_132)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_99),
.Y(n_137)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_57),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_103),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_49),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_52),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_55),
.B1(n_46),
.B2(n_52),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_109),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_55),
.B1(n_46),
.B2(n_38),
.Y(n_109)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_83),
.C(n_71),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_121),
.C(n_91),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_122),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_74),
.B(n_66),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_2),
.B(n_3),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_74),
.C(n_66),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_85),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_134),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_70),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_129),
.Y(n_155)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_85),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_86),
.B(n_37),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_64),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_136),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_107),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_90),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_105),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_121),
.C(n_131),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_110),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_140),
.B(n_141),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_91),
.B(n_67),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_95),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_132),
.A2(n_69),
.B1(n_76),
.B2(n_46),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_154),
.B1(n_130),
.B2(n_123),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_106),
.B(n_97),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_160),
.B(n_125),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_97),
.B1(n_99),
.B2(n_68),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_145),
.A2(n_152),
.B1(n_161),
.B2(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_75),
.C(n_15),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_153),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_150),
.B(n_158),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_68),
.B1(n_88),
.B2(n_89),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_89),
.B1(n_113),
.B2(n_93),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_43),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_159),
.B(n_162),
.Y(n_173)
);

HAxp5_ASAP7_75t_SL g160 ( 
.A(n_115),
.B(n_19),
.CON(n_160),
.SN(n_160)
);

XNOR2x1_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_136),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_136),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_172),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_167),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_170),
.C(n_179),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_157),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_114),
.C(n_122),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_175),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_114),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_176),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_162),
.B(n_127),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_153),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_128),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_116),
.C(n_129),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_181),
.A2(n_148),
.B1(n_149),
.B2(n_156),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_123),
.C(n_124),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_183),
.C(n_152),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_124),
.C(n_38),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_169),
.A2(n_134),
.B1(n_98),
.B2(n_92),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_198),
.B1(n_44),
.B2(n_3),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_154),
.B1(n_148),
.B2(n_155),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_188),
.A2(n_196),
.B1(n_197),
.B2(n_175),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_190),
.B(n_2),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_200),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_201),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_172),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_144),
.B1(n_140),
.B2(n_160),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_128),
.B1(n_113),
.B2(n_92),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_168),
.B1(n_182),
.B2(n_179),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_26),
.B1(n_24),
.B2(n_19),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_26),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_44),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_206),
.B1(n_211),
.B2(n_197),
.Y(n_220)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_209),
.B1(n_196),
.B2(n_7),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_173),
.B1(n_44),
.B2(n_26),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_14),
.C(n_4),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_212),
.C(n_213),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_14),
.C(n_5),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_4),
.C(n_5),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_4),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_214),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_205),
.B(n_191),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_218),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_193),
.C(n_184),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_220),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_188),
.C(n_191),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_223),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_185),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_222),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_200),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_224),
.A2(n_6),
.B(n_7),
.Y(n_231)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_215),
.B(n_208),
.CI(n_213),
.CON(n_226),
.SN(n_226)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_230),
.Y(n_233)
);

INVx11_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_231),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_203),
.B(n_212),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_227),
.A2(n_217),
.B1(n_216),
.B2(n_9),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_217),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_237),
.Y(n_241)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_230),
.A2(n_6),
.B(n_7),
.Y(n_238)
);

AOI21xp33_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_6),
.B(n_9),
.Y(n_240)
);

AO221x1_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_226),
.B1(n_228),
.B2(n_225),
.C(n_232),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_239),
.A2(n_236),
.B(n_233),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_237),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_233),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_245),
.B1(n_242),
.B2(n_226),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_232),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_246),
.B(n_10),
.Y(n_249)
);

XNOR2x2_ASAP7_75t_SL g250 ( 
.A(n_249),
.B(n_12),
.Y(n_250)
);


endmodule