module real_jpeg_25332_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_1),
.A2(n_27),
.B1(n_39),
.B2(n_42),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_1),
.A2(n_27),
.B1(n_51),
.B2(n_52),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_1),
.A2(n_27),
.B1(n_67),
.B2(n_68),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_3),
.A2(n_51),
.B1(n_52),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_3),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_3),
.A2(n_67),
.B1(n_68),
.B2(n_85),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_39),
.B1(n_42),
.B2(n_85),
.Y(n_134)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_7),
.A2(n_67),
.B1(n_68),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_72),
.Y(n_126)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_39),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_9),
.A2(n_49),
.B1(n_67),
.B2(n_68),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_10),
.A2(n_39),
.B1(n_42),
.B2(n_58),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_36),
.B1(n_58),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_58),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_10),
.A2(n_58),
.B1(n_67),
.B2(n_68),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_11),
.B(n_30),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_11),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_11),
.B(n_38),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_11),
.B(n_52),
.C(n_54),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_11),
.A2(n_39),
.B1(n_42),
.B2(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_11),
.B(n_109),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_159),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_11),
.B(n_67),
.C(n_80),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_11),
.A2(n_69),
.B(n_218),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_12),
.A2(n_36),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_12),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_12),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_12),
.A2(n_44),
.B1(n_67),
.B2(n_68),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_14),
.A2(n_67),
.B1(n_68),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_14),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_15),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_15),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_15),
.A2(n_51),
.B1(n_52),
.B2(n_66),
.Y(n_94)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_16),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_144),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_142),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_20),
.B(n_121),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_86),
.C(n_98),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_21),
.A2(n_22),
.B1(n_86),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_62),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_46),
.B2(n_47),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_25),
.B(n_46),
.C(n_62),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_38),
.B2(n_43),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_26),
.Y(n_100)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g111 ( 
.A1(n_31),
.A2(n_35),
.A3(n_42),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_31),
.A2(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_32),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_32),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_32),
.A2(n_139),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_42),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_34),
.B(n_39),
.Y(n_113)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_37),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_37),
.B(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_42),
.B1(n_54),
.B2(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_39),
.B(n_184),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_43),
.Y(n_136)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B(n_56),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_48),
.A2(n_50),
.B1(n_60),
.B2(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_50),
.A2(n_56),
.B(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_52),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_52),
.B(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_57),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_59),
.A2(n_107),
.B1(n_109),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_60),
.A2(n_106),
.B(n_108),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_60),
.A2(n_108),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_76),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_63),
.B(n_76),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_115),
.B1(n_116),
.B2(n_118),
.Y(n_114)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_70),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_68),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_68),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_71),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_73),
.B(n_88),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_69),
.A2(n_117),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_69),
.B(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_69),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_70),
.Y(n_219)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_75),
.B(n_159),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_77),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_77),
.A2(n_206),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_94),
.B1(n_95),
.B2(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_78),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_78),
.A2(n_95),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_82),
.A2(n_83),
.B(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_82),
.A2(n_155),
.B(n_191),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_82),
.B(n_159),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_86),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_91),
.A2(n_115),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_95),
.B(n_156),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_98),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.C(n_110),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_99),
.B(n_105),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_110),
.B(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_114),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_118),
.A2(n_186),
.B(n_187),
.Y(n_185)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_141),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_140),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_130),
.Y(n_140)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B(n_138),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_176),
.B(n_260),
.C(n_265),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_170),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_170),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_161),
.C(n_162),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_147),
.A2(n_148),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_157),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_153),
.C(n_157),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_161),
.B(n_162),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_167),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_200),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_169),
.A2(n_231),
.B(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_171),
.B(n_174),
.C(n_175),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_254),
.B(n_259),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_207),
.B(n_253),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_196),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_181),
.B(n_196),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_189),
.C(n_193),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_182),
.B(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_185),
.Y(n_203)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_189),
.A2(n_193),
.B1(n_194),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_197),
.B(n_203),
.C(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_247),
.B(n_252),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_227),
.B(n_246),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_221),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_221),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_215),
.C(n_216),
.Y(n_251)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_225),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_235),
.B(n_245),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_233),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_240),
.B(n_244),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_258),
.Y(n_259)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);


endmodule