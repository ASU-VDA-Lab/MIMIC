module fake_jpeg_7854_n_172 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_21),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_31),
.A2(n_29),
.B1(n_22),
.B2(n_25),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_29),
.B1(n_22),
.B2(n_25),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_45),
.B1(n_38),
.B2(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_47),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_38),
.B1(n_39),
.B2(n_29),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_30),
.B1(n_20),
.B2(n_16),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_31),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_66),
.B1(n_70),
.B2(n_43),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_63),
.B1(n_43),
.B2(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_20),
.B1(n_30),
.B2(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_23),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_73),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_30),
.B1(n_31),
.B2(n_16),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_23),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_8),
.C(n_14),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_47),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_75),
.B(n_79),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_56),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_62),
.B(n_71),
.C(n_18),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_54),
.B1(n_41),
.B2(n_37),
.Y(n_99)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_84),
.Y(n_103)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_87),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_83),
.B1(n_64),
.B2(n_46),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_46),
.B1(n_41),
.B2(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_51),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_51),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_104),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_79),
.B(n_85),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_84),
.B1(n_75),
.B2(n_86),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_105),
.B1(n_77),
.B2(n_26),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_87),
.B1(n_19),
.B2(n_78),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_62),
.B(n_37),
.C(n_26),
.D(n_51),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_26),
.B1(n_69),
.B2(n_2),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_76),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_69),
.C(n_27),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_19),
.C(n_27),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_86),
.C(n_78),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_121),
.C(n_107),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_81),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_118),
.B1(n_123),
.B2(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_89),
.C(n_8),
.Y(n_121)
);

NOR2xp67_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_0),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_122),
.A2(n_124),
.B1(n_101),
.B2(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_1),
.Y(n_124)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_126),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_135),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_111),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_136),
.B(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_140),
.B(n_136),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_143),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_127),
.C(n_133),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_117),
.B1(n_102),
.B2(n_105),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_142),
.A2(n_146),
.B1(n_1),
.B2(n_2),
.Y(n_152)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_145),
.B(n_128),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_117),
.B1(n_105),
.B2(n_97),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_153),
.C(n_151),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_139),
.A2(n_135),
.B(n_105),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_146),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_144),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_154),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_152),
.B(n_142),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_2),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_3),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_155),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_4),
.B(n_5),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_158),
.B(n_159),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_153),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_160),
.B(n_7),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_157),
.B(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_162),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_165),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_156),
.B1(n_6),
.B2(n_7),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_5),
.C(n_7),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_170),
.C(n_168),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_167),
.Y(n_172)
);


endmodule