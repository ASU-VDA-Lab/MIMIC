module fake_netlist_1_10697_n_642 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_642);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_642;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_494;
wire n_223;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_20), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_55), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_59), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_4), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_57), .Y(n_90) );
INVx2_ASAP7_75t_SL g91 ( .A(n_17), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_46), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_43), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_4), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_38), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_75), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_8), .Y(n_97) );
INVx3_ASAP7_75t_L g98 ( .A(n_45), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_66), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_36), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_64), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_3), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_10), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_44), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_77), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_39), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_9), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_6), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_35), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_62), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_1), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_50), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_23), .Y(n_113) );
INVx3_ASAP7_75t_L g114 ( .A(n_13), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_56), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_33), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_8), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_18), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_0), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_28), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_10), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_12), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_34), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_7), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_12), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_27), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_7), .Y(n_127) );
INVxp67_ASAP7_75t_SL g128 ( .A(n_81), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_30), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_51), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_114), .Y(n_132) );
INVx6_ASAP7_75t_L g133 ( .A(n_113), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_99), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_114), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_91), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_92), .B(n_2), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_114), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_114), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_98), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_125), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_125), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_98), .B(n_3), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_125), .B(n_5), .Y(n_144) );
INVx4_ASAP7_75t_L g145 ( .A(n_98), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_125), .B(n_5), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_87), .B(n_6), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_91), .B(n_9), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_97), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_113), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_91), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_87), .B(n_11), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_97), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_97), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_93), .B(n_11), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_119), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_151), .B(n_88), .Y(n_159) );
OR2x6_ASAP7_75t_L g160 ( .A(n_148), .B(n_89), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
NAND2x1p5_ASAP7_75t_L g162 ( .A(n_144), .B(n_88), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_144), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_133), .Y(n_164) );
INVx4_ASAP7_75t_L g165 ( .A(n_145), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_141), .B(n_95), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_148), .B(n_96), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_150), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_142), .B(n_95), .Y(n_170) );
NAND2xp33_ASAP7_75t_L g171 ( .A(n_146), .B(n_100), .Y(n_171) );
OR2x2_ASAP7_75t_L g172 ( .A(n_137), .B(n_146), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_132), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_132), .B(n_113), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_150), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_133), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_131), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_144), .B(n_119), .Y(n_179) );
INVxp67_ASAP7_75t_SL g180 ( .A(n_135), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_131), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_148), .B(n_123), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_138), .B(n_104), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_138), .B(n_119), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_139), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_133), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_140), .Y(n_188) );
INVx5_ASAP7_75t_L g189 ( .A(n_165), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_160), .B(n_136), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_160), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_172), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_182), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_160), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_160), .A2(n_143), .B1(n_147), .B2(n_152), .Y(n_195) );
NAND2x1p5_ASAP7_75t_L g196 ( .A(n_165), .B(n_139), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_172), .A2(n_155), .B(n_156), .C(n_154), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_172), .B(n_165), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_168), .B(n_134), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_160), .A2(n_108), .B1(n_89), .B2(n_94), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
BUFx2_ASAP7_75t_L g202 ( .A(n_160), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_183), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_163), .A2(n_133), .B1(n_140), .B2(n_118), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_182), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_163), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_162), .B(n_104), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_180), .A2(n_109), .B(n_101), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_164), .Y(n_209) );
NAND3xp33_ASAP7_75t_SL g210 ( .A(n_162), .B(n_134), .C(n_115), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_182), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_182), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_180), .B(n_101), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_162), .B(n_105), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
NAND2x1p5_ASAP7_75t_L g216 ( .A(n_163), .B(n_105), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_173), .B(n_109), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_182), .Y(n_218) );
NAND2xp33_ASAP7_75t_L g219 ( .A(n_163), .B(n_93), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_179), .B(n_94), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_182), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_164), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_182), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_178), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_179), .B(n_106), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_179), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_173), .B(n_149), .Y(n_227) );
BUFx2_ASAP7_75t_L g228 ( .A(n_184), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_178), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_178), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_192), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_200), .A2(n_167), .B(n_159), .C(n_184), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_215), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_228), .B(n_171), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_SL g235 ( .A1(n_208), .A2(n_159), .B(n_167), .C(n_175), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_203), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_191), .B(n_158), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_215), .A2(n_130), .B1(n_161), .B2(n_158), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_215), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_190), .A2(n_161), .B1(n_181), .B2(n_186), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_215), .Y(n_241) );
AND3x1_ASAP7_75t_SL g242 ( .A(n_210), .B(n_127), .C(n_102), .Y(n_242) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_197), .A2(n_186), .B(n_181), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_191), .B(n_188), .Y(n_244) );
INVx2_ASAP7_75t_SL g245 ( .A(n_228), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_206), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_226), .B(n_185), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_194), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_219), .A2(n_170), .B(n_187), .Y(n_249) );
INVx4_ASAP7_75t_L g250 ( .A(n_189), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_208), .A2(n_170), .B(n_188), .C(n_185), .Y(n_251) );
BUFx8_ASAP7_75t_SL g252 ( .A(n_190), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_224), .Y(n_253) );
INVx4_ASAP7_75t_L g254 ( .A(n_189), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_200), .A2(n_185), .B(n_188), .C(n_154), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_206), .Y(n_256) );
INVx5_ASAP7_75t_L g257 ( .A(n_201), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_206), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_189), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_206), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_202), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_190), .A2(n_149), .B1(n_156), .B2(n_153), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_226), .B(n_187), .Y(n_263) );
AO32x2_ASAP7_75t_L g264 ( .A1(n_194), .A2(n_187), .A3(n_166), .B1(n_153), .B2(n_174), .Y(n_264) );
INVx4_ASAP7_75t_L g265 ( .A(n_189), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_202), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_189), .B(n_187), .Y(n_267) );
BUFx2_ASAP7_75t_SL g268 ( .A(n_189), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_209), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_213), .B(n_86), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_190), .A2(n_127), .B1(n_102), .B2(n_118), .Y(n_271) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_243), .A2(n_216), .B(n_193), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_245), .B(n_213), .Y(n_273) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_249), .A2(n_216), .B(n_193), .Y(n_274) );
CKINVDCx16_ASAP7_75t_R g275 ( .A(n_266), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_253), .Y(n_276) );
OAI22x1_ASAP7_75t_L g277 ( .A1(n_231), .A2(n_195), .B1(n_216), .B2(n_220), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_251), .A2(n_193), .B(n_212), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_232), .A2(n_195), .B(n_198), .Y(n_279) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_253), .A2(n_211), .B(n_218), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_244), .A2(n_211), .B(n_218), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_262), .B(n_220), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_232), .A2(n_224), .B(n_230), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_244), .A2(n_211), .B(n_218), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_252), .A2(n_220), .B1(n_199), .B2(n_225), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_236), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_252), .B(n_220), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_267), .A2(n_221), .B(n_205), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_239), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_262), .B(n_217), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_238), .B(n_217), .Y(n_291) );
OAI21xp33_ASAP7_75t_L g292 ( .A1(n_270), .A2(n_234), .B(n_255), .Y(n_292) );
OAI21xp5_ASAP7_75t_L g293 ( .A1(n_255), .A2(n_224), .B(n_230), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_246), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_256), .Y(n_295) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_235), .A2(n_240), .B(n_230), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_258), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_241), .B(n_229), .Y(n_298) );
OAI21x1_ASAP7_75t_L g299 ( .A1(n_267), .A2(n_205), .B(n_212), .Y(n_299) );
AOI21x1_ASAP7_75t_L g300 ( .A1(n_237), .A2(n_169), .B(n_174), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_247), .A2(n_227), .B1(n_196), .B2(n_201), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_261), .B(n_229), .Y(n_302) );
AO21x2_ASAP7_75t_L g303 ( .A1(n_235), .A2(n_227), .B(n_207), .Y(n_303) );
AO31x2_ASAP7_75t_L g304 ( .A1(n_271), .A2(n_157), .A3(n_169), .B(n_174), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_257), .B(n_233), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_276), .Y(n_306) );
OAI22xp33_ASAP7_75t_L g307 ( .A1(n_275), .A2(n_266), .B1(n_257), .B2(n_248), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_301), .A2(n_237), .B(n_214), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_282), .B(n_229), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_277), .A2(n_257), .B1(n_268), .B2(n_260), .Y(n_310) );
INVx11_ASAP7_75t_L g311 ( .A(n_286), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_301), .A2(n_242), .B1(n_122), .B2(n_103), .Y(n_312) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_290), .A2(n_263), .B(n_204), .Y(n_313) );
OAI22xp33_ASAP7_75t_SL g314 ( .A1(n_291), .A2(n_124), .B1(n_117), .B2(n_121), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_282), .B(n_229), .Y(n_315) );
AOI22xp33_ASAP7_75t_SL g316 ( .A1(n_275), .A2(n_257), .B1(n_265), .B2(n_259), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_277), .A2(n_265), .B1(n_259), .B2(n_254), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_276), .B(n_250), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_276), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_273), .B(n_250), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_274), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_294), .Y(n_322) );
OAI22xp5_ASAP7_75t_SL g323 ( .A1(n_287), .A2(n_111), .B1(n_108), .B2(n_107), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_280), .Y(n_324) );
OAI21x1_ASAP7_75t_SL g325 ( .A1(n_283), .A2(n_254), .B(n_201), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_279), .B(n_196), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_291), .A2(n_248), .B1(n_269), .B2(n_201), .Y(n_327) );
AOI21xp33_ASAP7_75t_L g328 ( .A1(n_292), .A2(n_248), .B(n_269), .Y(n_328) );
NOR2xp33_ASAP7_75t_SL g329 ( .A(n_305), .B(n_248), .Y(n_329) );
OR2x6_ASAP7_75t_L g330 ( .A(n_305), .B(n_196), .Y(n_330) );
OAI22x1_ASAP7_75t_SL g331 ( .A1(n_285), .A2(n_107), .B1(n_106), .B2(n_129), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_305), .Y(n_332) );
BUFx3_ASAP7_75t_L g333 ( .A(n_305), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_279), .A2(n_209), .B1(n_222), .B2(n_110), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_306), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_319), .B(n_283), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_319), .B(n_296), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_314), .B(n_289), .Y(n_338) );
BUFx2_ASAP7_75t_SL g339 ( .A(n_332), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_306), .B(n_296), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_306), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_326), .B(n_293), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_326), .B(n_293), .Y(n_343) );
INVxp67_ASAP7_75t_L g344 ( .A(n_318), .Y(n_344) );
OAI321xp33_ASAP7_75t_L g345 ( .A1(n_312), .A2(n_292), .A3(n_126), .B1(n_129), .B2(n_116), .C(n_112), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_324), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_322), .B(n_278), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_322), .B(n_294), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_321), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_332), .B(n_304), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_309), .Y(n_351) );
INVx2_ASAP7_75t_SL g352 ( .A(n_330), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_309), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_315), .B(n_295), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_324), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_315), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_332), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_318), .B(n_278), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_314), .B(n_302), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_333), .B(n_295), .Y(n_360) );
AND2x4_ASAP7_75t_SL g361 ( .A(n_330), .B(n_302), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_324), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_347), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_350), .B(n_333), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_347), .Y(n_365) );
AOI22xp33_ASAP7_75t_SL g366 ( .A1(n_338), .A2(n_323), .B1(n_333), .B2(n_329), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_342), .B(n_321), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_346), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_352), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_350), .B(n_321), .Y(n_370) );
AOI21xp5_ASAP7_75t_SL g371 ( .A1(n_352), .A2(n_330), .B(n_327), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_336), .B(n_310), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_344), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_342), .B(n_321), .Y(n_374) );
AOI33xp33_ASAP7_75t_L g375 ( .A1(n_351), .A2(n_126), .A3(n_112), .B1(n_116), .B2(n_120), .B3(n_110), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_346), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_342), .B(n_321), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_338), .B(n_323), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_336), .B(n_304), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_343), .B(n_321), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_336), .B(n_304), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_347), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_359), .A2(n_312), .B1(n_307), .B2(n_330), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_343), .B(n_304), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_350), .B(n_330), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_343), .B(n_304), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_335), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_346), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_351), .B(n_304), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_353), .B(n_303), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_352), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_355), .Y(n_393) );
BUFx8_ASAP7_75t_L g394 ( .A(n_357), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_339), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_358), .B(n_303), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_373), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_367), .B(n_358), .Y(n_398) );
BUFx2_ASAP7_75t_SL g399 ( .A(n_395), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_367), .B(n_358), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_363), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_374), .B(n_337), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_363), .B(n_353), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_374), .B(n_337), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_365), .B(n_349), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_365), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_364), .B(n_355), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_377), .B(n_337), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_382), .B(n_356), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_395), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_382), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_364), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_370), .B(n_362), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_392), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_394), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_377), .B(n_362), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_370), .B(n_385), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_385), .B(n_362), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_380), .B(n_340), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_372), .B(n_356), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_387), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_378), .B(n_311), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_394), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_368), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_387), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_392), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_393), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_380), .B(n_340), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_396), .B(n_349), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_368), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_366), .B(n_311), .Y(n_431) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_371), .B(n_339), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_393), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_372), .B(n_335), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_389), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_389), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_368), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_384), .B(n_344), .Y(n_438) );
OR2x6_ASAP7_75t_SL g439 ( .A(n_379), .B(n_360), .Y(n_439) );
OAI211xp5_ASAP7_75t_L g440 ( .A1(n_366), .A2(n_316), .B(n_359), .C(n_354), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_379), .B(n_335), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_376), .Y(n_442) );
OAI211xp5_ASAP7_75t_L g443 ( .A1(n_383), .A2(n_354), .B(n_360), .C(n_317), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_384), .B(n_340), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_398), .B(n_396), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_398), .B(n_386), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_397), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_439), .B(n_386), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_400), .B(n_381), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_401), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_415), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_421), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_406), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_411), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_439), .B(n_381), .Y(n_455) );
NOR2x1_ASAP7_75t_L g456 ( .A(n_432), .B(n_371), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_400), .B(n_376), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_402), .B(n_376), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_435), .B(n_390), .Y(n_459) );
AO221x1_ASAP7_75t_L g460 ( .A1(n_423), .A2(n_394), .B1(n_325), .B2(n_388), .C(n_341), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_414), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_417), .B(n_388), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_402), .B(n_369), .Y(n_463) );
XNOR2x2_ASAP7_75t_L g464 ( .A(n_410), .B(n_390), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_436), .B(n_369), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_404), .B(n_388), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_412), .B(n_369), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_420), .B(n_391), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_425), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_420), .B(n_391), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_431), .B(n_375), .C(n_394), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_424), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_444), .B(n_391), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_414), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_405), .B(n_357), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_417), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_426), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_444), .B(n_341), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_404), .B(n_341), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_408), .B(n_357), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_427), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g482 ( .A(n_440), .B(n_345), .C(n_120), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_408), .B(n_348), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_424), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_433), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_430), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_405), .B(n_361), .Y(n_487) );
INVx1_ASAP7_75t_SL g488 ( .A(n_415), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_438), .B(n_348), .Y(n_489) );
NAND2x1p5_ASAP7_75t_L g490 ( .A(n_407), .B(n_329), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_403), .B(n_361), .Y(n_491) );
XNOR2x1_ASAP7_75t_L g492 ( .A(n_422), .B(n_13), .Y(n_492) );
INVx3_ASAP7_75t_L g493 ( .A(n_429), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_407), .B(n_361), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_430), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_409), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_399), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_434), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_441), .B(n_14), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_441), .B(n_14), .Y(n_500) );
AOI221x1_ASAP7_75t_SL g501 ( .A1(n_405), .A2(n_331), .B1(n_93), .B2(n_17), .C(n_18), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_434), .B(n_15), .Y(n_502) );
OAI22xp33_ASAP7_75t_L g503 ( .A1(n_471), .A2(n_418), .B1(n_413), .B2(n_437), .Y(n_503) );
OAI211xp5_ASAP7_75t_L g504 ( .A1(n_456), .A2(n_443), .B(n_418), .C(n_413), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_445), .B(n_419), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_452), .Y(n_506) );
OAI221xp5_ASAP7_75t_L g507 ( .A1(n_501), .A2(n_399), .B1(n_90), .B2(n_128), .C(n_442), .Y(n_507) );
INVxp67_ASAP7_75t_L g508 ( .A(n_452), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_469), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_469), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_498), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_447), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_482), .A2(n_345), .B(n_320), .C(n_331), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_450), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_449), .B(n_419), .Y(n_515) );
AOI31xp33_ASAP7_75t_L g516 ( .A1(n_451), .A2(n_429), .A3(n_416), .B(n_428), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_455), .A2(n_428), .B1(n_429), .B2(n_416), .C(n_442), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_449), .B(n_303), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_460), .A2(n_328), .B(n_325), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_453), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_482), .A2(n_334), .B1(n_297), .B2(n_308), .Y(n_521) );
XNOR2x1_ASAP7_75t_L g522 ( .A(n_492), .B(n_15), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_448), .A2(n_297), .B1(n_313), .B2(n_166), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_472), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_496), .B(n_16), .Y(n_525) );
OAI22xp33_ASAP7_75t_L g526 ( .A1(n_497), .A2(n_298), .B1(n_264), .B2(n_300), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_502), .A2(n_298), .B(n_169), .C(n_176), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_493), .Y(n_528) );
OAI221xp5_ASAP7_75t_L g529 ( .A1(n_492), .A2(n_176), .B1(n_157), .B2(n_166), .C(n_21), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_454), .Y(n_530) );
O2A1O1Ixp5_ASAP7_75t_L g531 ( .A1(n_487), .A2(n_176), .B(n_157), .C(n_300), .Y(n_531) );
NOR2x1_ASAP7_75t_L g532 ( .A(n_488), .B(n_16), .Y(n_532) );
INVxp67_ASAP7_75t_SL g533 ( .A(n_500), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_477), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_476), .B(n_19), .Y(n_535) );
OAI21xp33_ASAP7_75t_L g536 ( .A1(n_473), .A2(n_166), .B(n_274), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_446), .B(n_19), .Y(n_537) );
INVxp67_ASAP7_75t_L g538 ( .A(n_499), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_481), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_445), .B(n_20), .Y(n_540) );
NOR3xp33_ASAP7_75t_SL g541 ( .A(n_468), .B(n_21), .C(n_22), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_483), .B(n_166), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_457), .B(n_264), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_458), .B(n_166), .Y(n_544) );
NAND2xp33_ASAP7_75t_L g545 ( .A(n_493), .B(n_166), .Y(n_545) );
OAI31xp33_ASAP7_75t_L g546 ( .A1(n_490), .A2(n_264), .A3(n_177), .B(n_164), .Y(n_546) );
INVxp67_ASAP7_75t_L g547 ( .A(n_461), .Y(n_547) );
AOI221xp5_ASAP7_75t_L g548 ( .A1(n_470), .A2(n_177), .B1(n_212), .B2(n_221), .C(n_205), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_485), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_457), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_478), .B(n_272), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_458), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_474), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_517), .B(n_466), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_505), .B(n_466), .Y(n_555) );
OAI21xp33_ASAP7_75t_L g556 ( .A1(n_516), .A2(n_463), .B(n_480), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_550), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_552), .B(n_493), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_515), .B(n_479), .Y(n_559) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_504), .A2(n_465), .B(n_467), .Y(n_560) );
OAI322xp33_ASAP7_75t_L g561 ( .A1(n_538), .A2(n_489), .A3(n_464), .B1(n_462), .B2(n_459), .C1(n_491), .C2(n_494), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_SL g562 ( .A1(n_529), .A2(n_495), .B(n_486), .C(n_484), .Y(n_562) );
XNOR2xp5_ASAP7_75t_L g563 ( .A(n_522), .B(n_487), .Y(n_563) );
AND2x4_ASAP7_75t_L g564 ( .A(n_528), .B(n_487), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_518), .B(n_495), .Y(n_565) );
NAND2x1p5_ASAP7_75t_L g566 ( .A(n_532), .B(n_475), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_506), .B(n_486), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_509), .B(n_484), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_547), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_524), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_503), .A2(n_475), .B1(n_490), .B2(n_472), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_541), .B(n_475), .C(n_464), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_547), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_510), .B(n_272), .Y(n_574) );
O2A1O1Ixp33_ASAP7_75t_L g575 ( .A1(n_507), .A2(n_222), .B(n_209), .C(n_177), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_553), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_528), .B(n_264), .Y(n_577) );
XNOR2x1_ASAP7_75t_L g578 ( .A(n_537), .B(n_24), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_533), .B(n_299), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_553), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_533), .A2(n_222), .B1(n_223), .B2(n_288), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_514), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_508), .B(n_299), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_520), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_530), .Y(n_585) );
OAI311xp33_ASAP7_75t_L g586 ( .A1(n_540), .A2(n_25), .A3(n_26), .B1(n_29), .C1(n_31), .Y(n_586) );
OAI21xp5_ASAP7_75t_SL g587 ( .A1(n_513), .A2(n_32), .B(n_37), .Y(n_587) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_545), .B(n_223), .C(n_221), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_569), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_587), .A2(n_519), .B(n_508), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_557), .Y(n_591) );
OAI221xp5_ASAP7_75t_L g592 ( .A1(n_587), .A2(n_538), .B1(n_535), .B2(n_546), .C(n_527), .Y(n_592) );
OA21x2_ASAP7_75t_L g593 ( .A1(n_572), .A2(n_512), .B(n_511), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_556), .A2(n_534), .B1(n_549), .B2(n_539), .Y(n_594) );
XNOR2xp5_ASAP7_75t_L g595 ( .A(n_563), .B(n_525), .Y(n_595) );
NAND3xp33_ASAP7_75t_SL g596 ( .A(n_566), .B(n_523), .C(n_536), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_573), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_554), .B(n_542), .Y(n_598) );
AOI221x1_ASAP7_75t_L g599 ( .A1(n_572), .A2(n_544), .B1(n_543), .B2(n_526), .C(n_531), .Y(n_599) );
OAI211xp5_ASAP7_75t_L g600 ( .A1(n_562), .A2(n_521), .B(n_551), .C(n_548), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_576), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_580), .B(n_288), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_560), .A2(n_284), .B1(n_281), .B2(n_531), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_L g604 ( .A1(n_575), .A2(n_561), .B(n_586), .C(n_585), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_582), .Y(n_605) );
OAI211xp5_ASAP7_75t_L g606 ( .A1(n_571), .A2(n_284), .B(n_281), .C(n_280), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_578), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_584), .B(n_40), .Y(n_608) );
AOI21xp33_ASAP7_75t_L g609 ( .A1(n_579), .A2(n_41), .B(n_42), .Y(n_609) );
OAI21xp33_ASAP7_75t_SL g610 ( .A1(n_558), .A2(n_47), .B(n_48), .Y(n_610) );
NOR2xp67_ASAP7_75t_L g611 ( .A(n_590), .B(n_564), .Y(n_611) );
OAI321xp33_ASAP7_75t_L g612 ( .A1(n_592), .A2(n_577), .A3(n_581), .B1(n_583), .B2(n_574), .C(n_561), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_594), .A2(n_565), .B1(n_567), .B2(n_568), .C(n_559), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_598), .A2(n_564), .B1(n_570), .B2(n_555), .Y(n_614) );
AOI321xp33_ASAP7_75t_L g615 ( .A1(n_604), .A2(n_586), .A3(n_588), .B1(n_53), .B2(n_54), .C(n_58), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_592), .A2(n_588), .B1(n_223), .B2(n_60), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_590), .A2(n_223), .B1(n_52), .B2(n_61), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_589), .B(n_49), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_605), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_595), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_610), .A2(n_223), .B1(n_65), .B2(n_67), .C(n_68), .Y(n_621) );
AOI211xp5_ASAP7_75t_L g622 ( .A1(n_600), .A2(n_223), .B(n_69), .C(n_70), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_619), .B(n_614), .Y(n_623) );
BUFx2_ASAP7_75t_L g624 ( .A(n_620), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_611), .A2(n_593), .B1(n_596), .B2(n_607), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_613), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g627 ( .A(n_612), .B(n_608), .C(n_609), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_618), .Y(n_628) );
NOR2x1_ASAP7_75t_L g629 ( .A(n_617), .B(n_593), .Y(n_629) );
NOR3xp33_ASAP7_75t_L g630 ( .A(n_624), .B(n_622), .C(n_621), .Y(n_630) );
NOR3xp33_ASAP7_75t_SL g631 ( .A(n_626), .B(n_615), .C(n_606), .Y(n_631) );
AND3x4_ASAP7_75t_L g632 ( .A(n_629), .B(n_618), .C(n_599), .Y(n_632) );
OAI221xp5_ASAP7_75t_L g633 ( .A1(n_625), .A2(n_616), .B1(n_601), .B2(n_597), .C(n_591), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_632), .A2(n_627), .B1(n_623), .B2(n_628), .Y(n_634) );
NAND4xp75_ASAP7_75t_L g635 ( .A(n_631), .B(n_603), .C(n_602), .D(n_72), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_633), .A2(n_63), .B(n_71), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_634), .A2(n_630), .B1(n_74), .B2(n_76), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_636), .B(n_73), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_637), .B(n_635), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_639), .A2(n_638), .B1(n_79), .B2(n_80), .Y(n_640) );
AOI22x1_ASAP7_75t_L g641 ( .A1(n_640), .A2(n_78), .B1(n_82), .B2(n_83), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_641), .A2(n_84), .B(n_85), .Y(n_642) );
endmodule