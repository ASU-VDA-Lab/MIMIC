module fake_aes_12_n_720 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_720);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_720;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_46), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_17), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_68), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_26), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_71), .Y(n_84) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_34), .Y(n_85) );
CKINVDCx16_ASAP7_75t_R g86 ( .A(n_15), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_0), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_76), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_56), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_47), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_22), .Y(n_91) );
BUFx3_ASAP7_75t_L g92 ( .A(n_7), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_33), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_16), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_61), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_30), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_12), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_5), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_74), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_59), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_77), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_4), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_55), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_54), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_51), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_69), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_50), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_38), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_36), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_65), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_60), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_11), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_20), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_52), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_63), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_53), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_66), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_9), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_48), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_6), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_23), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_45), .Y(n_124) );
INVxp33_ASAP7_75t_SL g125 ( .A(n_40), .Y(n_125) );
OR2x2_ASAP7_75t_L g126 ( .A(n_8), .B(n_29), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_5), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_39), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_86), .B(n_0), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_92), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_80), .B(n_1), .Y(n_132) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_127), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_92), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_127), .B(n_1), .Y(n_135) );
AND2x6_ASAP7_75t_L g136 ( .A(n_90), .B(n_28), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
AOI22xp5_ASAP7_75t_L g138 ( .A1(n_84), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_101), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_81), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_108), .B(n_3), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_113), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_113), .Y(n_143) );
INVx6_ASAP7_75t_L g144 ( .A(n_108), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_98), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_93), .Y(n_146) );
BUFx2_ASAP7_75t_L g147 ( .A(n_107), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_87), .B(n_6), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_103), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_94), .B(n_7), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_105), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_93), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_84), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_93), .B(n_8), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_106), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_109), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_93), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_97), .B(n_9), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_112), .B(n_10), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_123), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_114), .B(n_10), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_111), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_123), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_117), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_119), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_124), .Y(n_167) );
NOR2xp67_ASAP7_75t_L g168 ( .A(n_126), .B(n_11), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_116), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_82), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_123), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_85), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_133), .A2(n_125), .B1(n_110), .B2(n_104), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_134), .Y(n_174) );
INVx5_ASAP7_75t_L g175 ( .A(n_136), .Y(n_175) );
BUFx8_ASAP7_75t_SL g176 ( .A(n_153), .Y(n_176) );
OAI22xp33_ASAP7_75t_L g177 ( .A1(n_138), .A2(n_102), .B1(n_120), .B2(n_122), .Y(n_177) );
INVx4_ASAP7_75t_L g178 ( .A(n_141), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_158), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_134), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g181 ( .A1(n_147), .A2(n_110), .B1(n_104), .B2(n_85), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_170), .B(n_89), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_147), .B(n_88), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_134), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_145), .B(n_88), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_130), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_141), .B(n_139), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_158), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_167), .B(n_128), .Y(n_189) );
AND2x6_ASAP7_75t_L g190 ( .A(n_141), .B(n_125), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_158), .A2(n_100), .B1(n_115), .B2(n_128), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_158), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_161), .Y(n_193) );
AND2x6_ASAP7_75t_L g194 ( .A(n_141), .B(n_96), .Y(n_194) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_161), .B(n_96), .Y(n_195) );
INVx6_ASAP7_75t_L g196 ( .A(n_144), .Y(n_196) );
INVx1_ASAP7_75t_SL g197 ( .A(n_130), .Y(n_197) );
BUFx10_ASAP7_75t_L g198 ( .A(n_161), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_170), .B(n_121), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_161), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_146), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_167), .B(n_118), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_139), .B(n_95), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
INVx1_ASAP7_75t_SL g205 ( .A(n_135), .Y(n_205) );
NAND3xp33_ASAP7_75t_SL g206 ( .A(n_138), .B(n_99), .C(n_91), .Y(n_206) );
BUFx10_ASAP7_75t_L g207 ( .A(n_149), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_137), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_149), .B(n_83), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_137), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_151), .B(n_42), .Y(n_211) );
INVx1_ASAP7_75t_SL g212 ( .A(n_148), .Y(n_212) );
INVxp33_ASAP7_75t_L g213 ( .A(n_168), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_131), .Y(n_214) );
OR2x6_ASAP7_75t_L g215 ( .A(n_168), .B(n_13), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_151), .B(n_43), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_134), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_144), .Y(n_218) );
INVx1_ASAP7_75t_SL g219 ( .A(n_148), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_131), .Y(n_220) );
INVx4_ASAP7_75t_SL g221 ( .A(n_136), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_129), .Y(n_222) );
AND2x6_ASAP7_75t_L g223 ( .A(n_159), .B(n_44), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_169), .B(n_15), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_144), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_169), .A2(n_16), .B(n_18), .C(n_19), .Y(n_226) );
AND2x2_ASAP7_75t_SL g227 ( .A(n_159), .B(n_21), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_155), .B(n_24), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_146), .Y(n_229) );
AND3x2_ASAP7_75t_L g230 ( .A(n_132), .B(n_25), .C(n_27), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_137), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_140), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_155), .A2(n_79), .B1(n_32), .B2(n_35), .Y(n_233) );
AO22x2_ASAP7_75t_L g234 ( .A1(n_156), .A2(n_31), .B1(n_37), .B2(n_41), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_144), .Y(n_235) );
AND2x6_ASAP7_75t_L g236 ( .A(n_129), .B(n_49), .Y(n_236) );
AOI22xp33_ASAP7_75t_SL g237 ( .A1(n_227), .A2(n_150), .B1(n_140), .B2(n_143), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_181), .B(n_150), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_207), .B(n_166), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_188), .A2(n_156), .B(n_166), .C(n_165), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_217), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_207), .B(n_165), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_192), .A2(n_162), .B(n_142), .C(n_143), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_173), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_205), .B(n_162), .Y(n_245) );
AND3x1_ASAP7_75t_L g246 ( .A(n_185), .B(n_172), .C(n_142), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_204), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_198), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_199), .B(n_162), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_222), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_204), .Y(n_251) );
NAND2xp33_ASAP7_75t_L g252 ( .A(n_190), .B(n_136), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_208), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_218), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_208), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_203), .B(n_172), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_210), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_199), .B(n_182), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_176), .Y(n_260) );
INVx4_ASAP7_75t_L g261 ( .A(n_178), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_182), .B(n_129), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_177), .A2(n_154), .B(n_142), .C(n_140), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_209), .B(n_140), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_210), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_202), .B(n_143), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_202), .B(n_143), .Y(n_267) );
NAND2x1p5_ASAP7_75t_L g268 ( .A(n_227), .B(n_142), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_212), .B(n_144), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_219), .B(n_136), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_189), .B(n_136), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_191), .B(n_136), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_196), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_191), .B(n_136), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_223), .A2(n_136), .B1(n_164), .B2(n_152), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_213), .B(n_164), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_213), .B(n_164), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_197), .B(n_160), .Y(n_278) );
NAND2x1_ASAP7_75t_L g279 ( .A(n_178), .B(n_164), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_224), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_183), .B(n_160), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_223), .A2(n_160), .B1(n_152), .B2(n_171), .Y(n_282) );
BUFx3_ASAP7_75t_L g283 ( .A(n_196), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_203), .B(n_163), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_228), .B(n_163), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_193), .B(n_152), .Y(n_286) );
BUFx12f_ASAP7_75t_L g287 ( .A(n_215), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_195), .A2(n_171), .B1(n_163), .B2(n_157), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_225), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_190), .B(n_171), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_223), .A2(n_171), .B1(n_163), .B2(n_157), .Y(n_291) );
BUFx6f_ASAP7_75t_SL g292 ( .A(n_194), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_179), .B(n_171), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_214), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_186), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_190), .B(n_171), .Y(n_296) );
O2A1O1Ixp5_ASAP7_75t_L g297 ( .A1(n_187), .A2(n_163), .B(n_157), .C(n_146), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_190), .B(n_163), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_223), .A2(n_157), .B1(n_146), .B2(n_62), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_215), .B(n_57), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_179), .B(n_58), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_190), .B(n_157), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_220), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_206), .B(n_157), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_200), .B(n_146), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_271), .A2(n_187), .B(n_200), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_252), .A2(n_239), .B(n_242), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_261), .Y(n_308) );
OAI21x1_ASAP7_75t_L g309 ( .A1(n_297), .A2(n_211), .B(n_174), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_259), .B(n_195), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_294), .A2(n_228), .B(n_216), .C(n_231), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g312 ( .A1(n_240), .A2(n_180), .B(n_184), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_238), .A2(n_177), .B(n_206), .C(n_215), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_268), .A2(n_234), .B1(n_233), .B2(n_194), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_280), .B(n_194), .Y(n_315) );
NOR2x1_ASAP7_75t_L g316 ( .A(n_300), .B(n_216), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_295), .B(n_194), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_268), .A2(n_234), .B1(n_233), .B2(n_194), .Y(n_318) );
A2O1A1Ixp33_ASAP7_75t_L g319 ( .A1(n_303), .A2(n_232), .B(n_226), .C(n_211), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_285), .A2(n_175), .B(n_226), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_300), .B(n_223), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_261), .Y(n_322) );
NOR2xp33_ASAP7_75t_R g323 ( .A(n_287), .B(n_198), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_254), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_278), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_272), .A2(n_175), .B(n_235), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_262), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_248), .B(n_236), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_248), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_274), .A2(n_175), .B(n_234), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_289), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_257), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_264), .Y(n_333) );
NOR2xp33_ASAP7_75t_R g334 ( .A(n_260), .B(n_236), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_270), .A2(n_221), .B(n_229), .Y(n_335) );
NOR3xp33_ASAP7_75t_SL g336 ( .A(n_244), .B(n_176), .C(n_230), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_237), .B(n_221), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_284), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_269), .Y(n_339) );
AOI21x1_ASAP7_75t_L g340 ( .A1(n_290), .A2(n_302), .B(n_296), .Y(n_340) );
AOI22x1_ASAP7_75t_L g341 ( .A1(n_304), .A2(n_146), .B1(n_229), .B2(n_201), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_245), .B(n_196), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_286), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_247), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_237), .A2(n_236), .B1(n_221), .B2(n_230), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_286), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_249), .A2(n_229), .B(n_201), .Y(n_347) );
NOR3xp33_ASAP7_75t_L g348 ( .A(n_263), .B(n_236), .C(n_67), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_275), .B(n_229), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_288), .B(n_201), .Y(n_350) );
OAI21x1_ASAP7_75t_L g351 ( .A1(n_297), .A2(n_236), .B(n_201), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_256), .B(n_64), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_298), .A2(n_266), .B(n_267), .Y(n_353) );
NOR2xp33_ASAP7_75t_R g354 ( .A(n_292), .B(n_70), .Y(n_354) );
INVx4_ASAP7_75t_L g355 ( .A(n_292), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_275), .B(n_72), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_256), .A2(n_73), .B1(n_75), .B2(n_78), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_282), .B(n_301), .Y(n_358) );
OAI21xp33_ASAP7_75t_L g359 ( .A1(n_281), .A2(n_246), .B(n_243), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_325), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_327), .Y(n_361) );
NOR2xp33_ASAP7_75t_SL g362 ( .A(n_321), .B(n_257), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_310), .B(n_241), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_351), .A2(n_291), .B(n_282), .Y(n_364) );
A2O1A1Ixp33_ASAP7_75t_L g365 ( .A1(n_313), .A2(n_281), .B(n_276), .C(n_277), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_333), .B(n_276), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_307), .A2(n_305), .B(n_293), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_326), .A2(n_305), .B(n_293), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_310), .B(n_265), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_321), .B(n_251), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_323), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_323), .Y(n_372) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_314), .A2(n_253), .B1(n_255), .B2(n_258), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_SL g374 ( .A1(n_319), .A2(n_277), .B(n_279), .C(n_250), .Y(n_374) );
NOR2x1_ASAP7_75t_SL g375 ( .A(n_355), .B(n_257), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_352), .B(n_273), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_344), .Y(n_377) );
BUFx2_ASAP7_75t_SL g378 ( .A(n_355), .Y(n_378) );
AOI22xp33_ASAP7_75t_SL g379 ( .A1(n_318), .A2(n_283), .B1(n_291), .B2(n_299), .Y(n_379) );
O2A1O1Ixp33_ASAP7_75t_L g380 ( .A1(n_359), .A2(n_257), .B(n_299), .C(n_315), .Y(n_380) );
AO31x2_ASAP7_75t_L g381 ( .A1(n_330), .A2(n_311), .A3(n_345), .B(n_353), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_338), .Y(n_382) );
O2A1O1Ixp33_ASAP7_75t_SL g383 ( .A1(n_337), .A2(n_349), .B(n_328), .C(n_358), .Y(n_383) );
NAND3xp33_ASAP7_75t_SL g384 ( .A(n_336), .B(n_357), .C(n_317), .Y(n_384) );
A2O1A1Ixp33_ASAP7_75t_L g385 ( .A1(n_339), .A2(n_348), .B(n_306), .C(n_346), .Y(n_385) );
NOR2xp33_ASAP7_75t_SL g386 ( .A(n_316), .B(n_332), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_329), .Y(n_387) );
INVx4_ASAP7_75t_L g388 ( .A(n_332), .Y(n_388) );
OAI21x1_ASAP7_75t_L g389 ( .A1(n_347), .A2(n_341), .B(n_309), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_L g390 ( .A1(n_343), .A2(n_337), .B(n_348), .C(n_312), .Y(n_390) );
A2O1A1Ixp33_ASAP7_75t_L g391 ( .A1(n_320), .A2(n_342), .B(n_357), .C(n_324), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_L g392 ( .A1(n_358), .A2(n_349), .B(n_342), .C(n_350), .Y(n_392) );
OAI21x1_ASAP7_75t_L g393 ( .A1(n_335), .A2(n_340), .B(n_356), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_361), .B(n_329), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_371), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_377), .Y(n_396) );
OAI21x1_ASAP7_75t_L g397 ( .A1(n_389), .A2(n_393), .B(n_364), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_372), .A2(n_308), .B1(n_322), .B2(n_331), .Y(n_398) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_372), .A2(n_366), .B1(n_360), .B2(n_369), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_363), .B(n_336), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_385), .A2(n_332), .B(n_334), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_384), .A2(n_334), .B1(n_354), .B2(n_332), .Y(n_402) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_388), .B(n_354), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_381), .Y(n_404) );
AO21x2_ASAP7_75t_L g405 ( .A1(n_373), .A2(n_383), .B(n_391), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_382), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_378), .Y(n_407) );
BUFx4f_ASAP7_75t_SL g408 ( .A(n_370), .Y(n_408) );
AOI22xp33_ASAP7_75t_SL g409 ( .A1(n_362), .A2(n_386), .B1(n_375), .B2(n_376), .Y(n_409) );
INVx3_ASAP7_75t_L g410 ( .A(n_388), .Y(n_410) );
INVx4_ASAP7_75t_SL g411 ( .A(n_381), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_390), .A2(n_374), .B(n_367), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_380), .A2(n_392), .B(n_368), .Y(n_413) );
OA21x2_ASAP7_75t_L g414 ( .A1(n_365), .A2(n_381), .B(n_387), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_370), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_386), .Y(n_416) );
INVx4_ASAP7_75t_SL g417 ( .A(n_362), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_379), .B(n_333), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_389), .Y(n_419) );
NOR4xp25_ASAP7_75t_L g420 ( .A(n_384), .B(n_313), .C(n_359), .D(n_365), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_385), .A2(n_390), .B(n_383), .Y(n_421) );
OA21x2_ASAP7_75t_L g422 ( .A1(n_389), .A2(n_330), .B(n_393), .Y(n_422) );
HB1xp67_ASAP7_75t_SL g423 ( .A(n_407), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_420), .B(n_418), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_406), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_410), .Y(n_426) );
OAI21x1_ASAP7_75t_L g427 ( .A1(n_397), .A2(n_412), .B(n_421), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_414), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_414), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_417), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_410), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_417), .B(n_411), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_406), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_420), .B(n_418), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_396), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_419), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_419), .Y(n_437) );
INVxp67_ASAP7_75t_SL g438 ( .A(n_399), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_400), .A2(n_414), .B1(n_396), .B2(n_395), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_414), .B(n_404), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_404), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_394), .B(n_415), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_404), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_394), .B(n_415), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_410), .B(n_400), .Y(n_445) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_397), .A2(n_413), .B(n_419), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_416), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_416), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_405), .B(n_411), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_411), .B(n_410), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_422), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_408), .A2(n_403), .B1(n_405), .B2(n_401), .Y(n_452) );
BUFx3_ASAP7_75t_L g453 ( .A(n_403), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_422), .Y(n_454) );
NAND2x1p5_ASAP7_75t_L g455 ( .A(n_422), .B(n_417), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_411), .Y(n_456) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_405), .A2(n_398), .B(n_411), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_422), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_440), .B(n_443), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_441), .Y(n_460) );
INVx3_ASAP7_75t_L g461 ( .A(n_432), .Y(n_461) );
INVx4_ASAP7_75t_L g462 ( .A(n_453), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_440), .B(n_443), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_424), .B(n_417), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_441), .Y(n_465) );
NOR2x1_ASAP7_75t_SL g466 ( .A(n_453), .B(n_417), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_440), .B(n_403), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_447), .B(n_402), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_424), .B(n_409), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_432), .B(n_456), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_423), .A2(n_438), .B1(n_434), .B2(n_445), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_447), .B(n_448), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_434), .B(n_445), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_425), .B(n_433), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_448), .B(n_428), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_428), .B(n_429), .Y(n_476) );
OAI221xp5_ASAP7_75t_L g477 ( .A1(n_438), .A2(n_439), .B1(n_452), .B2(n_444), .C(n_442), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_423), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_453), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g480 ( .A(n_450), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_425), .B(n_433), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_429), .B(n_439), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_435), .Y(n_483) );
INVx1_ASAP7_75t_SL g484 ( .A(n_426), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_435), .B(n_450), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_427), .A2(n_452), .B(n_444), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_450), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_432), .B(n_456), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_451), .B(n_458), .Y(n_489) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_427), .A2(n_449), .B(n_458), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_436), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_442), .B(n_426), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_436), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_437), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_426), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_437), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_426), .B(n_431), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_451), .B(n_458), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_431), .B(n_454), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_451), .B(n_454), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_427), .A2(n_454), .B(n_449), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_446), .Y(n_502) );
INVx2_ASAP7_75t_SL g503 ( .A(n_432), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_432), .B(n_446), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_446), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_446), .B(n_457), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_446), .B(n_457), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_459), .B(n_457), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_474), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_459), .B(n_431), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_459), .B(n_431), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_489), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_478), .B(n_430), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_470), .B(n_430), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_463), .B(n_457), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_460), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_473), .B(n_463), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_460), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_463), .B(n_455), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_474), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_489), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_485), .B(n_455), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_485), .B(n_455), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_472), .B(n_455), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_472), .B(n_475), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_470), .B(n_488), .Y(n_526) );
INVx3_ASAP7_75t_L g527 ( .A(n_462), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_470), .B(n_488), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_465), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_499), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_480), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_473), .B(n_480), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_472), .B(n_475), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_479), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_479), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_469), .A2(n_471), .B1(n_477), .B2(n_467), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_475), .B(n_482), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_465), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_489), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_470), .B(n_488), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_476), .B(n_492), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_470), .B(n_488), .Y(n_542) );
OA21x2_ASAP7_75t_L g543 ( .A1(n_501), .A2(n_486), .B(n_505), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_499), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_467), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_498), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_483), .B(n_481), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_482), .B(n_476), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_483), .B(n_481), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_491), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_479), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_482), .B(n_476), .Y(n_552) );
INVxp67_ASAP7_75t_SL g553 ( .A(n_491), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_467), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_469), .A2(n_471), .B1(n_477), .B2(n_487), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_492), .B(n_468), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_498), .B(n_500), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_487), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_468), .B(n_500), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_496), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_496), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_468), .B(n_500), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_498), .Y(n_563) );
NOR2xp67_ASAP7_75t_L g564 ( .A(n_462), .B(n_461), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_488), .B(n_503), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_462), .B(n_487), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_557), .B(n_504), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_512), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_557), .B(n_504), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_509), .B(n_464), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_508), .B(n_504), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_520), .B(n_464), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_516), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_525), .B(n_462), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_525), .B(n_507), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_517), .B(n_503), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_508), .B(n_507), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_516), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_512), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_521), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g581 ( .A1(n_555), .A2(n_486), .B(n_497), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_518), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_533), .B(n_507), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_518), .Y(n_584) );
AND2x4_ASAP7_75t_L g585 ( .A(n_526), .B(n_503), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_529), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_515), .B(n_506), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_529), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_538), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_538), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_521), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_551), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_517), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_541), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_559), .B(n_502), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_562), .B(n_502), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_533), .B(n_506), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_541), .B(n_461), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_553), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_530), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_537), .B(n_506), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_548), .B(n_461), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_548), .B(n_461), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_552), .B(n_494), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_550), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_515), .B(n_501), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_552), .B(n_493), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_539), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_539), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_537), .B(n_490), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_546), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_556), .B(n_493), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_531), .B(n_495), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_544), .B(n_493), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_551), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_546), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_550), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_563), .B(n_494), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_519), .B(n_490), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_519), .B(n_524), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g621 ( .A1(n_581), .A2(n_536), .B(n_564), .Y(n_621) );
NAND2x1p5_ASAP7_75t_L g622 ( .A(n_592), .B(n_527), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_600), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_606), .B(n_561), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_594), .Y(n_625) );
NAND2x1_ASAP7_75t_L g626 ( .A(n_585), .B(n_527), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_567), .B(n_528), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_575), .B(n_554), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_584), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_567), .B(n_526), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_584), .Y(n_631) );
NOR2xp33_ASAP7_75t_SL g632 ( .A(n_615), .B(n_535), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_593), .B(n_532), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_569), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_569), .B(n_540), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_586), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_620), .B(n_531), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_576), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_586), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_583), .B(n_532), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_577), .B(n_549), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_605), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_605), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_620), .B(n_540), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_617), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_614), .Y(n_646) );
OR2x6_ASAP7_75t_L g647 ( .A(n_585), .B(n_527), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_597), .B(n_511), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_606), .B(n_561), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_571), .B(n_540), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_617), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_576), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_613), .A2(n_566), .B(n_513), .C(n_558), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_601), .B(n_595), .Y(n_654) );
INVx2_ASAP7_75t_SL g655 ( .A(n_585), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_573), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_610), .B(n_547), .Y(n_657) );
INVxp67_ASAP7_75t_L g658 ( .A(n_595), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_621), .A2(n_574), .B(n_599), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_629), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_646), .Y(n_661) );
AOI21xp33_ASAP7_75t_L g662 ( .A1(n_621), .A2(n_543), .B(n_572), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_658), .A2(n_619), .B1(n_610), .B2(n_542), .Y(n_663) );
O2A1O1Ixp33_ASAP7_75t_L g664 ( .A1(n_623), .A2(n_570), .B(n_598), .C(n_596), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_632), .A2(n_534), .B(n_571), .Y(n_665) );
BUFx2_ASAP7_75t_L g666 ( .A(n_647), .Y(n_666) );
INVxp67_ASAP7_75t_SL g667 ( .A(n_622), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_631), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_646), .B(n_577), .Y(n_669) );
AOI21xp33_ASAP7_75t_L g670 ( .A1(n_632), .A2(n_543), .B(n_578), .Y(n_670) );
OAI32xp33_ASAP7_75t_L g671 ( .A1(n_622), .A2(n_598), .A3(n_603), .B1(n_602), .B2(n_596), .Y(n_671) );
AOI21xp33_ASAP7_75t_L g672 ( .A1(n_626), .A2(n_543), .B(n_582), .Y(n_672) );
INVx1_ASAP7_75t_SL g673 ( .A(n_644), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_636), .Y(n_674) );
OAI21xp5_ASAP7_75t_SL g675 ( .A1(n_653), .A2(n_542), .B(n_528), .Y(n_675) );
OAI31xp33_ASAP7_75t_L g676 ( .A1(n_637), .A2(n_619), .A3(n_565), .B(n_587), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_625), .A2(n_587), .B1(n_590), .B2(n_588), .C(n_589), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_634), .B(n_580), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_624), .B(n_568), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g680 ( .A1(n_633), .A2(n_603), .B(n_602), .C(n_612), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_639), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_642), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_675), .A2(n_652), .B1(n_655), .B2(n_638), .Y(n_683) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_676), .A2(n_647), .B1(n_624), .B2(n_649), .C(n_657), .Y(n_684) );
O2A1O1Ixp33_ASAP7_75t_L g685 ( .A1(n_662), .A2(n_649), .B(n_640), .C(n_657), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_661), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_671), .A2(n_641), .B1(n_656), .B2(n_651), .C(n_645), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_659), .A2(n_647), .B1(n_650), .B2(n_630), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_666), .A2(n_654), .B1(n_628), .B2(n_635), .Y(n_689) );
XOR2x2_ASAP7_75t_L g690 ( .A(n_665), .B(n_627), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_671), .A2(n_618), .B(n_466), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_663), .A2(n_666), .B1(n_677), .B2(n_667), .Y(n_692) );
OAI31xp33_ASAP7_75t_L g693 ( .A1(n_661), .A2(n_542), .A3(n_528), .B(n_526), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_664), .A2(n_466), .B(n_565), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_670), .A2(n_643), .B(n_648), .Y(n_695) );
OAI21x1_ASAP7_75t_SL g696 ( .A1(n_680), .A2(n_604), .B(n_607), .Y(n_696) );
OAI221xp5_ASAP7_75t_SL g697 ( .A1(n_693), .A2(n_673), .B1(n_669), .B2(n_679), .C(n_545), .Y(n_697) );
O2A1O1Ixp5_ASAP7_75t_SL g698 ( .A1(n_686), .A2(n_672), .B(n_660), .C(n_681), .Y(n_698) );
NAND3xp33_ASAP7_75t_SL g699 ( .A(n_687), .B(n_682), .C(n_674), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_685), .A2(n_668), .B1(n_678), .B2(n_616), .C(n_611), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_692), .A2(n_678), .B1(n_565), .B2(n_514), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_684), .A2(n_514), .B1(n_524), .B2(n_522), .Y(n_702) );
AOI321xp33_ASAP7_75t_L g703 ( .A1(n_683), .A2(n_514), .A3(n_522), .B1(n_510), .B2(n_523), .C(n_616), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_695), .A2(n_568), .B1(n_609), .B2(n_608), .C(n_591), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_699), .A2(n_696), .B1(n_689), .B2(n_691), .C(n_688), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_701), .Y(n_706) );
NAND4xp25_ASAP7_75t_L g707 ( .A(n_697), .B(n_694), .C(n_690), .D(n_495), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_698), .B(n_579), .C(n_609), .Y(n_708) );
INVxp67_ASAP7_75t_SL g709 ( .A(n_700), .Y(n_709) );
NOR3xp33_ASAP7_75t_L g710 ( .A(n_707), .B(n_704), .C(n_703), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_705), .B(n_702), .Y(n_711) );
AND4x1_ASAP7_75t_L g712 ( .A(n_708), .B(n_560), .C(n_607), .D(n_604), .Y(n_712) );
AND2x4_ASAP7_75t_L g713 ( .A(n_711), .B(n_706), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_710), .A2(n_709), .B(n_611), .Y(n_714) );
NAND3x1_ASAP7_75t_L g715 ( .A(n_714), .B(n_712), .C(n_495), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_715), .Y(n_716) );
NOR3xp33_ASAP7_75t_L g717 ( .A(n_716), .B(n_713), .C(n_608), .Y(n_717) );
OAI21xp5_ASAP7_75t_SL g718 ( .A1(n_717), .A2(n_591), .B(n_580), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_718), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_719), .A2(n_579), .B(n_484), .Y(n_720) );
endmodule