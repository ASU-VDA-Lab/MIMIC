module fake_jpeg_6899_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_38),
.B1(n_25),
.B2(n_20),
.Y(n_44)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_42),
.B(n_2),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_21),
.Y(n_43)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_46),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_52),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_20),
.B1(n_15),
.B2(n_37),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_32),
.A2(n_20),
.B1(n_25),
.B2(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_25),
.B1(n_15),
.B2(n_31),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_18),
.B1(n_31),
.B2(n_21),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_61),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_30),
.B(n_28),
.C(n_26),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_40),
.B(n_38),
.C(n_23),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_32),
.A2(n_30),
.B1(n_22),
.B2(n_28),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_26),
.B1(n_24),
.B2(n_22),
.Y(n_62)
);

AO22x1_ASAP7_75t_SL g68 ( 
.A1(n_62),
.A2(n_19),
.B1(n_29),
.B2(n_16),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_69),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_57),
.B1(n_32),
.B2(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_72),
.Y(n_83)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_60),
.Y(n_93)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_81),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_80),
.A2(n_58),
.B1(n_57),
.B2(n_47),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_67),
.B1(n_55),
.B2(n_79),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_98),
.B1(n_77),
.B2(n_74),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_48),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_87),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_99),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_70),
.B(n_76),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_96),
.B(n_83),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_57),
.B1(n_41),
.B2(n_34),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_39),
.C(n_40),
.Y(n_99)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_105),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_110),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_69),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_65),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_122),
.B1(n_100),
.B2(n_73),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_116),
.A2(n_23),
.B(n_19),
.Y(n_143)
);

AOI22x1_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_64),
.B1(n_48),
.B2(n_40),
.Y(n_117)
);

OAI22x1_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_39),
.B1(n_41),
.B2(n_34),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_59),
.B(n_74),
.Y(n_120)
);

OA21x2_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_73),
.B(n_92),
.Y(n_142)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_91),
.B(n_86),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_127),
.B(n_107),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_92),
.B(n_100),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_131),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_141),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_101),
.C(n_95),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_138),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_97),
.C(n_39),
.Y(n_138)
);

AOI221xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_120),
.B1(n_116),
.B2(n_111),
.C(n_113),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_105),
.B1(n_117),
.B2(n_119),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_142),
.B1(n_144),
.B2(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_104),
.B(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_149),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_153),
.B(n_106),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_155),
.Y(n_164)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_161),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_120),
.B1(n_115),
.B2(n_124),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_163),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_136),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_133),
.C(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_125),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_115),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_144),
.Y(n_172)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_SL g165 ( 
.A(n_153),
.B(n_126),
.C(n_143),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_178),
.Y(n_189)
);

XNOR2x1_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_131),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_172),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_169),
.C(n_174),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_134),
.C(n_135),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_137),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_171),
.B(n_176),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g173 ( 
.A(n_161),
.Y(n_173)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_128),
.C(n_142),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_162),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_13),
.C(n_41),
.Y(n_178)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_175),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_160),
.C(n_150),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_190),
.C(n_41),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_2),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_188),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_167),
.B(n_163),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_174),
.C(n_166),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_179),
.A2(n_123),
.B1(n_50),
.B2(n_19),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_191),
.B(n_192),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_19),
.B1(n_29),
.B2(n_16),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_190),
.A2(n_177),
.B(n_165),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_3),
.B(n_7),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_195),
.B(n_200),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_178),
.B(n_59),
.C(n_50),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_201),
.B(n_34),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_7),
.C(n_8),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_184),
.B(n_3),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_29),
.B(n_34),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_189),
.B1(n_185),
.B2(n_181),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_206),
.Y(n_211)
);

AOI31xp33_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_181),
.A3(n_29),
.B(n_6),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_204),
.A2(n_205),
.B(n_207),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_197),
.A2(n_12),
.B1(n_4),
.B2(n_6),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_194),
.B(n_3),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_210),
.C(n_201),
.Y(n_214)
);

OAI221xp5_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_198),
.B1(n_195),
.B2(n_199),
.C(n_202),
.Y(n_212)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_215),
.C(n_216),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_9),
.B(n_10),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_9),
.B(n_10),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_206),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_219),
.A2(n_220),
.B(n_11),
.Y(n_222)
);

AOI21x1_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_203),
.B(n_10),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_9),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_218),
.B(n_12),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_223),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_11),
.B(n_12),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_224),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_225),
.Y(n_227)
);


endmodule