module fake_jpeg_29123_n_104 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_3),
.B(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_17),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_33),
.B1(n_36),
.B2(n_44),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_62),
.B1(n_48),
.B2(n_52),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_4),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_63),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_43),
.B(n_52),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_23),
.C(n_24),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_69),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_4),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_73),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_75),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_5),
.Y(n_75)
);

AOI32xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_19),
.A3(n_31),
.B1(n_7),
.B2(n_8),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_88),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_82),
.B1(n_29),
.B2(n_32),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_18),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_27),
.C(n_28),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_86),
.A2(n_88),
.B(n_85),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_89),
.B(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

AOI22x1_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_85),
.B1(n_87),
.B2(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_95),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_98),
.B(n_93),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_94),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_100),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_97),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_78),
.B(n_96),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_89),
.Y(n_104)
);


endmodule