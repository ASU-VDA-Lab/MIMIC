module fake_jpeg_17887_n_166 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_166);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

INVx8_ASAP7_75t_SL g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_0),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_55),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_68),
.Y(n_71)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_45),
.B1(n_60),
.B2(n_41),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_80),
.B1(n_53),
.B2(n_44),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_59),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_79),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_56),
.B1(n_47),
.B2(n_54),
.Y(n_80)
);

INVx5_ASAP7_75t_SL g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

CKINVDCx6p67_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_47),
.B1(n_52),
.B2(n_51),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_106),
.B1(n_109),
.B2(n_8),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_94),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_71),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_79),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_110),
.C(n_7),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_0),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_1),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_2),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_107),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_42),
.B1(n_53),
.B2(n_40),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_3),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_6),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_29),
.B1(n_38),
.B2(n_37),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_3),
.B(n_4),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_6),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_89),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_118),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_119),
.A2(n_103),
.B(n_89),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_129),
.Y(n_134)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_125),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_133),
.B(n_128),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_132),
.A2(n_125),
.B1(n_114),
.B2(n_120),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_136),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_127),
.B(n_117),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_137),
.A2(n_124),
.B(n_119),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_139),
.B(n_141),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_140),
.B(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_98),
.B1(n_96),
.B2(n_107),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_147),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_97),
.C(n_95),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_138),
.C(n_130),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_151),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_146),
.C(n_12),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_149),
.A2(n_145),
.B1(n_132),
.B2(n_112),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_153),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_11),
.C(n_15),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_18),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_39),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_20),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_22),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_23),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_24),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_26),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_28),
.C(n_30),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_31),
.Y(n_166)
);


endmodule