module fake_jpeg_24875_n_37 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_37);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NAND3xp33_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_0),
.C(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_12),
.B(n_4),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_12),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_17),
.A2(n_22),
.B(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_19),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_16),
.C(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_32),
.B(n_24),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_18),
.B(n_30),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_34),
.C(n_32),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_30),
.B(n_23),
.Y(n_37)
);


endmodule