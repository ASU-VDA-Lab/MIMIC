module fake_ariane_1596_n_1725 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1725);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1725;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_153),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_55),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_65),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_66),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_31),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_3),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_107),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_23),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_18),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_128),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_120),
.Y(n_175)
);

BUFx8_ASAP7_75t_SL g176 ( 
.A(n_93),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_11),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_68),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_76),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_96),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_18),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_97),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_72),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_6),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_40),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_79),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_81),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_31),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_48),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_89),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_143),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_29),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_57),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_91),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_25),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_17),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_32),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_67),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_25),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_124),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_155),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_43),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_99),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_73),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_149),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_58),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_11),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_46),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_34),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_112),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_104),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_122),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_43),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_74),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_5),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_105),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_88),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_34),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_60),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_21),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_52),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_134),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_129),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_111),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_119),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_37),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_98),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_29),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_114),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_82),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_100),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_20),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_59),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_48),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_44),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_152),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_141),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_55),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_8),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_37),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_108),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_84),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_109),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_136),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_130),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_61),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_6),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_62),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_32),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_28),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_27),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_101),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_158),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_142),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_75),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_85),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_54),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_28),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_110),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_95),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_2),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_148),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_16),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_20),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_53),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_103),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_10),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_24),
.Y(n_273)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_19),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_80),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_137),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_106),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_10),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_14),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_42),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_132),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_21),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_83),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_154),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_53),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_50),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_19),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_144),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_77),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_14),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_23),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_24),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_113),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_87),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_35),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_70),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_116),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_159),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_147),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_8),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_64),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_71),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_78),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_42),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_133),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_69),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_2),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_63),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_45),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_39),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_102),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_15),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_13),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_146),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_176),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_209),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_200),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_184),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_200),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_178),
.B(n_1),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_200),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_173),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_204),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_200),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_200),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_166),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_200),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_166),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_276),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_175),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_200),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_223),
.B(n_4),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_263),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_175),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_266),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_212),
.B(n_5),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_312),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_310),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_263),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_R g340 ( 
.A(n_187),
.B(n_121),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_263),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_263),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_162),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_187),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_194),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_263),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_169),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_263),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_223),
.B(n_7),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_268),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_194),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_218),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_268),
.B(n_7),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_263),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_170),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_184),
.B(n_9),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_274),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_188),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_189),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_272),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_192),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_197),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_196),
.B(n_9),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_274),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_227),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_227),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_198),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_203),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_274),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_274),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_210),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_274),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_218),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_289),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_304),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_274),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_289),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_221),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_274),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_196),
.B(n_234),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_272),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_311),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_234),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_224),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_314),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_164),
.B(n_12),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_311),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_314),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_272),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_237),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_272),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_243),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_272),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_172),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_193),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_172),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_304),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_230),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_193),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_230),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_244),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_252),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_240),
.Y(n_403)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_317),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_342),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_342),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_317),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_319),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_240),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_323),
.B(n_262),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_385),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_385),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_388),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_398),
.B(n_262),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_319),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_321),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_321),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_400),
.B(n_276),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_324),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_324),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_383),
.B(n_276),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_325),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_337),
.A2(n_291),
.B1(n_280),
.B2(n_245),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_316),
.B(n_292),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_L g431 ( 
.A(n_340),
.B(n_314),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_360),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_393),
.B(n_165),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_325),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_329),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g436 ( 
.A(n_327),
.B(n_257),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_327),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_331),
.B(n_167),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_331),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_333),
.B(n_183),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_333),
.A2(n_251),
.B(n_220),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_323),
.B(n_191),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_339),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_339),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_341),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_341),
.B(n_195),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_346),
.B(n_199),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_360),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_323),
.B(n_318),
.Y(n_449)
);

OA21x2_ASAP7_75t_L g450 ( 
.A1(n_381),
.A2(n_251),
.B(n_220),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_383),
.B(n_191),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_395),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_391),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_346),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_320),
.B(n_332),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_348),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_348),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_380),
.B(n_204),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_332),
.B(n_201),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_354),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_354),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_357),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_357),
.B(n_205),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_364),
.B(n_206),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_364),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_369),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_369),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_353),
.B(n_201),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_375),
.B(n_219),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_353),
.B(n_208),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_370),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_370),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_372),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_372),
.B(n_208),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_376),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_376),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_379),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_379),
.B(n_303),
.Y(n_478)
);

INVxp33_ASAP7_75t_SL g479 ( 
.A(n_315),
.Y(n_479)
);

OA21x2_ASAP7_75t_L g480 ( 
.A1(n_381),
.A2(n_217),
.B(n_207),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_389),
.Y(n_481)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_406),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_458),
.B(n_350),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_413),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_421),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_413),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_413),
.Y(n_487)
);

OAI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_430),
.A2(n_336),
.B1(n_349),
.B2(n_386),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_469),
.B(n_347),
.C(n_343),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_469),
.B(n_316),
.Y(n_490)
);

INVxp33_ASAP7_75t_L g491 ( 
.A(n_406),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_421),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_427),
.B(n_355),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_449),
.B(n_358),
.Y(n_494)
);

CKINVDCx6p67_ASAP7_75t_R g495 ( 
.A(n_452),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_413),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_427),
.B(n_352),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_427),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_421),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_415),
.Y(n_500)
);

OAI22xp33_ASAP7_75t_L g501 ( 
.A1(n_430),
.A2(n_245),
.B1(n_280),
.B2(n_273),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_415),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_451),
.B(n_359),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_428),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_451),
.B(n_361),
.Y(n_505)
);

INVxp33_ASAP7_75t_L g506 ( 
.A(n_429),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_431),
.A2(n_291),
.B1(n_273),
.B2(n_356),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_421),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_426),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_426),
.Y(n_510)
);

BUFx6f_ASAP7_75t_SL g511 ( 
.A(n_451),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_428),
.Y(n_512)
);

NAND3xp33_ASAP7_75t_L g513 ( 
.A(n_431),
.B(n_367),
.C(n_362),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_426),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_449),
.B(n_459),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_452),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_415),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_428),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_415),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_458),
.B(n_394),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_459),
.B(n_368),
.Y(n_521)
);

INVx4_ASAP7_75t_SL g522 ( 
.A(n_436),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_414),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_419),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_419),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_L g526 ( 
.A(n_428),
.B(n_314),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_459),
.B(n_468),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_419),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_426),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_445),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_459),
.B(n_371),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_428),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_419),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_445),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_445),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_414),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_424),
.B(n_373),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_420),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_459),
.B(n_378),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_R g540 ( 
.A(n_435),
.B(n_322),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_420),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_445),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_468),
.B(n_470),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_428),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_435),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_454),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_451),
.B(n_384),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_428),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_468),
.B(n_390),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_424),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_468),
.A2(n_363),
.B1(n_397),
.B2(n_177),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_414),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_420),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_405),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_420),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_408),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_408),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_441),
.A2(n_238),
.B(n_226),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_405),
.B(n_401),
.C(n_392),
.Y(n_559)
);

OAI21xp33_ASAP7_75t_SL g560 ( 
.A1(n_455),
.A2(n_441),
.B(n_418),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_429),
.B(n_338),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_408),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_451),
.B(n_402),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_468),
.B(n_389),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_443),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_455),
.B(n_225),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_408),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_470),
.A2(n_232),
.B1(n_256),
.B2(n_307),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_SL g569 ( 
.A(n_470),
.B(n_309),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_436),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_454),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_470),
.B(n_442),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_454),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_454),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_411),
.B(n_394),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_458),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_433),
.B(n_470),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_407),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_414),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_443),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_442),
.B(n_391),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_407),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_409),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_412),
.B(n_403),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_409),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_474),
.A2(n_309),
.B1(n_313),
.B2(n_254),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_443),
.Y(n_587)
);

OR2x6_ASAP7_75t_L g588 ( 
.A(n_412),
.B(n_403),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_R g589 ( 
.A(n_479),
.B(n_326),
.Y(n_589)
);

INVxp33_ASAP7_75t_L g590 ( 
.A(n_411),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_412),
.A2(n_216),
.B1(n_295),
.B2(n_279),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_410),
.Y(n_592)
);

OAI22xp33_ASAP7_75t_L g593 ( 
.A1(n_479),
.A2(n_286),
.B1(n_313),
.B2(n_278),
.Y(n_593)
);

AOI22x1_ASAP7_75t_L g594 ( 
.A1(n_457),
.A2(n_287),
.B1(n_269),
.B2(n_270),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_407),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_442),
.B(n_160),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_407),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_443),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_442),
.B(n_303),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_412),
.B(n_181),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_410),
.Y(n_601)
);

INVx5_ASAP7_75t_L g602 ( 
.A(n_436),
.Y(n_602)
);

INVxp33_ASAP7_75t_L g603 ( 
.A(n_411),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_407),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_414),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_414),
.Y(n_606)
);

NOR2x1p5_ASAP7_75t_L g607 ( 
.A(n_418),
.B(n_255),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_442),
.A2(n_478),
.B1(n_480),
.B2(n_474),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_474),
.B(n_228),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_422),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_443),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_478),
.A2(n_185),
.B1(n_285),
.B2(n_300),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_422),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_423),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_414),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_423),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_418),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_478),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_478),
.A2(n_290),
.B1(n_211),
.B2(n_239),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_443),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_478),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_425),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_416),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_474),
.B(n_247),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_425),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_434),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_474),
.B(n_257),
.Y(n_627)
);

BUFx10_ASAP7_75t_L g628 ( 
.A(n_434),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_437),
.B(n_298),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_433),
.B(n_242),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_416),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_577),
.B(n_457),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_556),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_556),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_557),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_494),
.B(n_330),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_506),
.A2(n_344),
.B1(n_345),
.B2(n_334),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_550),
.A2(n_480),
.B1(n_450),
.B2(n_440),
.Y(n_638)
);

AND2x4_ASAP7_75t_SL g639 ( 
.A(n_497),
.B(n_351),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_554),
.Y(n_640)
);

BUFx6f_ASAP7_75t_SL g641 ( 
.A(n_483),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_628),
.B(n_457),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_583),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_550),
.B(n_457),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_628),
.B(n_457),
.Y(n_645)
);

BUFx6f_ASAP7_75t_SL g646 ( 
.A(n_483),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_557),
.Y(n_647)
);

BUFx6f_ASAP7_75t_SL g648 ( 
.A(n_483),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_589),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_515),
.B(n_461),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_628),
.B(n_488),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_566),
.B(n_461),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_488),
.B(n_461),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_537),
.B(n_365),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_490),
.B(n_366),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_536),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_630),
.B(n_461),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_617),
.B(n_461),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_498),
.A2(n_439),
.B1(n_437),
.B2(n_444),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_618),
.B(n_462),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_617),
.B(n_462),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_527),
.B(n_462),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_618),
.B(n_462),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_498),
.A2(n_465),
.B1(n_439),
.B2(n_456),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_543),
.B(n_462),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_629),
.B(n_471),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_516),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_562),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_572),
.B(n_471),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_609),
.B(n_471),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_537),
.B(n_374),
.Y(n_671)
);

NOR2xp67_ASAP7_75t_SL g672 ( 
.A(n_489),
.B(n_513),
.Y(n_672)
);

AND2x2_ASAP7_75t_SL g673 ( 
.A(n_507),
.B(n_480),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_624),
.B(n_520),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_497),
.B(n_377),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_536),
.B(n_471),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_562),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_482),
.B(n_382),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_536),
.B(n_471),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_607),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_491),
.B(n_387),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_507),
.A2(n_551),
.B1(n_511),
.B2(n_608),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_567),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_520),
.B(n_575),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_567),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_520),
.B(n_477),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_484),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_575),
.B(n_477),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_522),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_536),
.B(n_477),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_576),
.B(n_477),
.Y(n_691)
);

O2A1O1Ixp5_ASAP7_75t_L g692 ( 
.A1(n_523),
.A2(n_565),
.B(n_512),
.C(n_596),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_L g693 ( 
.A(n_559),
.B(n_453),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_484),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_585),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_592),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_621),
.B(n_477),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_545),
.B(n_399),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_621),
.B(n_444),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_607),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_590),
.B(n_292),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_552),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_516),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_L g704 ( 
.A(n_552),
.B(n_443),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_486),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_486),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_495),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_487),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_603),
.B(n_456),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_495),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_552),
.B(n_460),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_592),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_601),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_601),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_561),
.B(n_292),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_610),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_487),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_561),
.B(n_438),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_610),
.B(n_460),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_588),
.B(n_441),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_521),
.A2(n_472),
.B1(n_476),
.B2(n_475),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_493),
.B(n_465),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_579),
.B(n_466),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_613),
.B(n_466),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_579),
.B(n_467),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_613),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_511),
.A2(n_569),
.B1(n_539),
.B2(n_549),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_614),
.B(n_467),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_531),
.A2(n_476),
.B1(n_475),
.B2(n_473),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_579),
.B(n_472),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_540),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_579),
.B(n_443),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_511),
.A2(n_440),
.B1(n_446),
.B2(n_464),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_616),
.B(n_446),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_594),
.B(n_447),
.C(n_464),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_588),
.B(n_447),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_503),
.B(n_463),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_568),
.B(n_463),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_574),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_496),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_599),
.A2(n_547),
.B1(n_563),
.B2(n_505),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_599),
.A2(n_160),
.B1(n_174),
.B2(n_179),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_599),
.A2(n_480),
.B1(n_450),
.B2(n_453),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_622),
.B(n_416),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_605),
.B(n_414),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_568),
.B(n_282),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_593),
.B(n_417),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_622),
.B(n_416),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_599),
.A2(n_480),
.B1(n_450),
.B2(n_453),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_496),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_625),
.B(n_416),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_625),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_605),
.B(n_417),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_626),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_605),
.B(n_417),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_600),
.B(n_417),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_626),
.B(n_432),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_605),
.B(n_417),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_600),
.B(n_588),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_600),
.B(n_417),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_594),
.B(n_586),
.C(n_612),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_584),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_599),
.B(n_432),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_606),
.B(n_417),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_600),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_599),
.A2(n_480),
.B1(n_450),
.B2(n_453),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_599),
.B(n_432),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_588),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_581),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_606),
.B(n_448),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_512),
.B(n_174),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_564),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_500),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_500),
.Y(n_774)
);

NOR2xp67_ASAP7_75t_L g775 ( 
.A(n_623),
.B(n_453),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_502),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_578),
.B(n_448),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_574),
.Y(n_778)
);

INVx8_ASAP7_75t_L g779 ( 
.A(n_627),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_502),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_517),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_517),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_578),
.Y(n_783)
);

NOR3xp33_ASAP7_75t_L g784 ( 
.A(n_560),
.B(n_565),
.C(n_512),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_519),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_606),
.B(n_448),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_619),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_519),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_485),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_636),
.B(n_623),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_632),
.A2(n_565),
.B(n_504),
.Y(n_791)
);

A2O1A1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_737),
.A2(n_631),
.B(n_535),
.C(n_534),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_643),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_761),
.A2(n_631),
.B(n_535),
.C(n_534),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_689),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_736),
.A2(n_627),
.B1(n_485),
.B2(n_492),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_718),
.B(n_591),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_639),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_735),
.A2(n_650),
.B(n_662),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_657),
.A2(n_532),
.B(n_518),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_674),
.B(n_492),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_738),
.B(n_499),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_739),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_695),
.Y(n_804)
);

BUFx6f_ASAP7_75t_SL g805 ( 
.A(n_680),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_734),
.A2(n_548),
.B(n_544),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_652),
.A2(n_548),
.B(n_544),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_673),
.A2(n_627),
.B1(n_571),
.B2(n_529),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_736),
.B(n_508),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_666),
.A2(n_580),
.B(n_548),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_653),
.A2(n_546),
.B(n_509),
.C(n_510),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_736),
.B(n_508),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_696),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_L g814 ( 
.A(n_702),
.B(n_784),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_665),
.A2(n_510),
.B(n_509),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_709),
.B(n_514),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_712),
.A2(n_542),
.B1(n_529),
.B2(n_530),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_722),
.B(n_514),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_768),
.B(n_606),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_691),
.B(n_530),
.Y(n_820)
);

INVxp67_ASAP7_75t_SL g821 ( 
.A(n_720),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_699),
.B(n_542),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_SL g823 ( 
.A(n_731),
.B(n_627),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_688),
.B(n_546),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_772),
.B(n_571),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_739),
.Y(n_826)
);

CKINVDCx10_ASAP7_75t_R g827 ( 
.A(n_641),
.Y(n_827)
);

AO21x1_ASAP7_75t_L g828 ( 
.A1(n_653),
.A2(n_573),
.B(n_526),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_669),
.A2(n_573),
.B(n_525),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_745),
.A2(n_598),
.B(n_587),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_747),
.A2(n_595),
.B(n_582),
.C(n_597),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_713),
.A2(n_595),
.B(n_582),
.C(n_597),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_715),
.B(n_587),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_714),
.A2(n_598),
.B1(n_620),
.B2(n_611),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_719),
.A2(n_604),
.B(n_481),
.C(n_448),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_762),
.B(n_604),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_651),
.B(n_703),
.C(n_667),
.Y(n_837)
);

CKINVDCx10_ASAP7_75t_R g838 ( 
.A(n_641),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_739),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_741),
.B(n_615),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_753),
.A2(n_615),
.B(n_528),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_676),
.A2(n_524),
.B(n_525),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_716),
.A2(n_615),
.B1(n_524),
.B2(n_528),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_755),
.A2(n_615),
.B(n_533),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_724),
.A2(n_526),
.B(n_533),
.C(n_555),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_639),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_682),
.B(n_538),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_689),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_676),
.A2(n_541),
.B(n_553),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_759),
.Y(n_850)
);

NAND2x1_ASAP7_75t_L g851 ( 
.A(n_689),
.B(n_541),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_654),
.B(n_553),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_755),
.A2(n_615),
.B(n_555),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_733),
.B(n_627),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_779),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_759),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_758),
.A2(n_558),
.B(n_450),
.Y(n_857)
);

AO21x1_ASAP7_75t_L g858 ( 
.A1(n_651),
.A2(n_253),
.B(n_248),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_758),
.A2(n_558),
.B(n_450),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_728),
.A2(n_284),
.B(n_261),
.C(n_299),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_726),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_710),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_671),
.B(n_558),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_778),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_769),
.B(n_627),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_675),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_752),
.B(n_754),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_759),
.A2(n_648),
.B1(n_646),
.B2(n_673),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_701),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_686),
.B(n_640),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_764),
.A2(n_570),
.B(n_602),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_759),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_787),
.B(n_697),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_727),
.B(n_179),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_659),
.B(n_664),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_679),
.A2(n_627),
.B(n_436),
.Y(n_876)
);

OAI21xp33_ASAP7_75t_L g877 ( 
.A1(n_644),
.A2(n_186),
.B(n_308),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_778),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_649),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_702),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_658),
.B(n_180),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_720),
.B(n_522),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_661),
.B(n_180),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_670),
.B(n_182),
.Y(n_884)
);

OAI21xp33_ASAP7_75t_SL g885 ( 
.A1(n_642),
.A2(n_645),
.B(n_660),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_756),
.A2(n_294),
.B(n_182),
.C(n_308),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_721),
.A2(n_12),
.B(n_13),
.C(n_16),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_778),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_679),
.A2(n_602),
.B(n_570),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_765),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_646),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_742),
.B(n_186),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_690),
.A2(n_436),
.B(n_570),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_690),
.A2(n_732),
.B(n_723),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_789),
.A2(n_306),
.B1(n_305),
.B2(n_602),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_789),
.B(n_305),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_720),
.B(n_306),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_760),
.A2(n_602),
.B(n_570),
.C(n_190),
.Y(n_898)
);

INVx11_ASAP7_75t_L g899 ( 
.A(n_648),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_678),
.Y(n_900)
);

O2A1O1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_729),
.A2(n_17),
.B(n_22),
.C(n_26),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_771),
.B(n_522),
.Y(n_902)
);

NOR2xp67_ASAP7_75t_L g903 ( 
.A(n_681),
.B(n_602),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_779),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_779),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_732),
.A2(n_602),
.B(n_570),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_700),
.B(n_570),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_707),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_711),
.A2(n_436),
.B(n_404),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_725),
.A2(n_168),
.B(n_171),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_744),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_702),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_779),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_730),
.A2(n_163),
.B(n_161),
.Y(n_914)
);

INVx11_ASAP7_75t_L g915 ( 
.A(n_698),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_730),
.A2(n_202),
.B(n_213),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_783),
.Y(n_917)
);

AO21x1_ASAP7_75t_L g918 ( 
.A1(n_660),
.A2(n_314),
.B(n_288),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_704),
.A2(n_264),
.B(n_215),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_663),
.A2(n_260),
.B(n_222),
.C(n_302),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_663),
.B(n_672),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_655),
.B(n_22),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_748),
.A2(n_751),
.B(n_757),
.C(n_692),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_704),
.A2(n_265),
.B(n_229),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_770),
.A2(n_267),
.B(n_231),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_746),
.B(n_788),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_687),
.B(n_259),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_R g928 ( 
.A(n_763),
.B(n_235),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_786),
.A2(n_275),
.B(n_233),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_694),
.B(n_271),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_656),
.B(n_404),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_702),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_777),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_637),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_705),
.A2(n_277),
.B(n_236),
.C(n_301),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_706),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_706),
.B(n_258),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_775),
.A2(n_788),
.B(n_785),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_708),
.A2(n_283),
.B(n_241),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_656),
.B(n_404),
.Y(n_940)
);

INVx6_ASAP7_75t_L g941 ( 
.A(n_656),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_693),
.A2(n_214),
.B1(n_246),
.B2(n_249),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_638),
.A2(n_436),
.B(n_404),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_708),
.A2(n_785),
.B(n_782),
.C(n_781),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_717),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_767),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_717),
.B(n_297),
.Y(n_947)
);

NOR2x2_ASAP7_75t_L g948 ( 
.A(n_740),
.B(n_26),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_750),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_750),
.A2(n_436),
.B1(n_257),
.B2(n_288),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_773),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_774),
.A2(n_782),
.B(n_781),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_SL g953 ( 
.A1(n_774),
.A2(n_27),
.B(n_30),
.C(n_33),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_922),
.A2(n_780),
.B(n_776),
.C(n_634),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_922),
.A2(n_780),
.B(n_776),
.C(n_634),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_SL g956 ( 
.A(n_887),
.B(n_901),
.C(n_885),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_821),
.A2(n_633),
.B(n_635),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_821),
.A2(n_766),
.B1(n_749),
.B2(n_743),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_790),
.A2(n_685),
.B(n_683),
.C(n_677),
.Y(n_959)
);

INVx3_ASAP7_75t_SL g960 ( 
.A(n_948),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_873),
.B(n_685),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_818),
.A2(n_683),
.B(n_677),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_790),
.A2(n_833),
.B(n_875),
.C(n_860),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_867),
.A2(n_668),
.B1(n_647),
.B2(n_293),
.Y(n_964)
);

AND2x2_ASAP7_75t_SL g965 ( 
.A(n_808),
.B(n_288),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_926),
.B(n_668),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_814),
.A2(n_647),
.B(n_250),
.Y(n_967)
);

OAI22x1_ASAP7_75t_L g968 ( 
.A1(n_934),
.A2(n_281),
.B1(n_296),
.B2(n_36),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_850),
.B(n_404),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_900),
.B(n_38),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_899),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_902),
.A2(n_288),
.B(n_257),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_795),
.Y(n_973)
);

O2A1O1Ixp5_ASAP7_75t_L g974 ( 
.A1(n_799),
.A2(n_314),
.B(n_436),
.C(n_41),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_802),
.A2(n_404),
.B1(n_288),
.B2(n_41),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_791),
.A2(n_404),
.B(n_436),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_890),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_824),
.A2(n_404),
.B(n_94),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_921),
.B(n_880),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_797),
.B(n_38),
.Y(n_980)
);

BUFx12f_ASAP7_75t_L g981 ( 
.A(n_798),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_846),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_852),
.B(n_39),
.Y(n_983)
);

NAND3xp33_ASAP7_75t_SL g984 ( 
.A(n_887),
.B(n_44),
.C(n_45),
.Y(n_984)
);

AO22x1_ASAP7_75t_L g985 ( 
.A1(n_891),
.A2(n_404),
.B1(n_47),
.B2(n_49),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_833),
.A2(n_314),
.B(n_47),
.C(n_49),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_917),
.B(n_46),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_793),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_SL g989 ( 
.A1(n_868),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_837),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_917),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_800),
.A2(n_125),
.B(n_150),
.Y(n_992)
);

AOI21x1_ASAP7_75t_L g993 ( 
.A1(n_857),
.A2(n_86),
.B(n_92),
.Y(n_993)
);

AND2x2_ASAP7_75t_SL g994 ( 
.A(n_808),
.B(n_115),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_807),
.A2(n_118),
.B(n_126),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_SL g996 ( 
.A1(n_835),
.A2(n_131),
.B(n_138),
.C(n_139),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_848),
.Y(n_997)
);

INVxp67_ASAP7_75t_SL g998 ( 
.A(n_850),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_869),
.B(n_157),
.Y(n_999)
);

BUFx2_ASAP7_75t_SL g1000 ( 
.A(n_805),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_923),
.A2(n_815),
.B(n_810),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_859),
.A2(n_952),
.B(n_844),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_856),
.B(n_872),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_838),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_915),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_805),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_R g1007 ( 
.A(n_823),
.B(n_855),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_SL g1008 ( 
.A1(n_879),
.A2(n_891),
.B1(n_862),
.B2(n_908),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_863),
.B(n_856),
.Y(n_1009)
);

BUFx8_ASAP7_75t_L g1010 ( 
.A(n_880),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_804),
.B(n_813),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_936),
.Y(n_1012)
);

AO32x1_ASAP7_75t_L g1013 ( 
.A1(n_843),
.A2(n_834),
.A3(n_817),
.B1(n_861),
.B2(n_945),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_847),
.A2(n_816),
.B1(n_822),
.B2(n_801),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_928),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_872),
.B(n_870),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_896),
.B(n_809),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_812),
.B(n_897),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_841),
.A2(n_853),
.B(n_806),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_825),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_880),
.B(n_912),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_SL g1022 ( 
.A(n_904),
.B(n_905),
.Y(n_1022)
);

AOI21x1_ASAP7_75t_L g1023 ( 
.A1(n_858),
.A2(n_874),
.B(n_894),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_949),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_795),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_803),
.Y(n_1026)
);

OR2x6_ASAP7_75t_L g1027 ( 
.A(n_795),
.B(n_904),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_911),
.B(n_933),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_884),
.A2(n_883),
.B1(n_881),
.B2(n_820),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_946),
.B(n_826),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_839),
.B(n_864),
.Y(n_1031)
);

OR2x6_ASAP7_75t_L g1032 ( 
.A(n_795),
.B(n_905),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_796),
.A2(n_792),
.B1(n_941),
.B2(n_932),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_951),
.B(n_878),
.Y(n_1034)
);

NOR3xp33_ASAP7_75t_SL g1035 ( 
.A(n_920),
.B(n_877),
.C(n_886),
.Y(n_1035)
);

BUFx8_ASAP7_75t_SL g1036 ( 
.A(n_912),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_951),
.B(n_888),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_836),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_794),
.A2(n_831),
.B(n_845),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_912),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_892),
.A2(n_854),
.B1(n_895),
.B2(n_882),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_865),
.B(n_907),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_912),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_830),
.A2(n_845),
.B(n_811),
.Y(n_1044)
);

INVxp67_ASAP7_75t_L g1045 ( 
.A(n_819),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_932),
.A2(n_832),
.B1(n_942),
.B2(n_937),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_882),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_944),
.A2(n_829),
.B(n_849),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_931),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_835),
.B(n_855),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_927),
.A2(n_947),
.B1(n_930),
.B2(n_928),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_931),
.B(n_940),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_940),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_913),
.B(n_842),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_851),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_938),
.A2(n_944),
.B(n_939),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_935),
.B(n_950),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_903),
.B(n_924),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_876),
.Y(n_1059)
);

OR2x6_ASAP7_75t_L g1060 ( 
.A(n_943),
.B(n_889),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_SL g1061 ( 
.A(n_909),
.B(n_893),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_898),
.B(n_919),
.Y(n_1062)
);

NOR3xp33_ASAP7_75t_L g1063 ( 
.A(n_953),
.B(n_929),
.C(n_925),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_910),
.B(n_914),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_916),
.B(n_906),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_R g1066 ( 
.A(n_871),
.B(n_589),
.Y(n_1066)
);

AOI21x1_ASAP7_75t_L g1067 ( 
.A1(n_840),
.A2(n_859),
.B(n_857),
.Y(n_1067)
);

NOR2xp67_ASAP7_75t_SL g1068 ( 
.A(n_862),
.B(n_498),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_821),
.A2(n_875),
.B1(n_684),
.B2(n_682),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_900),
.B(n_506),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_873),
.B(n_718),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_873),
.B(n_718),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_866),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_873),
.B(n_718),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_821),
.A2(n_632),
.B(n_657),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_793),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_821),
.A2(n_632),
.B(n_657),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_857),
.A2(n_859),
.B(n_952),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_821),
.A2(n_632),
.B(n_657),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_793),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_827),
.Y(n_1081)
);

NAND3xp33_ASAP7_75t_L g1082 ( 
.A(n_922),
.B(n_636),
.C(n_469),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_793),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_821),
.A2(n_632),
.B(n_657),
.Y(n_1084)
);

AND2x4_ASAP7_75t_SL g1085 ( 
.A(n_891),
.B(n_452),
.Y(n_1085)
);

BUFx4f_ASAP7_75t_L g1086 ( 
.A(n_960),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_988),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1076),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1075),
.A2(n_1079),
.B(n_1077),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1084),
.A2(n_1001),
.B(n_963),
.Y(n_1090)
);

INVxp67_ASAP7_75t_SL g1091 ( 
.A(n_991),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1080),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_SL g1093 ( 
.A1(n_986),
.A2(n_1050),
.B(n_996),
.C(n_1029),
.Y(n_1093)
);

OR2x6_ASAP7_75t_L g1094 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_1005),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1083),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_1036),
.Y(n_1097)
);

INVxp67_ASAP7_75t_L g1098 ( 
.A(n_991),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1014),
.B(n_1069),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1044),
.A2(n_994),
.B(n_1065),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_1085),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_1071),
.A2(n_1072),
.B(n_1074),
.C(n_987),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_994),
.A2(n_1039),
.B(n_1062),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_1070),
.B(n_1073),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_981),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1070),
.B(n_960),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_965),
.A2(n_989),
.B1(n_1009),
.B2(n_1018),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1014),
.B(n_965),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1056),
.A2(n_1048),
.B(n_993),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1004),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_972),
.A2(n_1023),
.B(n_962),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_977),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1015),
.B(n_970),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1054),
.A2(n_957),
.B(n_1058),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_999),
.B(n_1053),
.Y(n_1115)
);

INVx3_ASAP7_75t_SL g1116 ( 
.A(n_1081),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1020),
.B(n_1017),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_992),
.A2(n_995),
.B(n_979),
.Y(n_1118)
);

NAND2xp33_ASAP7_75t_L g1119 ( 
.A(n_956),
.B(n_1035),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1011),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_1010),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1060),
.A2(n_1064),
.B(n_1028),
.Y(n_1122)
);

INVxp67_ASAP7_75t_L g1123 ( 
.A(n_982),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1033),
.A2(n_978),
.B(n_1046),
.Y(n_1124)
);

OR2x6_ASAP7_75t_L g1125 ( 
.A(n_1003),
.B(n_1008),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1022),
.A2(n_958),
.B(n_955),
.Y(n_1126)
);

CKINVDCx11_ASAP7_75t_R g1127 ( 
.A(n_973),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_954),
.A2(n_1013),
.B(n_1061),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_973),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1013),
.A2(n_1021),
.B(n_959),
.Y(n_1130)
);

AOI221x1_ASAP7_75t_L g1131 ( 
.A1(n_1063),
.A2(n_975),
.B1(n_968),
.B2(n_980),
.C(n_1057),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1013),
.A2(n_1051),
.B(n_967),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_976),
.A2(n_974),
.B(n_1055),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_1003),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_961),
.B(n_1016),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_956),
.A2(n_990),
.B1(n_983),
.B2(n_1035),
.Y(n_1136)
);

BUFx10_ASAP7_75t_L g1137 ( 
.A(n_1006),
.Y(n_1137)
);

AOI221x1_ASAP7_75t_L g1138 ( 
.A1(n_1063),
.A2(n_1016),
.B1(n_964),
.B2(n_1009),
.C(n_1042),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1041),
.A2(n_1051),
.B1(n_998),
.B2(n_966),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1038),
.B(n_1030),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1026),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_1027),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1010),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1045),
.A2(n_1026),
.B(n_1047),
.C(n_971),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_973),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1047),
.B(n_1031),
.Y(n_1146)
);

AOI221xp5_ASAP7_75t_SL g1147 ( 
.A1(n_1045),
.A2(n_1034),
.B1(n_1037),
.B2(n_1024),
.C(n_1000),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1040),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_969),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1059),
.B(n_1025),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1059),
.A2(n_1043),
.B(n_1025),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1068),
.B(n_1066),
.Y(n_1152)
);

AO21x2_ASAP7_75t_L g1153 ( 
.A1(n_1007),
.A2(n_1066),
.B(n_973),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_997),
.A2(n_1027),
.B1(n_1032),
.B2(n_985),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1007),
.A2(n_1067),
.B(n_1078),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1075),
.A2(n_821),
.B(n_1077),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_965),
.A2(n_506),
.B1(n_501),
.B2(n_429),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1052),
.B(n_1049),
.Y(n_1158)
);

BUFx8_ASAP7_75t_L g1159 ( 
.A(n_971),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_977),
.Y(n_1160)
);

BUFx10_ASAP7_75t_L g1161 ( 
.A(n_1004),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_988),
.Y(n_1162)
);

AO21x2_ASAP7_75t_L g1163 ( 
.A1(n_1067),
.A2(n_1078),
.B(n_1019),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1004),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_988),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1075),
.A2(n_821),
.B(n_1077),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1012),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1067),
.A2(n_1078),
.B(n_1002),
.Y(n_1168)
);

AO22x1_ASAP7_75t_L g1169 ( 
.A1(n_960),
.A2(n_506),
.B1(n_922),
.B2(n_429),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1067),
.A2(n_1078),
.B(n_1002),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1070),
.B(n_654),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_SL g1172 ( 
.A1(n_963),
.A2(n_1082),
.B(n_921),
.C(n_986),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_SL g1173 ( 
.A(n_965),
.B(n_994),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1014),
.B(n_821),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1067),
.A2(n_1078),
.B(n_1002),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1004),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1067),
.A2(n_1078),
.B(n_1002),
.Y(n_1177)
);

INVx4_ASAP7_75t_L g1178 ( 
.A(n_1036),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_965),
.A2(n_506),
.B1(n_501),
.B2(n_429),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_988),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1082),
.A2(n_922),
.B1(n_636),
.B2(n_994),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_958),
.A2(n_918),
.A3(n_828),
.B(n_858),
.Y(n_1182)
);

NAND2x1p5_ASAP7_75t_L g1183 ( 
.A(n_1053),
.B(n_1049),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1014),
.B(n_821),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1075),
.A2(n_821),
.B(n_1077),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1067),
.A2(n_1078),
.B(n_1002),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1075),
.A2(n_821),
.B(n_1077),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1005),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1005),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1071),
.B(n_1072),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_963),
.A2(n_1082),
.B(n_1077),
.Y(n_1191)
);

CKINVDCx6p67_ASAP7_75t_R g1192 ( 
.A(n_960),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1075),
.A2(n_821),
.B(n_1077),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_SL g1194 ( 
.A(n_965),
.B(n_994),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1067),
.A2(n_1078),
.B(n_1002),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1075),
.A2(n_821),
.B(n_1077),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1082),
.A2(n_922),
.B1(n_636),
.B2(n_994),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1014),
.B(n_821),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_963),
.A2(n_1082),
.B(n_1077),
.Y(n_1199)
);

INVx2_ASAP7_75t_SL g1200 ( 
.A(n_1005),
.Y(n_1200)
);

OAI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1082),
.A2(n_507),
.B1(n_429),
.B2(n_506),
.Y(n_1201)
);

AOI221x1_ASAP7_75t_L g1202 ( 
.A1(n_984),
.A2(n_1082),
.B1(n_488),
.B2(n_986),
.C(n_963),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_958),
.A2(n_918),
.A3(n_828),
.B(n_858),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_977),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_977),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1075),
.A2(n_821),
.B(n_1077),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1075),
.A2(n_821),
.B(n_1077),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_958),
.A2(n_918),
.A3(n_828),
.B(n_858),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1073),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_1036),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1087),
.Y(n_1211)
);

CKINVDCx6p67_ASAP7_75t_R g1212 ( 
.A(n_1116),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1157),
.A2(n_1179),
.B1(n_1201),
.B2(n_1173),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1171),
.B(n_1104),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_1210),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1112),
.Y(n_1216)
);

CKINVDCx11_ASAP7_75t_R g1217 ( 
.A(n_1161),
.Y(n_1217)
);

INVx6_ASAP7_75t_L g1218 ( 
.A(n_1159),
.Y(n_1218)
);

INVx6_ASAP7_75t_L g1219 ( 
.A(n_1159),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1088),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_1153),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1127),
.Y(n_1222)
);

INVx1_ASAP7_75t_SL g1223 ( 
.A(n_1209),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1173),
.A2(n_1194),
.B1(n_1181),
.B2(n_1197),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1194),
.A2(n_1119),
.B1(n_1136),
.B2(n_1107),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1136),
.A2(n_1169),
.B1(n_1115),
.B2(n_1106),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1092),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1110),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1158),
.Y(n_1229)
);

CKINVDCx11_ASAP7_75t_R g1230 ( 
.A(n_1161),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1160),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1096),
.Y(n_1232)
);

BUFx12f_ASAP7_75t_L g1233 ( 
.A(n_1164),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1108),
.A2(n_1099),
.B1(n_1103),
.B2(n_1139),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1162),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1165),
.Y(n_1236)
);

BUFx2_ASAP7_75t_SL g1237 ( 
.A(n_1210),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1095),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1210),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1180),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1108),
.A2(n_1139),
.B1(n_1117),
.B2(n_1135),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1209),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1174),
.A2(n_1184),
.B1(n_1198),
.B2(n_1120),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1113),
.B(n_1098),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1174),
.A2(n_1184),
.B1(n_1198),
.B2(n_1140),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1152),
.A2(n_1101),
.B1(n_1125),
.B2(n_1154),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1140),
.A2(n_1191),
.B1(n_1199),
.B2(n_1167),
.Y(n_1247)
);

INVx5_ASAP7_75t_L g1248 ( 
.A(n_1142),
.Y(n_1248)
);

INVx6_ASAP7_75t_L g1249 ( 
.A(n_1142),
.Y(n_1249)
);

BUFx4f_ASAP7_75t_SL g1250 ( 
.A(n_1188),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1204),
.B(n_1205),
.Y(n_1251)
);

INVx6_ASAP7_75t_L g1252 ( 
.A(n_1142),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1094),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_1176),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1125),
.A2(n_1132),
.B1(n_1124),
.B2(n_1154),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1125),
.A2(n_1134),
.B1(n_1100),
.B2(n_1126),
.Y(n_1256)
);

INVx6_ASAP7_75t_L g1257 ( 
.A(n_1094),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1102),
.B(n_1134),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1189),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1183),
.A2(n_1141),
.B1(n_1149),
.B2(n_1128),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1146),
.A2(n_1094),
.B1(n_1090),
.B2(n_1148),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1146),
.B(n_1123),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1121),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1150),
.Y(n_1264)
);

CKINVDCx11_ASAP7_75t_R g1265 ( 
.A(n_1137),
.Y(n_1265)
);

INVx5_ASAP7_75t_L g1266 ( 
.A(n_1143),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1200),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1086),
.A2(n_1192),
.B1(n_1147),
.B2(n_1105),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1144),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1137),
.Y(n_1270)
);

BUFx12f_ASAP7_75t_L g1271 ( 
.A(n_1097),
.Y(n_1271)
);

BUFx4f_ASAP7_75t_SL g1272 ( 
.A(n_1097),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1114),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1183),
.A2(n_1122),
.B1(n_1130),
.B2(n_1086),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1178),
.B(n_1151),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1151),
.A2(n_1131),
.B1(n_1202),
.B2(n_1178),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1156),
.A2(n_1166),
.B1(n_1207),
.B2(n_1206),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1129),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1093),
.A2(n_1138),
.B1(n_1187),
.B2(n_1185),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1193),
.A2(n_1196),
.B1(n_1172),
.B2(n_1089),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1155),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1145),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1133),
.A2(n_1118),
.B1(n_1163),
.B2(n_1111),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1163),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1182),
.A2(n_1208),
.B1(n_1203),
.B2(n_1109),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1168),
.A2(n_1170),
.B(n_1175),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1203),
.A2(n_1208),
.B1(n_1186),
.B2(n_1195),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1177),
.Y(n_1288)
);

BUFx12f_ASAP7_75t_L g1289 ( 
.A(n_1161),
.Y(n_1289)
);

CKINVDCx11_ASAP7_75t_R g1290 ( 
.A(n_1116),
.Y(n_1290)
);

CKINVDCx8_ASAP7_75t_R g1291 ( 
.A(n_1210),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1087),
.Y(n_1292)
);

CKINVDCx11_ASAP7_75t_R g1293 ( 
.A(n_1116),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1110),
.Y(n_1294)
);

BUFx4f_ASAP7_75t_SL g1295 ( 
.A(n_1116),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1087),
.Y(n_1296)
);

INVx8_ASAP7_75t_L g1297 ( 
.A(n_1210),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1181),
.A2(n_1197),
.B1(n_1082),
.B2(n_965),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1181),
.A2(n_1197),
.B1(n_1082),
.B2(n_965),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1110),
.Y(n_1300)
);

CKINVDCx6p67_ASAP7_75t_R g1301 ( 
.A(n_1116),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1087),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1157),
.A2(n_1179),
.B1(n_506),
.B2(n_1201),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1087),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1173),
.A2(n_1194),
.B1(n_330),
.B2(n_328),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1127),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1173),
.A2(n_1194),
.B1(n_330),
.B2(n_328),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1157),
.A2(n_1179),
.B1(n_506),
.B2(n_1201),
.Y(n_1308)
);

INVx5_ASAP7_75t_L g1309 ( 
.A(n_1142),
.Y(n_1309)
);

BUFx12f_ASAP7_75t_L g1310 ( 
.A(n_1161),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_1161),
.Y(n_1311)
);

BUFx2_ASAP7_75t_SL g1312 ( 
.A(n_1210),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1087),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1157),
.A2(n_1179),
.B1(n_506),
.B2(n_1201),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1087),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1098),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1171),
.B(n_1104),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1190),
.B(n_1117),
.Y(n_1318)
);

INVxp67_ASAP7_75t_SL g1319 ( 
.A(n_1091),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1173),
.A2(n_1194),
.B1(n_1197),
.B2(n_1181),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_1104),
.Y(n_1321)
);

INVxp67_ASAP7_75t_SL g1322 ( 
.A(n_1091),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1190),
.B(n_1117),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1190),
.B(n_1117),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1265),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1211),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1220),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1319),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_SL g1329 ( 
.A(n_1291),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1303),
.A2(n_1308),
.B1(n_1314),
.B2(n_1213),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1227),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1297),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1322),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1232),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1235),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1285),
.A2(n_1277),
.B(n_1287),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1264),
.B(n_1245),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1236),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1265),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1275),
.B(n_1215),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1286),
.A2(n_1277),
.B(n_1283),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1240),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1292),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1316),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1296),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1302),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1304),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1318),
.B(n_1323),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1313),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1315),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1225),
.A2(n_1224),
.B1(n_1299),
.B2(n_1298),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1297),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1254),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1234),
.B(n_1245),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1321),
.B(n_1267),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1324),
.B(n_1262),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1234),
.B(n_1243),
.Y(n_1357)
);

AOI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1284),
.A2(n_1288),
.B(n_1281),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1216),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1258),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1231),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1243),
.B(n_1241),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1248),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1213),
.A2(n_1308),
.B1(n_1314),
.B2(n_1303),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1241),
.B(n_1247),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1273),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1221),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1221),
.Y(n_1368)
);

AO21x1_ASAP7_75t_L g1369 ( 
.A1(n_1320),
.A2(n_1226),
.B(n_1269),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1247),
.Y(n_1370)
);

AO31x2_ASAP7_75t_L g1371 ( 
.A1(n_1278),
.A2(n_1282),
.A3(n_1279),
.B(n_1280),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1223),
.Y(n_1372)
);

OR2x6_ASAP7_75t_L g1373 ( 
.A(n_1253),
.B(n_1257),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1242),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1263),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1251),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1244),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1214),
.B(n_1317),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1224),
.B(n_1225),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1246),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1276),
.B(n_1229),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1261),
.B(n_1255),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1260),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1276),
.B(n_1229),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1256),
.B(n_1274),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1238),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1305),
.A2(n_1307),
.B1(n_1253),
.B2(n_1257),
.Y(n_1387)
);

BUFx8_ASAP7_75t_SL g1388 ( 
.A(n_1254),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1238),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_1290),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1333),
.B(n_1222),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1338),
.Y(n_1392)
);

BUFx4f_ASAP7_75t_L g1393 ( 
.A(n_1363),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1356),
.B(n_1268),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1336),
.B(n_1306),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1328),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1353),
.B(n_1250),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1336),
.B(n_1306),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1388),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1336),
.B(n_1222),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1336),
.B(n_1239),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1338),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1341),
.A2(n_1270),
.B(n_1252),
.Y(n_1403)
);

A2O1A1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1330),
.A2(n_1259),
.B(n_1266),
.C(n_1312),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1333),
.B(n_1237),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1344),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1389),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_SL g1408 ( 
.A1(n_1353),
.A2(n_1290),
.B(n_1293),
.C(n_1230),
.Y(n_1408)
);

OAI211xp5_ASAP7_75t_L g1409 ( 
.A1(n_1351),
.A2(n_1217),
.B(n_1230),
.C(n_1293),
.Y(n_1409)
);

INVxp67_ASAP7_75t_L g1410 ( 
.A(n_1355),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1340),
.B(n_1248),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1360),
.B(n_1259),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1364),
.A2(n_1218),
.B1(n_1219),
.B2(n_1272),
.Y(n_1413)
);

NOR2x1_ASAP7_75t_R g1414 ( 
.A(n_1390),
.B(n_1218),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1361),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1354),
.A2(n_1294),
.B(n_1300),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1342),
.B(n_1343),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1343),
.B(n_1212),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1348),
.B(n_1301),
.Y(n_1419)
);

OA21x2_ASAP7_75t_L g1420 ( 
.A1(n_1341),
.A2(n_1249),
.B(n_1309),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1365),
.A2(n_1218),
.B1(n_1219),
.B2(n_1250),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1377),
.B(n_1219),
.Y(n_1422)
);

OAI211xp5_ASAP7_75t_L g1423 ( 
.A1(n_1354),
.A2(n_1217),
.B(n_1228),
.C(n_1272),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1345),
.B(n_1271),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1345),
.B(n_1271),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1357),
.A2(n_1295),
.B(n_1289),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_R g1427 ( 
.A(n_1390),
.B(n_1295),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1346),
.B(n_1310),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1347),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1382),
.A2(n_1310),
.B(n_1311),
.C(n_1249),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1347),
.B(n_1311),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1349),
.B(n_1233),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1340),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1372),
.B(n_1374),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1349),
.B(n_1350),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1369),
.A2(n_1379),
.B1(n_1382),
.B2(n_1357),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1350),
.B(n_1326),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1337),
.B(n_1362),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1327),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1379),
.A2(n_1385),
.B(n_1370),
.C(n_1383),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1378),
.B(n_1359),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1331),
.B(n_1334),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1385),
.A2(n_1383),
.B(n_1384),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1335),
.B(n_1376),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1392),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1392),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1443),
.A2(n_1395),
.B1(n_1398),
.B2(n_1400),
.Y(n_1447)
);

OAI222xp33_ASAP7_75t_L g1448 ( 
.A1(n_1436),
.A2(n_1380),
.B1(n_1381),
.B2(n_1378),
.C1(n_1387),
.C2(n_1373),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1402),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1438),
.B(n_1371),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1436),
.A2(n_1329),
.B1(n_1386),
.B2(n_1375),
.Y(n_1451)
);

INVx4_ASAP7_75t_L g1452 ( 
.A(n_1393),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1396),
.B(n_1371),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1407),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1406),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1438),
.B(n_1371),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1391),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1417),
.B(n_1371),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1415),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1395),
.B(n_1371),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1398),
.B(n_1400),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1433),
.Y(n_1462)
);

AOI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1401),
.A2(n_1358),
.B(n_1367),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1433),
.B(n_1366),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1417),
.B(n_1366),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1429),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1435),
.B(n_1437),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1437),
.B(n_1442),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1411),
.B(n_1368),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1401),
.B(n_1367),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1444),
.B(n_1368),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1439),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1439),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1444),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1434),
.B(n_1359),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1466),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1466),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1467),
.B(n_1403),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1463),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1445),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1458),
.B(n_1441),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1459),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1458),
.B(n_1403),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1459),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1467),
.B(n_1403),
.Y(n_1486)
);

INVx5_ASAP7_75t_L g1487 ( 
.A(n_1460),
.Y(n_1487)
);

NAND4xp25_ASAP7_75t_L g1488 ( 
.A(n_1451),
.B(n_1409),
.C(n_1416),
.D(n_1418),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1455),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1445),
.Y(n_1490)
);

CKINVDCx14_ASAP7_75t_R g1491 ( 
.A(n_1475),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1470),
.Y(n_1492)
);

NOR2xp67_ASAP7_75t_L g1493 ( 
.A(n_1453),
.B(n_1423),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1455),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1446),
.Y(n_1495)
);

NAND3xp33_ASAP7_75t_SL g1496 ( 
.A(n_1453),
.B(n_1440),
.C(n_1391),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1467),
.B(n_1403),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1450),
.B(n_1405),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_R g1499 ( 
.A(n_1452),
.B(n_1399),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1470),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1465),
.B(n_1412),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1447),
.A2(n_1394),
.B1(n_1410),
.B2(n_1404),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1461),
.B(n_1420),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1446),
.Y(n_1504)
);

OAI31xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1460),
.A2(n_1413),
.A3(n_1424),
.B(n_1425),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1450),
.B(n_1456),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1461),
.B(n_1420),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1470),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1449),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1509),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1509),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1480),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1487),
.B(n_1462),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1487),
.B(n_1461),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1480),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1487),
.B(n_1462),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1487),
.B(n_1460),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1483),
.Y(n_1518)
);

NOR3xp33_ASAP7_75t_SL g1519 ( 
.A(n_1488),
.B(n_1399),
.C(n_1339),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1482),
.B(n_1468),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1490),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1487),
.B(n_1471),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1483),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1485),
.B(n_1472),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1485),
.B(n_1489),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1489),
.B(n_1472),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1487),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1487),
.B(n_1471),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1478),
.B(n_1474),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1478),
.B(n_1457),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1494),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1482),
.B(n_1468),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1486),
.B(n_1457),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1486),
.B(n_1464),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1508),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1490),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1482),
.B(n_1498),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1494),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1495),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1498),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1486),
.B(n_1464),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1495),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1497),
.B(n_1464),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1476),
.B(n_1473),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1503),
.B(n_1469),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1504),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1517),
.B(n_1491),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1512),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1527),
.A2(n_1502),
.B(n_1481),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1534),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1520),
.B(n_1498),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1520),
.B(n_1532),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1512),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1532),
.B(n_1493),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1537),
.B(n_1476),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1534),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1518),
.B(n_1493),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1515),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1515),
.Y(n_1559)
);

OA21x2_ASAP7_75t_L g1560 ( 
.A1(n_1510),
.A2(n_1479),
.B(n_1484),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1535),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1535),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1517),
.B(n_1514),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1535),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1521),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1518),
.B(n_1497),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1521),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1517),
.B(n_1491),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1537),
.B(n_1477),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1513),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1540),
.B(n_1477),
.Y(n_1571)
);

OAI31xp33_ASAP7_75t_L g1572 ( 
.A1(n_1530),
.A2(n_1502),
.A3(n_1448),
.B(n_1484),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1530),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1519),
.A2(n_1481),
.B1(n_1492),
.B2(n_1447),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1519),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1530),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1538),
.B(n_1497),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1536),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1534),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1525),
.B(n_1538),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1533),
.A2(n_1496),
.B1(n_1488),
.B2(n_1450),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1541),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1536),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1533),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1539),
.Y(n_1585)
);

AOI311xp33_ASAP7_75t_L g1586 ( 
.A1(n_1510),
.A2(n_1408),
.A3(n_1504),
.B(n_1397),
.C(n_1448),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1525),
.B(n_1506),
.Y(n_1587)
);

INVx4_ASAP7_75t_L g1588 ( 
.A(n_1513),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1527),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1550),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1552),
.B(n_1524),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1554),
.B(n_1581),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1548),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1557),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1552),
.B(n_1524),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1581),
.B(n_1523),
.Y(n_1596)
);

AOI221x1_ASAP7_75t_SL g1597 ( 
.A1(n_1574),
.A2(n_1511),
.B1(n_1526),
.B2(n_1545),
.C(n_1419),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1547),
.B(n_1514),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1550),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1548),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1549),
.B(n_1531),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_1580),
.B(n_1421),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1580),
.B(n_1533),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1551),
.B(n_1500),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1547),
.B(n_1514),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1551),
.B(n_1526),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1555),
.B(n_1500),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1575),
.B(n_1325),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1556),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1587),
.B(n_1511),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1568),
.B(n_1545),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1568),
.B(n_1545),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1587),
.B(n_1501),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1555),
.B(n_1569),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1553),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1586),
.B(n_1479),
.C(n_1505),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1569),
.B(n_1529),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1571),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1571),
.B(n_1501),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1573),
.B(n_1529),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1553),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1586),
.B(n_1527),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1573),
.B(n_1544),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1572),
.A2(n_1496),
.B(n_1503),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1573),
.A2(n_1456),
.B1(n_1503),
.B2(n_1507),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1593),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1616),
.A2(n_1624),
.B1(n_1592),
.B2(n_1622),
.Y(n_1627)
);

AOI221xp5_ASAP7_75t_L g1628 ( 
.A1(n_1597),
.A2(n_1577),
.B1(n_1566),
.B2(n_1479),
.C(n_1562),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1600),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1608),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1615),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1618),
.B(n_1558),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1602),
.Y(n_1633)
);

AOI221xp5_ASAP7_75t_L g1634 ( 
.A1(n_1596),
.A2(n_1594),
.B1(n_1622),
.B2(n_1601),
.C(n_1621),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1602),
.A2(n_1584),
.B1(n_1576),
.B2(n_1556),
.Y(n_1635)
);

NAND2x1p5_ASAP7_75t_L g1636 ( 
.A(n_1608),
.B(n_1588),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1614),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1591),
.B(n_1576),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1610),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1602),
.A2(n_1456),
.B1(n_1507),
.B2(n_1560),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1590),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1603),
.A2(n_1560),
.B(n_1505),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1590),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1599),
.Y(n_1644)
);

OAI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1625),
.A2(n_1506),
.B1(n_1576),
.B2(n_1584),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1599),
.B(n_1558),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1594),
.B(n_1584),
.Y(n_1647)
);

OAI31xp33_ASAP7_75t_L g1648 ( 
.A1(n_1595),
.A2(n_1506),
.A3(n_1507),
.B(n_1561),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1598),
.B(n_1588),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1598),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1611),
.B(n_1579),
.Y(n_1651)
);

AOI21xp33_ASAP7_75t_L g1652 ( 
.A1(n_1627),
.A2(n_1609),
.B(n_1623),
.Y(n_1652)
);

NAND2xp33_ASAP7_75t_L g1653 ( 
.A(n_1636),
.B(n_1637),
.Y(n_1653)
);

INVxp67_ASAP7_75t_L g1654 ( 
.A(n_1633),
.Y(n_1654)
);

AOI311xp33_ASAP7_75t_L g1655 ( 
.A1(n_1634),
.A2(n_1620),
.A3(n_1604),
.B(n_1583),
.C(n_1578),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1650),
.B(n_1609),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1642),
.A2(n_1589),
.B(n_1606),
.Y(n_1657)
);

AOI222xp33_ASAP7_75t_L g1658 ( 
.A1(n_1628),
.A2(n_1617),
.B1(n_1564),
.B2(n_1561),
.C1(n_1562),
.C2(n_1607),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1640),
.B(n_1588),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1635),
.A2(n_1589),
.B(n_1611),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1641),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1639),
.B(n_1613),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1647),
.B(n_1619),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1643),
.Y(n_1664)
);

AOI222xp33_ASAP7_75t_L g1665 ( 
.A1(n_1635),
.A2(n_1561),
.B1(n_1562),
.B2(n_1564),
.C1(n_1578),
.C2(n_1567),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1636),
.A2(n_1612),
.B1(n_1579),
.B2(n_1582),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1651),
.B(n_1582),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1630),
.A2(n_1560),
.B1(n_1564),
.B2(n_1612),
.Y(n_1668)
);

AOI21xp33_ASAP7_75t_L g1669 ( 
.A1(n_1632),
.A2(n_1560),
.B(n_1559),
.Y(n_1669)
);

AOI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1645),
.A2(n_1585),
.B1(n_1583),
.B2(n_1559),
.C(n_1567),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1644),
.Y(n_1671)
);

OA22x2_ASAP7_75t_L g1672 ( 
.A1(n_1657),
.A2(n_1649),
.B1(n_1632),
.B2(n_1626),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1653),
.Y(n_1673)
);

A2O1A1Ixp33_ASAP7_75t_SL g1674 ( 
.A1(n_1669),
.A2(n_1629),
.B(n_1631),
.C(n_1646),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1654),
.B(n_1638),
.Y(n_1675)
);

NAND2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1671),
.B(n_1414),
.Y(n_1676)
);

O2A1O1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1652),
.A2(n_1654),
.B(n_1664),
.C(n_1661),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1656),
.B(n_1646),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1662),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1663),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1667),
.B(n_1648),
.Y(n_1681)
);

AOI21xp33_ASAP7_75t_L g1682 ( 
.A1(n_1665),
.A2(n_1658),
.B(n_1668),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1660),
.Y(n_1683)
);

AOI31xp33_ASAP7_75t_SL g1684 ( 
.A1(n_1655),
.A2(n_1414),
.A3(n_1427),
.B(n_1325),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1675),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_SL g1686 ( 
.A(n_1674),
.B(n_1670),
.C(n_1666),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1678),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1677),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1682),
.A2(n_1659),
.B1(n_1605),
.B2(n_1421),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1680),
.B(n_1605),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1679),
.Y(n_1691)
);

OR2x6_ASAP7_75t_L g1692 ( 
.A(n_1676),
.B(n_1339),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1673),
.B(n_1563),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1672),
.A2(n_1585),
.B(n_1565),
.Y(n_1694)
);

NOR3xp33_ASAP7_75t_L g1695 ( 
.A(n_1688),
.B(n_1685),
.C(n_1686),
.Y(n_1695)
);

O2A1O1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1687),
.A2(n_1683),
.B(n_1684),
.C(n_1691),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1694),
.A2(n_1681),
.B1(n_1684),
.B2(n_1565),
.C(n_1570),
.Y(n_1697)
);

NOR3xp33_ASAP7_75t_SL g1698 ( 
.A(n_1690),
.B(n_1426),
.C(n_1430),
.Y(n_1698)
);

AOI211xp5_ASAP7_75t_L g1699 ( 
.A1(n_1693),
.A2(n_1570),
.B(n_1563),
.C(n_1432),
.Y(n_1699)
);

AOI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1695),
.A2(n_1689),
.B1(n_1692),
.B2(n_1570),
.C(n_1588),
.Y(n_1700)
);

OAI211xp5_ASAP7_75t_L g1701 ( 
.A1(n_1696),
.A2(n_1692),
.B(n_1570),
.C(n_1499),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1699),
.B(n_1697),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1698),
.A2(n_1432),
.B1(n_1431),
.B2(n_1428),
.C(n_1425),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1695),
.Y(n_1704)
);

NOR3xp33_ASAP7_75t_L g1705 ( 
.A(n_1695),
.B(n_1424),
.C(n_1428),
.Y(n_1705)
);

NAND4xp75_ASAP7_75t_L g1706 ( 
.A(n_1700),
.B(n_1431),
.C(n_1418),
.D(n_1516),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_L g1707 ( 
.A(n_1704),
.B(n_1701),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1702),
.Y(n_1708)
);

NAND4xp75_ASAP7_75t_L g1709 ( 
.A(n_1703),
.B(n_1516),
.C(n_1528),
.D(n_1522),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1705),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1707),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1708),
.B(n_1710),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1706),
.A2(n_1545),
.B1(n_1541),
.B2(n_1543),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1711),
.A2(n_1709),
.B1(n_1545),
.B2(n_1543),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1714),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1715),
.B(n_1712),
.Y(n_1716)
);

INVx3_ASAP7_75t_SL g1717 ( 
.A(n_1715),
.Y(n_1717)
);

AO22x2_ASAP7_75t_L g1718 ( 
.A1(n_1716),
.A2(n_1717),
.B1(n_1713),
.B2(n_1546),
.Y(n_1718)
);

INVx6_ASAP7_75t_L g1719 ( 
.A(n_1716),
.Y(n_1719)
);

OA21x2_ASAP7_75t_L g1720 ( 
.A1(n_1719),
.A2(n_1544),
.B(n_1542),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1720),
.B(n_1718),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1721),
.Y(n_1722)
);

AOI22x1_ASAP7_75t_L g1723 ( 
.A1(n_1722),
.A2(n_1546),
.B1(n_1539),
.B2(n_1542),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1723),
.A2(n_1422),
.B1(n_1541),
.B2(n_1543),
.C(n_1529),
.Y(n_1724)
);

AOI211xp5_ASAP7_75t_L g1725 ( 
.A1(n_1724),
.A2(n_1499),
.B(n_1332),
.C(n_1352),
.Y(n_1725)
);


endmodule