module real_aes_9082_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_182;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g581 ( .A1(n_0), .A2(n_160), .B(n_582), .C(n_585), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_1), .B(n_526), .Y(n_586) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g194 ( .A(n_3), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_4), .B(n_152), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_5), .A2(n_495), .B(n_520), .Y(n_519) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_6), .A2(n_137), .B(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_7), .A2(n_35), .B1(n_146), .B2(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_8), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_9), .B(n_137), .Y(n_163) );
AND2x6_ASAP7_75t_L g161 ( .A(n_10), .B(n_162), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_11), .A2(n_161), .B(n_485), .C(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g108 ( .A(n_12), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_12), .B(n_36), .Y(n_447) );
INVx1_ASAP7_75t_L g142 ( .A(n_13), .Y(n_142) );
INVx1_ASAP7_75t_L g187 ( .A(n_14), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_15), .B(n_150), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_16), .B(n_152), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_17), .B(n_138), .Y(n_199) );
AO32x2_ASAP7_75t_L g221 ( .A1(n_18), .A2(n_137), .A3(n_167), .B1(n_178), .B2(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_19), .B(n_146), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_20), .B(n_138), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_21), .A2(n_54), .B1(n_146), .B2(n_224), .Y(n_225) );
AOI22xp33_ASAP7_75t_SL g246 ( .A1(n_22), .A2(n_82), .B1(n_146), .B2(n_150), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_23), .B(n_146), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_24), .A2(n_178), .B(n_485), .C(n_546), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_25), .A2(n_178), .B(n_485), .C(n_514), .Y(n_513) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_26), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_27), .B(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_28), .A2(n_495), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_29), .B(n_180), .Y(n_218) );
INVx2_ASAP7_75t_L g148 ( .A(n_30), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_31), .A2(n_497), .B(n_505), .C(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_32), .B(n_146), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_33), .B(n_180), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_34), .B(n_232), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_36), .B(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_37), .B(n_544), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_38), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_39), .A2(n_78), .B1(n_462), .B2(n_463), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g463 ( .A(n_39), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_40), .B(n_152), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_41), .B(n_495), .Y(n_512) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_42), .A2(n_79), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_42), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_43), .A2(n_497), .B(n_499), .C(n_505), .Y(n_496) );
OAI22xp5_ASAP7_75t_SL g460 ( .A1(n_44), .A2(n_461), .B1(n_464), .B2(n_465), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_44), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_45), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g583 ( .A(n_46), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_47), .A2(n_91), .B1(n_224), .B2(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g500 ( .A(n_48), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_49), .B(n_146), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_50), .B(n_146), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_51), .B(n_124), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_51), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_52), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_53), .B(n_158), .Y(n_157) );
AOI22xp33_ASAP7_75t_SL g203 ( .A1(n_55), .A2(n_59), .B1(n_146), .B2(n_150), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_56), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_57), .B(n_146), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_58), .B(n_146), .Y(n_229) );
INVx1_ASAP7_75t_L g162 ( .A(n_60), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_61), .B(n_495), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_62), .B(n_526), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_63), .A2(n_158), .B(n_190), .C(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_64), .B(n_146), .Y(n_195) );
INVx1_ASAP7_75t_L g141 ( .A(n_65), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_66), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_67), .B(n_152), .Y(n_536) );
AO32x2_ASAP7_75t_L g242 ( .A1(n_68), .A2(n_137), .A3(n_178), .B1(n_243), .B2(n_247), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_69), .B(n_153), .Y(n_488) );
INVx1_ASAP7_75t_L g173 ( .A(n_70), .Y(n_173) );
INVx1_ASAP7_75t_L g213 ( .A(n_71), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g580 ( .A(n_72), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_73), .B(n_502), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_74), .A2(n_485), .B(n_505), .C(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_75), .B(n_150), .Y(n_214) );
CKINVDCx16_ASAP7_75t_R g521 ( .A(n_76), .Y(n_521) );
INVx1_ASAP7_75t_L g115 ( .A(n_77), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_78), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_79), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g468 ( .A1(n_79), .A2(n_128), .B1(n_129), .B2(n_439), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_80), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_81), .B(n_501), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_83), .B(n_224), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_84), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_85), .B(n_150), .Y(n_217) );
INVx2_ASAP7_75t_L g139 ( .A(n_86), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_87), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_88), .B(n_177), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_89), .B(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g112 ( .A(n_90), .Y(n_112) );
OR2x2_ASAP7_75t_L g444 ( .A(n_90), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g471 ( .A(n_90), .B(n_446), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_92), .A2(n_103), .B1(n_150), .B2(n_151), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_93), .B(n_495), .Y(n_532) );
INVx1_ASAP7_75t_L g535 ( .A(n_94), .Y(n_535) );
INVxp67_ASAP7_75t_L g524 ( .A(n_95), .Y(n_524) );
AOI222xp33_ASAP7_75t_SL g459 ( .A1(n_96), .A2(n_460), .B1(n_466), .B2(n_759), .C1(n_760), .C2(n_764), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_97), .A2(n_105), .B1(n_116), .B2(n_767), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_98), .B(n_150), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_99), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g481 ( .A(n_100), .Y(n_481) );
INVx1_ASAP7_75t_L g559 ( .A(n_101), .Y(n_559) );
AND2x2_ASAP7_75t_L g507 ( .A(n_102), .B(n_180), .Y(n_507) );
INVx2_ASAP7_75t_L g769 ( .A(n_105), .Y(n_769) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_112), .C(n_113), .Y(n_110) );
AND2x2_ASAP7_75t_L g446 ( .A(n_111), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g758 ( .A(n_112), .B(n_446), .Y(n_758) );
NOR2x2_ASAP7_75t_L g766 ( .A(n_112), .B(n_445), .Y(n_766) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AOI22x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B1(n_456), .B2(n_459), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g458 ( .A(n_120), .Y(n_458) );
AOI211xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_448), .B(n_449), .C(n_453), .Y(n_121) );
NOR3xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_440), .C(n_443), .Y(n_122) );
INVxp67_ASAP7_75t_L g450 ( .A(n_123), .Y(n_450) );
INVx1_ASAP7_75t_L g442 ( .A(n_124), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_129), .B2(n_439), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g439 ( .A(n_129), .Y(n_439) );
NAND2x1p5_ASAP7_75t_L g129 ( .A(n_130), .B(n_363), .Y(n_129) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_321), .Y(n_130) );
NOR4xp25_ASAP7_75t_L g131 ( .A(n_132), .B(n_261), .C(n_297), .D(n_311), .Y(n_131) );
OAI221xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_205), .B1(n_237), .B2(n_248), .C(n_252), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_133), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_181), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_164), .Y(n_135) );
AND2x2_ASAP7_75t_L g258 ( .A(n_136), .B(n_165), .Y(n_258) );
INVx3_ASAP7_75t_L g266 ( .A(n_136), .Y(n_266) );
AND2x2_ASAP7_75t_L g320 ( .A(n_136), .B(n_184), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_136), .B(n_183), .Y(n_356) );
AND2x2_ASAP7_75t_L g414 ( .A(n_136), .B(n_276), .Y(n_414) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_143), .B(n_163), .Y(n_136) );
INVx4_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_137), .A2(n_512), .B(n_513), .Y(n_511) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_137), .Y(n_518) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g167 ( .A(n_138), .Y(n_167) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_139), .B(n_140), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_155), .B(n_161), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_149), .B(n_152), .Y(n_144) );
INVx3_ASAP7_75t_L g212 ( .A(n_146), .Y(n_212) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_146), .Y(n_561) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g224 ( .A(n_147), .Y(n_224) );
BUFx3_ASAP7_75t_L g245 ( .A(n_147), .Y(n_245) );
AND2x6_ASAP7_75t_L g485 ( .A(n_147), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g151 ( .A(n_148), .Y(n_151) );
INVx1_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
INVx2_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_152), .A2(n_170), .B(n_171), .Y(n_169) );
O2A1O1Ixp5_ASAP7_75t_SL g211 ( .A1(n_152), .A2(n_212), .B(n_213), .C(n_214), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_152), .B(n_524), .Y(n_523) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g243 ( .A1(n_153), .A2(n_177), .B1(n_244), .B2(n_246), .Y(n_243) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_154), .Y(n_177) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
INVx1_ASAP7_75t_L g232 ( .A(n_154), .Y(n_232) );
AND2x2_ASAP7_75t_L g483 ( .A(n_154), .B(n_159), .Y(n_483) );
INVx1_ASAP7_75t_L g486 ( .A(n_154), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_160), .Y(n_155) );
INVx2_ASAP7_75t_L g174 ( .A(n_158), .Y(n_174) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_160), .A2(n_174), .B(n_194), .C(n_195), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_160), .A2(n_177), .B1(n_202), .B2(n_203), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_160), .A2(n_177), .B1(n_223), .B2(n_225), .Y(n_222) );
BUFx3_ASAP7_75t_L g178 ( .A(n_161), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_161), .A2(n_186), .B(n_193), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_161), .A2(n_211), .B(n_215), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_161), .A2(n_228), .B(n_233), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_161), .B(n_483), .Y(n_482) );
AND2x4_ASAP7_75t_L g495 ( .A(n_161), .B(n_483), .Y(n_495) );
INVx4_ASAP7_75t_SL g506 ( .A(n_161), .Y(n_506) );
AND2x2_ASAP7_75t_L g249 ( .A(n_164), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g263 ( .A(n_164), .B(n_184), .Y(n_263) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_165), .B(n_184), .Y(n_278) );
AND2x2_ASAP7_75t_L g290 ( .A(n_165), .B(n_266), .Y(n_290) );
OR2x2_ASAP7_75t_L g292 ( .A(n_165), .B(n_250), .Y(n_292) );
AND2x2_ASAP7_75t_L g327 ( .A(n_165), .B(n_250), .Y(n_327) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_165), .Y(n_372) );
INVx1_ASAP7_75t_L g380 ( .A(n_165), .Y(n_380) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_168), .B(n_179), .Y(n_165) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_166), .A2(n_185), .B(n_196), .Y(n_184) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_167), .B(n_491), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_178), .Y(n_168) );
O2A1O1Ixp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_175), .C(n_176), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_174), .A2(n_547), .B(n_548), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_176), .A2(n_234), .B(n_235), .Y(n_233) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx4_ASAP7_75t_L g584 ( .A(n_177), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g200 ( .A(n_178), .B(n_201), .C(n_204), .Y(n_200) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_180), .A2(n_210), .B(n_218), .Y(n_209) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_180), .A2(n_227), .B(n_236), .Y(n_226) );
INVx2_ASAP7_75t_L g247 ( .A(n_180), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_180), .A2(n_494), .B(n_496), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_180), .A2(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g552 ( .A(n_180), .Y(n_552) );
OAI221xp5_ASAP7_75t_L g297 ( .A1(n_181), .A2(n_298), .B1(n_302), .B2(n_306), .C(n_307), .Y(n_297) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g257 ( .A(n_182), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_197), .Y(n_182) );
INVx2_ASAP7_75t_L g256 ( .A(n_183), .Y(n_256) );
AND2x2_ASAP7_75t_L g309 ( .A(n_183), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g328 ( .A(n_183), .B(n_266), .Y(n_328) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g391 ( .A(n_184), .B(n_266), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_189), .C(n_190), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_188), .A2(n_488), .B(n_489), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_188), .A2(n_515), .B(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g558 ( .A1(n_190), .A2(n_559), .B(n_560), .C(n_561), .Y(n_558) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_191), .A2(n_216), .B(n_217), .Y(n_215) );
INVx4_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g502 ( .A(n_192), .Y(n_502) );
AND2x2_ASAP7_75t_L g313 ( .A(n_197), .B(n_258), .Y(n_313) );
OAI322xp33_ASAP7_75t_L g381 ( .A1(n_197), .A2(n_337), .A3(n_382), .B1(n_384), .B2(n_387), .C1(n_389), .C2(n_393), .Y(n_381) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2x1_ASAP7_75t_L g264 ( .A(n_198), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g277 ( .A(n_198), .Y(n_277) );
AND2x2_ASAP7_75t_L g386 ( .A(n_198), .B(n_266), .Y(n_386) );
AND2x2_ASAP7_75t_L g418 ( .A(n_198), .B(n_290), .Y(n_418) );
OR2x2_ASAP7_75t_L g421 ( .A(n_198), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
INVx1_ASAP7_75t_L g251 ( .A(n_199), .Y(n_251) );
AO21x1_ASAP7_75t_L g250 ( .A1(n_201), .A2(n_204), .B(n_251), .Y(n_250) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_204), .A2(n_480), .B(n_490), .Y(n_479) );
INVx3_ASAP7_75t_L g526 ( .A(n_204), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_204), .B(n_538), .Y(n_537) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_204), .A2(n_556), .B(n_563), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_204), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_219), .Y(n_206) );
INVx1_ASAP7_75t_L g434 ( .A(n_207), .Y(n_434) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g239 ( .A(n_208), .B(n_226), .Y(n_239) );
INVx2_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g296 ( .A(n_209), .Y(n_296) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_209), .Y(n_304) );
OR2x2_ASAP7_75t_L g428 ( .A(n_209), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g253 ( .A(n_219), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g293 ( .A(n_219), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g345 ( .A(n_219), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_226), .Y(n_219) );
AND2x2_ASAP7_75t_L g240 ( .A(n_220), .B(n_241), .Y(n_240) );
NOR2xp67_ASAP7_75t_L g300 ( .A(n_220), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g354 ( .A(n_220), .B(n_242), .Y(n_354) );
OR2x2_ASAP7_75t_L g362 ( .A(n_220), .B(n_296), .Y(n_362) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
BUFx2_ASAP7_75t_L g271 ( .A(n_221), .Y(n_271) );
AND2x2_ASAP7_75t_L g281 ( .A(n_221), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g305 ( .A(n_221), .B(n_226), .Y(n_305) );
AND2x2_ASAP7_75t_L g369 ( .A(n_221), .B(n_242), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_226), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_226), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g282 ( .A(n_226), .Y(n_282) );
INVx1_ASAP7_75t_L g287 ( .A(n_226), .Y(n_287) );
AND2x2_ASAP7_75t_L g299 ( .A(n_226), .B(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_226), .Y(n_377) );
INVx1_ASAP7_75t_L g429 ( .A(n_226), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .Y(n_228) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
AND2x2_ASAP7_75t_L g406 ( .A(n_238), .B(n_315), .Y(n_406) );
INVx2_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g333 ( .A(n_240), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g432 ( .A(n_240), .B(n_367), .Y(n_432) );
INVx1_ASAP7_75t_L g254 ( .A(n_241), .Y(n_254) );
AND2x2_ASAP7_75t_L g280 ( .A(n_241), .B(n_274), .Y(n_280) );
BUFx2_ASAP7_75t_L g339 ( .A(n_241), .Y(n_339) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_242), .Y(n_260) );
INVx1_ASAP7_75t_L g270 ( .A(n_242), .Y(n_270) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_245), .Y(n_504) );
INVx2_ASAP7_75t_L g585 ( .A(n_245), .Y(n_585) );
INVx1_ASAP7_75t_L g549 ( .A(n_247), .Y(n_549) );
NOR2xp67_ASAP7_75t_L g408 ( .A(n_248), .B(n_255), .Y(n_408) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI32xp33_ASAP7_75t_L g252 ( .A1(n_249), .A2(n_253), .A3(n_255), .B1(n_257), .B2(n_259), .Y(n_252) );
AND2x2_ASAP7_75t_L g392 ( .A(n_249), .B(n_265), .Y(n_392) );
AND2x2_ASAP7_75t_L g430 ( .A(n_249), .B(n_328), .Y(n_430) );
INVx1_ASAP7_75t_L g310 ( .A(n_250), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_254), .B(n_316), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_255), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_255), .B(n_258), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_255), .B(n_327), .Y(n_409) );
OR2x2_ASAP7_75t_L g423 ( .A(n_255), .B(n_292), .Y(n_423) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g350 ( .A(n_256), .B(n_258), .Y(n_350) );
OR2x2_ASAP7_75t_L g359 ( .A(n_256), .B(n_346), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_258), .B(n_309), .Y(n_331) );
INVx2_ASAP7_75t_L g346 ( .A(n_260), .Y(n_346) );
OR2x2_ASAP7_75t_L g361 ( .A(n_260), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g376 ( .A(n_260), .B(n_377), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_260), .A2(n_353), .B(n_434), .C(n_435), .Y(n_433) );
OAI321xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_267), .A3(n_272), .B1(n_275), .B2(n_279), .C(n_283), .Y(n_261) );
INVx1_ASAP7_75t_L g374 ( .A(n_262), .Y(n_374) );
NAND2x1p5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
AND2x2_ASAP7_75t_L g385 ( .A(n_263), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g337 ( .A(n_265), .Y(n_337) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_266), .B(n_380), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_267), .A2(n_405), .B1(n_407), .B2(n_409), .C(n_410), .Y(n_404) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
AND2x2_ASAP7_75t_L g342 ( .A(n_269), .B(n_316), .Y(n_342) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_270), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g315 ( .A(n_271), .Y(n_315) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_272), .A2(n_313), .B(n_358), .C(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g324 ( .A(n_274), .B(n_281), .Y(n_324) );
BUFx2_ASAP7_75t_L g334 ( .A(n_274), .Y(n_334) );
INVx1_ASAP7_75t_L g349 ( .A(n_274), .Y(n_349) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OR2x2_ASAP7_75t_L g355 ( .A(n_277), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g438 ( .A(n_277), .Y(n_438) );
INVx1_ASAP7_75t_L g431 ( .A(n_278), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AND2x2_ASAP7_75t_L g284 ( .A(n_280), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g388 ( .A(n_280), .B(n_305), .Y(n_388) );
INVx1_ASAP7_75t_L g317 ( .A(n_281), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_288), .B1(n_291), .B2(n_293), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_285), .B(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_L g353 ( .A(n_286), .B(n_354), .Y(n_353) );
BUFx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_SL g316 ( .A(n_287), .B(n_296), .Y(n_316) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g308 ( .A(n_290), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g318 ( .A(n_292), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OAI221xp5_ASAP7_75t_L g412 ( .A1(n_295), .A2(n_413), .B1(n_415), .B2(n_416), .C(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g301 ( .A(n_296), .Y(n_301) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_296), .Y(n_367) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_299), .B(n_418), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_300), .A2(n_305), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_303), .B(n_313), .Y(n_410) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g379 ( .A(n_304), .Y(n_379) );
AND2x2_ASAP7_75t_L g338 ( .A(n_305), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g427 ( .A(n_305), .Y(n_427) );
INVx1_ASAP7_75t_L g343 ( .A(n_308), .Y(n_343) );
INVx1_ASAP7_75t_L g398 ( .A(n_309), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_314), .B1(n_317), .B2(n_318), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_315), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g383 ( .A(n_316), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_316), .B(n_354), .Y(n_420) );
OR2x2_ASAP7_75t_L g393 ( .A(n_317), .B(n_346), .Y(n_393) );
INVx1_ASAP7_75t_L g332 ( .A(n_318), .Y(n_332) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_320), .B(n_371), .Y(n_370) );
NOR3xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_340), .C(n_351), .Y(n_321) );
OAI211xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_325), .B(n_329), .C(n_335), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_324), .A2(n_395), .B1(n_399), .B2(n_402), .C(n_404), .Y(n_394) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AND2x2_ASAP7_75t_L g336 ( .A(n_327), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g390 ( .A(n_327), .B(n_391), .Y(n_390) );
OAI211xp5_ASAP7_75t_L g375 ( .A1(n_328), .A2(n_376), .B(n_378), .C(n_380), .Y(n_375) );
INVx2_ASAP7_75t_L g422 ( .A(n_328), .Y(n_422) );
OAI21xp5_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_332), .B(n_333), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g401 ( .A(n_334), .B(n_354), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
OAI21xp5_ASAP7_75t_SL g340 ( .A1(n_341), .A2(n_343), .B(n_344), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OAI21xp5_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_347), .B(n_350), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_345), .B(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_350), .B(n_437), .Y(n_436) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B(n_357), .Y(n_351) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g378 ( .A(n_354), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND4x1_ASAP7_75t_L g363 ( .A(n_364), .B(n_394), .C(n_411), .D(n_433), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_381), .Y(n_364) );
OAI211xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_370), .B(n_373), .C(n_375), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_369), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_380), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g415 ( .A(n_390), .Y(n_415) );
INVx2_ASAP7_75t_SL g403 ( .A(n_391), .Y(n_403) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g416 ( .A(n_401), .Y(n_416) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NOR2xp33_ASAP7_75t_SL g411 ( .A(n_412), .B(n_419), .Y(n_411) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_421), .B1(n_423), .B2(n_424), .C(n_425), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_430), .B1(n_431), .B2(n_432), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVxp67_ASAP7_75t_L g451 ( .A(n_440), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g452 ( .A(n_444), .Y(n_452) );
BUFx2_ASAP7_75t_L g454 ( .A(n_444), .Y(n_454) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI211xp5_ASAP7_75t_L g449 ( .A1(n_448), .A2(n_450), .B(n_451), .C(n_452), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_453), .B(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_SL g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g759 ( .A(n_460), .Y(n_759) );
INVx1_ASAP7_75t_L g464 ( .A(n_461), .Y(n_464) );
OAI22xp5_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_469), .B1(n_472), .B2(n_756), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OAI22xp5_ASAP7_75t_SL g760 ( .A1(n_468), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_760) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g761 ( .A(n_470), .Y(n_761) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g762 ( .A(n_472), .Y(n_762) );
OR3x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_654), .C(n_719), .Y(n_472) );
NAND4xp25_ASAP7_75t_SL g473 ( .A(n_474), .B(n_595), .C(n_621), .D(n_644), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_527), .B1(n_565), .B2(n_572), .C(n_587), .Y(n_474) );
CKINVDCx14_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_476), .A2(n_588), .B1(n_612), .B2(n_743), .Y(n_742) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_508), .Y(n_476) );
INVx1_ASAP7_75t_SL g648 ( .A(n_477), .Y(n_648) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_492), .Y(n_477) );
OR2x2_ASAP7_75t_L g570 ( .A(n_478), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g590 ( .A(n_478), .B(n_509), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_478), .B(n_517), .Y(n_603) );
AND2x2_ASAP7_75t_L g620 ( .A(n_478), .B(n_492), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_478), .B(n_568), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_478), .B(n_619), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_478), .B(n_508), .Y(n_741) );
AOI211xp5_ASAP7_75t_SL g752 ( .A1(n_478), .A2(n_658), .B(n_753), .C(n_754), .Y(n_752) );
INVx5_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_479), .B(n_509), .Y(n_624) );
AND2x2_ASAP7_75t_L g627 ( .A(n_479), .B(n_510), .Y(n_627) );
OR2x2_ASAP7_75t_L g672 ( .A(n_479), .B(n_509), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_479), .B(n_517), .Y(n_681) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B(n_484), .Y(n_480) );
INVx5_ASAP7_75t_L g498 ( .A(n_485), .Y(n_498) );
INVx5_ASAP7_75t_SL g571 ( .A(n_492), .Y(n_571) );
AND2x2_ASAP7_75t_L g589 ( .A(n_492), .B(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_492), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g675 ( .A(n_492), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g707 ( .A(n_492), .B(n_517), .Y(n_707) );
OR2x2_ASAP7_75t_L g713 ( .A(n_492), .B(n_603), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_492), .B(n_663), .Y(n_722) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_507), .Y(n_492) );
BUFx2_ASAP7_75t_L g544 ( .A(n_495), .Y(n_544) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_498), .A2(n_506), .B(n_521), .C(n_522), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_SL g579 ( .A1(n_498), .A2(n_506), .B(n_580), .C(n_581), .Y(n_579) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B(n_503), .C(n_504), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_501), .A2(n_504), .B(n_535), .C(n_536), .Y(n_534) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_517), .Y(n_508) );
AND2x2_ASAP7_75t_L g604 ( .A(n_509), .B(n_571), .Y(n_604) );
INVx1_ASAP7_75t_SL g617 ( .A(n_509), .Y(n_617) );
OR2x2_ASAP7_75t_L g652 ( .A(n_509), .B(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g658 ( .A(n_509), .B(n_517), .Y(n_658) );
AND2x2_ASAP7_75t_L g716 ( .A(n_509), .B(n_568), .Y(n_716) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_510), .B(n_571), .Y(n_643) );
INVx3_ASAP7_75t_L g568 ( .A(n_517), .Y(n_568) );
OR2x2_ASAP7_75t_L g609 ( .A(n_517), .B(n_571), .Y(n_609) );
AND2x2_ASAP7_75t_L g619 ( .A(n_517), .B(n_617), .Y(n_619) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_517), .Y(n_667) );
AND2x2_ASAP7_75t_L g676 ( .A(n_517), .B(n_590), .Y(n_676) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_525), .Y(n_517) );
OA21x2_ASAP7_75t_L g577 ( .A1(n_526), .A2(n_578), .B(n_586), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_527), .A2(n_693), .B1(n_695), .B2(n_697), .C(n_700), .Y(n_692) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_539), .Y(n_528) );
AND2x2_ASAP7_75t_L g666 ( .A(n_529), .B(n_647), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_529), .B(n_725), .Y(n_729) );
OR2x2_ASAP7_75t_L g750 ( .A(n_529), .B(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_529), .B(n_755), .Y(n_754) );
BUFx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx5_ASAP7_75t_L g597 ( .A(n_530), .Y(n_597) );
AND2x2_ASAP7_75t_L g674 ( .A(n_530), .B(n_541), .Y(n_674) );
AND2x2_ASAP7_75t_L g735 ( .A(n_530), .B(n_614), .Y(n_735) );
AND2x2_ASAP7_75t_L g748 ( .A(n_530), .B(n_568), .Y(n_748) );
OR2x6_ASAP7_75t_L g530 ( .A(n_531), .B(n_537), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_553), .Y(n_539) );
AND2x4_ASAP7_75t_L g575 ( .A(n_540), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g593 ( .A(n_540), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g600 ( .A(n_540), .Y(n_600) );
AND2x2_ASAP7_75t_L g669 ( .A(n_540), .B(n_647), .Y(n_669) );
AND2x2_ASAP7_75t_L g679 ( .A(n_540), .B(n_597), .Y(n_679) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_540), .Y(n_687) );
AND2x2_ASAP7_75t_L g699 ( .A(n_540), .B(n_577), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_540), .B(n_631), .Y(n_703) );
AND2x2_ASAP7_75t_L g740 ( .A(n_540), .B(n_735), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_540), .B(n_614), .Y(n_751) );
OR2x2_ASAP7_75t_L g753 ( .A(n_540), .B(n_689), .Y(n_753) );
INVx5_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g639 ( .A(n_541), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g649 ( .A(n_541), .B(n_594), .Y(n_649) );
AND2x2_ASAP7_75t_L g661 ( .A(n_541), .B(n_577), .Y(n_661) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_541), .Y(n_691) );
AND2x4_ASAP7_75t_L g725 ( .A(n_541), .B(n_576), .Y(n_725) );
OR2x6_ASAP7_75t_L g541 ( .A(n_542), .B(n_550), .Y(n_541) );
AOI21xp5_ASAP7_75t_SL g542 ( .A1(n_543), .A2(n_545), .B(n_549), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
BUFx2_ASAP7_75t_L g574 ( .A(n_553), .Y(n_574) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g614 ( .A(n_554), .Y(n_614) );
AND2x2_ASAP7_75t_L g647 ( .A(n_554), .B(n_577), .Y(n_647) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g594 ( .A(n_555), .B(n_577), .Y(n_594) );
BUFx2_ASAP7_75t_L g640 ( .A(n_555), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_562), .Y(n_556) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_567), .B(n_648), .Y(n_727) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_568), .B(n_590), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_568), .B(n_571), .Y(n_629) );
AND2x2_ASAP7_75t_L g684 ( .A(n_568), .B(n_620), .Y(n_684) );
AOI221xp5_ASAP7_75t_SL g621 ( .A1(n_569), .A2(n_622), .B1(n_630), .B2(n_632), .C(n_636), .Y(n_621) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g616 ( .A(n_570), .B(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g657 ( .A(n_570), .B(n_658), .Y(n_657) );
OAI321xp33_ASAP7_75t_L g664 ( .A1(n_570), .A2(n_623), .A3(n_665), .B1(n_667), .B2(n_668), .C(n_670), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_571), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_574), .B(n_725), .Y(n_743) );
AND2x2_ASAP7_75t_L g630 ( .A(n_575), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_575), .B(n_634), .Y(n_633) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_576), .Y(n_606) );
AND2x2_ASAP7_75t_L g613 ( .A(n_576), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_576), .B(n_688), .Y(n_718) );
INVx1_ASAP7_75t_L g755 ( .A(n_576), .Y(n_755) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_591), .B(n_592), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
A2O1A1Ixp33_ASAP7_75t_L g747 ( .A1(n_589), .A2(n_699), .B(n_748), .C(n_749), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_590), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_590), .B(n_628), .Y(n_694) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g637 ( .A(n_594), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_594), .B(n_597), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_594), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_594), .B(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_598), .B1(n_610), .B2(n_615), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g611 ( .A(n_597), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g634 ( .A(n_597), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g646 ( .A(n_597), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_597), .B(n_640), .Y(n_682) );
OR2x2_ASAP7_75t_L g689 ( .A(n_597), .B(n_614), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_597), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g739 ( .A(n_597), .B(n_725), .Y(n_739) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .B1(n_605), .B2(n_607), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g645 ( .A(n_600), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
OAI22xp33_ASAP7_75t_L g685 ( .A1(n_603), .A2(n_618), .B1(n_686), .B2(n_690), .Y(n_685) );
INVx1_ASAP7_75t_L g733 ( .A(n_604), .Y(n_733) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_608), .A2(n_645), .B1(n_648), .B2(n_649), .C(n_650), .Y(n_644) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g623 ( .A(n_609), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_613), .B(n_679), .Y(n_711) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_614), .Y(n_631) );
INVx1_ASAP7_75t_L g635 ( .A(n_614), .Y(n_635) );
NAND2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx1_ASAP7_75t_L g653 ( .A(n_620), .Y(n_653) );
AND2x2_ASAP7_75t_L g662 ( .A(n_620), .B(n_663), .Y(n_662) );
NAND2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx2_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
AND2x4_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
AND2x2_ASAP7_75t_L g706 ( .A(n_627), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_630), .A2(n_656), .B1(n_659), .B2(n_662), .C(n_664), .Y(n_655) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_634), .B(n_691), .Y(n_690) );
AOI21xp33_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_638), .B(n_641), .Y(n_636) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
CKINVDCx16_ASAP7_75t_R g738 ( .A(n_641), .Y(n_738) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
OR2x2_ASAP7_75t_L g680 ( .A(n_643), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g701 ( .A(n_646), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_646), .B(n_706), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_649), .B(n_671), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_655), .B(n_673), .C(n_692), .D(n_705), .Y(n_654) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g663 ( .A(n_658), .Y(n_663) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g696 ( .A(n_667), .B(n_672), .Y(n_696) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B(n_677), .C(n_685), .Y(n_673) );
AOI211xp5_ASAP7_75t_L g744 ( .A1(n_675), .A2(n_717), .B(n_745), .C(n_752), .Y(n_744) );
INVx1_ASAP7_75t_SL g704 ( .A(n_676), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B1(n_682), .B2(n_683), .Y(n_677) );
INVx1_ASAP7_75t_L g708 ( .A(n_682), .Y(n_708) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_688), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_688), .B(n_699), .Y(n_732) );
INVx2_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g709 ( .A(n_699), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B(n_704), .Y(n_700) );
INVxp33_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI322xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_708), .A3(n_709), .B1(n_710), .B2(n_712), .C1(n_714), .C2(n_717), .Y(n_705) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND3xp33_ASAP7_75t_SL g719 ( .A(n_720), .B(n_737), .C(n_744), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_723), .B1(n_726), .B2(n_728), .C(n_730), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g736 ( .A(n_725), .Y(n_736) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI22xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_739), .B1(n_740), .B2(n_741), .C(n_742), .Y(n_737) );
NAND2xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVxp67_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g763 ( .A(n_757), .Y(n_763) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
endmodule