module fake_ibex_1793_n_849 (n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_849);

input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_849;

wire n_151;
wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_418;
wire n_256;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_840;
wire n_561;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_285;
wire n_379;
wire n_247;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_159;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_559;
wire n_425;

BUFx3_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_82),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_68),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_94),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_2),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_30),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_55),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_49),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_27),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_24),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_2),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVxp33_ASAP7_75t_SL g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_43),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_118),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_22),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_61),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_40),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_97),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_16),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_93),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_34),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_34),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_92),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_48),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_91),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_L g195 ( 
.A(n_59),
.B(n_26),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_71),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_13),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_12),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_150),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_19),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_13),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_37),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_105),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_21),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_32),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_19),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_41),
.Y(n_211)
);

BUFx2_ASAP7_75t_SL g212 ( 
.A(n_60),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_26),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_14),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_37),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_10),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_67),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_86),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_120),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_1),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_22),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_95),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_8),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_30),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_39),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_45),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_138),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_63),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_101),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_116),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_50),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_62),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_14),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_122),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_18),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_69),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_73),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_36),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_149),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_6),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_126),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_123),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_11),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_58),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_66),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_64),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_112),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_96),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_100),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_117),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_152),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_0),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_160),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_3),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_152),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_152),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_178),
.B(n_3),
.Y(n_259)
);

OA22x2_ASAP7_75t_SL g260 ( 
.A1(n_185),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_161),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_151),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_186),
.B(n_4),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_155),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_152),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_154),
.Y(n_267)
);

AND2x6_ASAP7_75t_L g268 ( 
.A(n_151),
.B(n_42),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_5),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_204),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_155),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_173),
.B(n_7),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_164),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_159),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_182),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_204),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_182),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_231),
.B(n_7),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_171),
.Y(n_279)
);

AND2x2_ASAP7_75t_SL g280 ( 
.A(n_162),
.B(n_44),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_190),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_189),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_204),
.Y(n_283)
);

AND2x4_ASAP7_75t_L g284 ( 
.A(n_206),
.B(n_8),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_205),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_211),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_190),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_211),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_228),
.B(n_9),
.Y(n_289)
);

OA21x2_ASAP7_75t_L g290 ( 
.A1(n_192),
.A2(n_81),
.B(n_148),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_209),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_192),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_196),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_196),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_215),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_228),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_173),
.B(n_9),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_172),
.B(n_10),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_158),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_215),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_213),
.Y(n_301)
);

BUFx8_ASAP7_75t_L g302 ( 
.A(n_221),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_216),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_221),
.B(n_11),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_217),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_218),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_161),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_230),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_223),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_230),
.Y(n_310)
);

INVx5_ASAP7_75t_L g311 ( 
.A(n_212),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_163),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_158),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_235),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_165),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_225),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_227),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_235),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_166),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_167),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_240),
.B(n_20),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_242),
.B(n_20),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_169),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_300),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_300),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_255),
.B(n_187),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_304),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_253),
.Y(n_329)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_268),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_300),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_280),
.A2(n_184),
.B1(n_174),
.B2(n_246),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_261),
.A2(n_176),
.B1(n_184),
.B2(n_174),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_284),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_279),
.Y(n_339)
);

NOR3xp33_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_208),
.C(n_188),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_265),
.B(n_176),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_261),
.B(n_157),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_310),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_254),
.A2(n_197),
.B1(n_198),
.B2(n_202),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_311),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_288),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_288),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_267),
.B(n_175),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_288),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_279),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_254),
.A2(n_210),
.B1(n_222),
.B2(n_226),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_296),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_280),
.A2(n_248),
.B1(n_170),
.B2(n_246),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_296),
.Y(n_357)
);

NOR3xp33_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_237),
.C(n_180),
.Y(n_358)
);

OR2x6_ASAP7_75t_L g359 ( 
.A(n_272),
.B(n_195),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_296),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_296),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_312),
.B(n_177),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_291),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_L g364 ( 
.A1(n_321),
.A2(n_245),
.B1(n_185),
.B2(n_248),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_291),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_297),
.B(n_232),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g369 ( 
.A(n_284),
.B(n_181),
.Y(n_369)
);

AND3x2_ASAP7_75t_L g370 ( 
.A(n_260),
.B(n_191),
.C(n_183),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_297),
.B(n_232),
.Y(n_371)
);

AND2x2_ASAP7_75t_SL g372 ( 
.A(n_289),
.B(n_193),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_302),
.B(n_233),
.Y(n_373)
);

OR2x6_ASAP7_75t_L g374 ( 
.A(n_259),
.B(n_170),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_289),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_262),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_303),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_257),
.Y(n_378)
);

AND3x2_ASAP7_75t_L g379 ( 
.A(n_259),
.B(n_200),
.C(n_194),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_289),
.Y(n_380)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_256),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_315),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_262),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_315),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_317),
.B(n_203),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_257),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_258),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_268),
.A2(n_244),
.B1(n_224),
.B2(n_251),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_258),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_274),
.B(n_241),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_320),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_320),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_258),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_258),
.Y(n_395)
);

NOR2x1p5_ASAP7_75t_L g396 ( 
.A(n_299),
.B(n_245),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_258),
.Y(n_397)
);

OR2x6_ASAP7_75t_L g398 ( 
.A(n_263),
.B(n_298),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_269),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_273),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_282),
.B(n_153),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_270),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_320),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_285),
.B(n_156),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_R g405 ( 
.A(n_299),
.B(n_168),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_372),
.A2(n_278),
.B1(n_322),
.B2(n_319),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_286),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_286),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_334),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_339),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_401),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_342),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_353),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_301),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_383),
.Y(n_415)
);

AOI221xp5_ASAP7_75t_L g416 ( 
.A1(n_364),
.A2(n_305),
.B1(n_316),
.B2(n_309),
.C(n_306),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_383),
.B(n_368),
.Y(n_417)
);

BUFx6f_ASAP7_75t_SL g418 ( 
.A(n_374),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_368),
.B(n_319),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_341),
.B(n_313),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_371),
.B(n_268),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_363),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_371),
.B(n_268),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_367),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_369),
.A2(n_320),
.B1(n_323),
.B2(n_308),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_369),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_342),
.B(n_264),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_377),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_L g429 ( 
.A(n_358),
.B(n_290),
.C(n_323),
.Y(n_429)
);

BUFx5_ASAP7_75t_L g430 ( 
.A(n_369),
.Y(n_430)
);

BUFx5_ASAP7_75t_L g431 ( 
.A(n_369),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_398),
.A2(n_323),
.B1(n_295),
.B2(n_294),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_400),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_398),
.A2(n_323),
.B1(n_295),
.B2(n_294),
.Y(n_434)
);

AND2x4_ASAP7_75t_SL g435 ( 
.A(n_374),
.B(n_264),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_400),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_330),
.B(n_179),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_365),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_327),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_376),
.B(n_199),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_365),
.B(n_271),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_328),
.B(n_207),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_324),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_328),
.B(n_219),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_336),
.B(n_239),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_333),
.B(n_336),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_340),
.A2(n_293),
.B1(n_292),
.B2(n_271),
.Y(n_449)
);

BUFx8_ASAP7_75t_L g450 ( 
.A(n_396),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_338),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_338),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_405),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_356),
.A2(n_335),
.B1(n_354),
.B2(n_346),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_359),
.B(n_275),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_338),
.A2(n_293),
.B1(n_292),
.B2(n_275),
.Y(n_456)
);

BUFx5_ASAP7_75t_L g457 ( 
.A(n_324),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_374),
.B(n_337),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_375),
.B(n_250),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_375),
.B(n_252),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_374),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_331),
.Y(n_462)
);

OAI22xp33_ASAP7_75t_L g463 ( 
.A1(n_359),
.A2(n_277),
.B1(n_287),
.B2(n_281),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_375),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_380),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_331),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_380),
.A2(n_290),
.B(n_287),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_359),
.B(n_351),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_385),
.B(n_277),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_373),
.B(n_214),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_362),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_404),
.B(n_220),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_389),
.B(n_229),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_347),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_347),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_379),
.B(n_234),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_414),
.B(n_359),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_438),
.B(n_370),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_406),
.A2(n_247),
.B1(n_236),
.B2(n_238),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_21),
.Y(n_480)
);

AO21x1_ASAP7_75t_L g481 ( 
.A1(n_467),
.A2(n_384),
.B(n_366),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_421),
.A2(n_392),
.B(n_386),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_423),
.A2(n_392),
.B(n_386),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_406),
.B(n_23),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_439),
.A2(n_403),
.B(n_393),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_426),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_448),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_411),
.B(n_23),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_443),
.Y(n_489)
);

NOR3xp33_ASAP7_75t_SL g490 ( 
.A(n_454),
.B(n_24),
.C(n_25),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_451),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_430),
.B(n_345),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_407),
.A2(n_326),
.B(n_325),
.Y(n_493)
);

AO22x1_ASAP7_75t_L g494 ( 
.A1(n_450),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_412),
.B(n_28),
.Y(n_495)
);

AO21x1_ASAP7_75t_L g496 ( 
.A1(n_463),
.A2(n_469),
.B(n_473),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_459),
.A2(n_460),
.B(n_452),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_464),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_462),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_427),
.B(n_29),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_430),
.B(n_348),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_461),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_465),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_419),
.B(n_31),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_442),
.A2(n_344),
.B(n_332),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_471),
.B(n_415),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_444),
.A2(n_343),
.B(n_332),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_409),
.Y(n_508)
);

OAI21xp33_ASAP7_75t_L g509 ( 
.A1(n_416),
.A2(n_349),
.B(n_360),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_458),
.A2(n_266),
.B1(n_361),
.B2(n_349),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_410),
.Y(n_511)
);

OA21x2_ASAP7_75t_L g512 ( 
.A1(n_456),
.A2(n_350),
.B(n_352),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_453),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_420),
.B(n_31),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_462),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_413),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_435),
.B(n_33),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_417),
.A2(n_355),
.B1(n_357),
.B2(n_266),
.Y(n_518)
);

OA21x2_ASAP7_75t_L g519 ( 
.A1(n_456),
.A2(n_357),
.B(n_355),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_418),
.A2(n_266),
.B1(n_270),
.B2(n_276),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_462),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_468),
.A2(n_266),
.B1(n_270),
.B2(n_276),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_408),
.B(n_35),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_R g524 ( 
.A(n_418),
.B(n_36),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_466),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_422),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_424),
.Y(n_527)
);

OR2x6_ASAP7_75t_SL g528 ( 
.A(n_450),
.B(n_38),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_455),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_428),
.Y(n_530)
);

CKINVDCx10_ASAP7_75t_R g531 ( 
.A(n_476),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_466),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_L g533 ( 
.A(n_430),
.B(n_283),
.Y(n_533)
);

O2A1O1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_470),
.A2(n_397),
.B(n_395),
.C(n_394),
.Y(n_534)
);

AO32x1_ASAP7_75t_L g535 ( 
.A1(n_433),
.A2(n_378),
.A3(n_390),
.B1(n_388),
.B2(n_387),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_449),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_445),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_432),
.B(n_434),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_440),
.Y(n_539)
);

INVx5_ASAP7_75t_L g540 ( 
.A(n_436),
.Y(n_540)
);

CKINVDCx10_ASAP7_75t_R g541 ( 
.A(n_449),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_437),
.A2(n_329),
.B(n_402),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_472),
.B(n_46),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_506),
.B(n_431),
.Y(n_544)
);

A2O1A1Ixp33_ASAP7_75t_L g545 ( 
.A1(n_490),
.A2(n_475),
.B(n_474),
.C(n_425),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_511),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_536),
.B(n_431),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_486),
.Y(n_548)
);

OAI21x1_ASAP7_75t_SL g549 ( 
.A1(n_496),
.A2(n_431),
.B(n_457),
.Y(n_549)
);

OA21x2_ASAP7_75t_L g550 ( 
.A1(n_481),
.A2(n_447),
.B(n_446),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_516),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_539),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_526),
.B(n_457),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_527),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_482),
.A2(n_457),
.B(n_51),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_483),
.A2(n_457),
.B(n_52),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_477),
.B(n_47),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_502),
.Y(n_558)
);

NAND3x1_ASAP7_75t_L g559 ( 
.A(n_528),
.B(n_53),
.C(n_54),
.Y(n_559)
);

NAND3x1_ASAP7_75t_L g560 ( 
.A(n_524),
.B(n_56),
.C(n_57),
.Y(n_560)
);

INVx8_ASAP7_75t_L g561 ( 
.A(n_540),
.Y(n_561)
);

AOI221x1_ASAP7_75t_L g562 ( 
.A1(n_479),
.A2(n_65),
.B1(n_72),
.B2(n_74),
.C(n_75),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_505),
.A2(n_77),
.B(n_78),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_507),
.A2(n_79),
.B(n_80),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_485),
.A2(n_83),
.B(n_84),
.Y(n_565)
);

OAI21x1_ASAP7_75t_SL g566 ( 
.A1(n_484),
.A2(n_85),
.B(n_87),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_530),
.B(n_88),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_500),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_480),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_487),
.A2(n_488),
.B(n_538),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_529),
.B(n_495),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_491),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_478),
.B(n_99),
.Y(n_573)
);

OAI22x1_ASAP7_75t_L g574 ( 
.A1(n_514),
.A2(n_102),
.B1(n_103),
.B2(n_108),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_517),
.B(n_110),
.Y(n_575)
);

CKINVDCx11_ASAP7_75t_R g576 ( 
.A(n_513),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_504),
.A2(n_113),
.B(n_115),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_537),
.B(n_503),
.Y(n_578)
);

AOI221x1_ASAP7_75t_L g579 ( 
.A1(n_522),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.C(n_129),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_541),
.B(n_141),
.Y(n_580)
);

A2O1A1Ixp33_ASAP7_75t_L g581 ( 
.A1(n_523),
.A2(n_144),
.B(n_145),
.C(n_146),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_541),
.B(n_489),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_510),
.B(n_498),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_543),
.B(n_515),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_493),
.A2(n_512),
.B(n_519),
.Y(n_585)
);

NOR2xp67_ASAP7_75t_L g586 ( 
.A(n_515),
.B(n_521),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_492),
.A2(n_501),
.B(n_535),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_521),
.Y(n_588)
);

NOR2xp67_ASAP7_75t_L g589 ( 
.A(n_525),
.B(n_518),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_535),
.A2(n_533),
.B(n_534),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_494),
.B(n_509),
.Y(n_591)
);

AO31x2_ASAP7_75t_L g592 ( 
.A1(n_520),
.A2(n_499),
.A3(n_532),
.B(n_531),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_532),
.B(n_531),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_506),
.B(n_414),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_486),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_477),
.B(n_374),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_542),
.A2(n_467),
.B(n_481),
.Y(n_597)
);

BUFx12f_ASAP7_75t_L g598 ( 
.A(n_513),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_524),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_490),
.B(n_514),
.C(n_429),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_508),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_539),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_508),
.Y(n_603)
);

OAI21xp33_ASAP7_75t_L g604 ( 
.A1(n_490),
.A2(n_414),
.B(n_514),
.Y(n_604)
);

OAI21x1_ASAP7_75t_L g605 ( 
.A1(n_542),
.A2(n_467),
.B(n_481),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_506),
.B(n_438),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_524),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_508),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_506),
.B(n_414),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_536),
.A2(n_454),
.B1(n_458),
.B2(n_418),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_506),
.B(n_438),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_506),
.A2(n_372),
.B1(n_335),
.B2(n_406),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_513),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_513),
.Y(n_614)
);

AO22x2_ASAP7_75t_L g615 ( 
.A1(n_479),
.A2(n_335),
.B1(n_454),
.B2(n_458),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_497),
.A2(n_429),
.B(n_467),
.Y(n_616)
);

OAI21x1_ASAP7_75t_L g617 ( 
.A1(n_542),
.A2(n_467),
.B(n_481),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_594),
.B(n_609),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_596),
.B(n_606),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_598),
.Y(n_620)
);

OA21x2_ASAP7_75t_L g621 ( 
.A1(n_585),
.A2(n_617),
.B(n_605),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_554),
.B(n_601),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_L g623 ( 
.A1(n_570),
.A2(n_600),
.B(n_545),
.Y(n_623)
);

AO21x2_ASAP7_75t_L g624 ( 
.A1(n_549),
.A2(n_590),
.B(n_597),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_608),
.B(n_568),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_551),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_558),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_561),
.B(n_593),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_604),
.A2(n_577),
.B(n_591),
.C(n_584),
.Y(n_629)
);

INVx4_ASAP7_75t_SL g630 ( 
.A(n_592),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_603),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_615),
.B(n_610),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_615),
.A2(n_583),
.B1(n_577),
.B2(n_569),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_572),
.B(n_544),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_561),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_611),
.Y(n_636)
);

AO31x2_ASAP7_75t_L g637 ( 
.A1(n_562),
.A2(n_579),
.A3(n_574),
.B(n_581),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_561),
.B(n_602),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_552),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_582),
.B(n_613),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_578),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_576),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_614),
.Y(n_643)
);

AO31x2_ASAP7_75t_L g644 ( 
.A1(n_555),
.A2(n_556),
.A3(n_563),
.B(n_564),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_580),
.B(n_575),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_547),
.B(n_553),
.Y(n_646)
);

CKINVDCx11_ASAP7_75t_R g647 ( 
.A(n_595),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_548),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_550),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_588),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_589),
.A2(n_567),
.B(n_557),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_599),
.Y(n_652)
);

INVx8_ASAP7_75t_L g653 ( 
.A(n_548),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_571),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_559),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_607),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_573),
.B(n_586),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_560),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_576),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_576),
.Y(n_660)
);

AO21x2_ASAP7_75t_L g661 ( 
.A1(n_585),
.A2(n_549),
.B(n_616),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_606),
.Y(n_662)
);

BUFx8_ASAP7_75t_L g663 ( 
.A(n_598),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_606),
.B(n_611),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_606),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_546),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_606),
.B(n_611),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_615),
.A2(n_612),
.B1(n_610),
.B2(n_536),
.Y(n_668)
);

AO21x2_ASAP7_75t_L g669 ( 
.A1(n_585),
.A2(n_549),
.B(n_616),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_606),
.B(n_611),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_546),
.Y(n_671)
);

AO31x2_ASAP7_75t_L g672 ( 
.A1(n_587),
.A2(n_481),
.A3(n_496),
.B(n_590),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_606),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_546),
.Y(n_674)
);

OAI22xp33_ASAP7_75t_L g675 ( 
.A1(n_612),
.A2(n_335),
.B1(n_356),
.B2(n_374),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_606),
.B(n_611),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_615),
.A2(n_612),
.B1(n_610),
.B2(n_536),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_606),
.B(n_611),
.Y(n_678)
);

OAI21x1_ASAP7_75t_SL g679 ( 
.A1(n_577),
.A2(n_565),
.B(n_566),
.Y(n_679)
);

INVx6_ASAP7_75t_L g680 ( 
.A(n_598),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_561),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_634),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_649),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_635),
.Y(n_684)
);

NAND2x1_ASAP7_75t_L g685 ( 
.A(n_679),
.B(n_658),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_SL g686 ( 
.A(n_659),
.B(n_663),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_622),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_665),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_653),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_622),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_630),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_658),
.B(n_630),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_632),
.B(n_668),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_676),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_632),
.B(n_668),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_677),
.A2(n_675),
.B1(n_619),
.B2(n_655),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_677),
.B(n_670),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_621),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_676),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_625),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_673),
.B(n_618),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_647),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_618),
.B(n_664),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_673),
.B(n_667),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_638),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_625),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_626),
.B(n_666),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_631),
.B(n_671),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_678),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_648),
.B(n_674),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_641),
.B(n_654),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_653),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_SL g713 ( 
.A1(n_633),
.A2(n_629),
.B(n_651),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_636),
.B(n_623),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_662),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_627),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_645),
.A2(n_640),
.B1(n_633),
.B2(n_639),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_661),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_648),
.B(n_681),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_681),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_669),
.B(n_638),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_646),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_653),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_638),
.B(n_672),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_672),
.B(n_628),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_650),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_643),
.Y(n_727)
);

AO21x2_ASAP7_75t_L g728 ( 
.A1(n_624),
.A2(n_651),
.B(n_657),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_672),
.B(n_628),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_628),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_650),
.B(n_637),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_714),
.B(n_637),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_702),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_693),
.B(n_642),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_703),
.B(n_620),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_709),
.Y(n_736)
);

NOR2x1_ASAP7_75t_L g737 ( 
.A(n_685),
.B(n_705),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_683),
.Y(n_738)
);

AND2x4_ASAP7_75t_SL g739 ( 
.A(n_692),
.B(n_689),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_698),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_701),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_692),
.B(n_644),
.Y(n_742)
);

NAND2x1_ASAP7_75t_L g743 ( 
.A(n_692),
.B(n_691),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_724),
.B(n_644),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_701),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_691),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_716),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_704),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_704),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_711),
.B(n_642),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_731),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_693),
.B(n_656),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_687),
.B(n_680),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_707),
.B(n_680),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_731),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_695),
.B(n_660),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_707),
.B(n_652),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_708),
.B(n_682),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_695),
.B(n_663),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_708),
.B(n_652),
.Y(n_760)
);

OAI33xp33_ASAP7_75t_L g761 ( 
.A1(n_688),
.A2(n_715),
.A3(n_697),
.B1(n_690),
.B2(n_700),
.B3(n_706),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_697),
.B(n_725),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_694),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_720),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_696),
.A2(n_717),
.B1(n_722),
.B2(n_700),
.Y(n_765)
);

OAI22xp33_ASAP7_75t_L g766 ( 
.A1(n_702),
.A2(n_686),
.B1(n_689),
.B2(n_706),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_684),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_744),
.B(n_728),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_740),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_744),
.B(n_728),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_762),
.B(n_725),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_747),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_742),
.B(n_721),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_738),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_762),
.B(n_729),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_732),
.B(n_718),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_758),
.B(n_690),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_741),
.B(n_729),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_751),
.B(n_721),
.Y(n_779)
);

OAI222xp33_ASAP7_75t_L g780 ( 
.A1(n_759),
.A2(n_730),
.B1(n_722),
.B2(n_699),
.C1(n_712),
.C2(n_723),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_776),
.B(n_748),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_773),
.B(n_742),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_772),
.B(n_749),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_777),
.B(n_745),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_780),
.B(n_759),
.Y(n_785)
);

NOR2x1_ASAP7_75t_L g786 ( 
.A(n_778),
.B(n_766),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_769),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_773),
.B(n_742),
.Y(n_788)
);

AND2x4_ASAP7_75t_SL g789 ( 
.A(n_773),
.B(n_746),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_768),
.B(n_755),
.Y(n_790)
);

HB1xp67_ASAP7_75t_SL g791 ( 
.A(n_773),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_776),
.B(n_758),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_768),
.B(n_755),
.Y(n_793)
);

INVxp67_ASAP7_75t_SL g794 ( 
.A(n_774),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_770),
.B(n_742),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_779),
.A2(n_765),
.B1(n_735),
.B2(n_761),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_781),
.B(n_771),
.Y(n_797)
);

NOR2x1p5_ASAP7_75t_L g798 ( 
.A(n_791),
.B(n_743),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_781),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_785),
.B(n_750),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_794),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_795),
.B(n_790),
.Y(n_802)
);

OAI211xp5_ASAP7_75t_L g803 ( 
.A1(n_785),
.A2(n_734),
.B(n_767),
.C(n_713),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_792),
.B(n_775),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_787),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_782),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_782),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_784),
.B(n_775),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_797),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_799),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_801),
.Y(n_811)
);

OAI211xp5_ASAP7_75t_L g812 ( 
.A1(n_803),
.A2(n_796),
.B(n_733),
.C(n_736),
.Y(n_812)
);

OAI21xp33_ASAP7_75t_SL g813 ( 
.A1(n_798),
.A2(n_786),
.B(n_737),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_807),
.B(n_806),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_800),
.A2(n_788),
.B1(n_782),
.B2(n_793),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_801),
.Y(n_816)
);

OAI322xp33_ASAP7_75t_L g817 ( 
.A1(n_800),
.A2(n_734),
.A3(n_783),
.B1(n_756),
.B2(n_778),
.C1(n_752),
.C2(n_713),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_805),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_808),
.Y(n_819)
);

OAI211xp5_ASAP7_75t_L g820 ( 
.A1(n_812),
.A2(n_756),
.B(n_765),
.C(n_806),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_814),
.B(n_806),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_815),
.A2(n_804),
.B1(n_752),
.B2(n_789),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_818),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_L g824 ( 
.A(n_822),
.B(n_818),
.Y(n_824)
);

NOR2xp67_ASAP7_75t_L g825 ( 
.A(n_820),
.B(n_813),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_SL g826 ( 
.A(n_822),
.B(n_817),
.Y(n_826)
);

NOR4xp25_ASAP7_75t_L g827 ( 
.A(n_824),
.B(n_812),
.C(n_816),
.D(n_811),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_825),
.Y(n_828)
);

NOR2xp67_ASAP7_75t_L g829 ( 
.A(n_828),
.B(n_823),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_827),
.Y(n_830)
);

NAND4xp25_ASAP7_75t_SL g831 ( 
.A(n_830),
.B(n_826),
.C(n_821),
.D(n_819),
.Y(n_831)
);

NOR3x2_ASAP7_75t_L g832 ( 
.A(n_829),
.B(n_684),
.C(n_727),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_832),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_831),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_833),
.Y(n_835)
);

OAI22x1_ASAP7_75t_L g836 ( 
.A1(n_834),
.A2(n_754),
.B1(n_753),
.B2(n_809),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_833),
.Y(n_837)
);

AO22x2_ASAP7_75t_L g838 ( 
.A1(n_837),
.A2(n_836),
.B1(n_757),
.B2(n_760),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_835),
.B(n_810),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_835),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_837),
.Y(n_841)
);

AO22x1_ASAP7_75t_L g842 ( 
.A1(n_841),
.A2(n_840),
.B1(n_839),
.B2(n_838),
.Y(n_842)
);

XNOR2xp5_ASAP7_75t_L g843 ( 
.A(n_841),
.B(n_720),
.Y(n_843)
);

AOI221xp5_ASAP7_75t_L g844 ( 
.A1(n_842),
.A2(n_719),
.B1(n_726),
.B2(n_763),
.C(n_710),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_SL g845 ( 
.A1(n_843),
.A2(n_739),
.B(n_726),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_844),
.B(n_719),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_845),
.B(n_710),
.Y(n_847)
);

OA21x2_ASAP7_75t_L g848 ( 
.A1(n_846),
.A2(n_847),
.B(n_805),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_848),
.A2(n_764),
.B1(n_802),
.B2(n_788),
.Y(n_849)
);


endmodule