module fake_netlist_6_3914_n_458 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_458);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_458;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_148;
wire n_208;
wire n_161;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_392;
wire n_442;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_443;
wire n_246;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_360;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_397;
wire n_155;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_381;
wire n_236;
wire n_172;
wire n_270;
wire n_239;
wire n_414;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_417;
wire n_446;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_293;
wire n_334;
wire n_370;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_456;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_406;
wire n_204;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_292;
wire n_164;
wire n_307;
wire n_433;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_136;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_418;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_328;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVxp67_ASAP7_75t_SL g127 ( 
.A(n_33),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_17),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_41),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_4),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_29),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

NOR2xp67_ASAP7_75t_L g134 ( 
.A(n_9),
.B(n_53),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_22),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_52),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_2),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_50),
.Y(n_140)
);

INVxp33_ASAP7_75t_SL g141 ( 
.A(n_99),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g142 ( 
.A(n_70),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_13),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_85),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_56),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_43),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_44),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_30),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_6),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_18),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_11),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_77),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_19),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_121),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_32),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_34),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_62),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_91),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_24),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_49),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_54),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_27),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_12),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_78),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_81),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_92),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_23),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_90),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_66),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_83),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_93),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_82),
.Y(n_185)
);

INVxp33_ASAP7_75t_SL g186 ( 
.A(n_89),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_123),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_68),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_61),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_16),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_58),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_71),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_1),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_57),
.Y(n_196)
);

INVxp67_ASAP7_75t_SL g197 ( 
.A(n_42),
.Y(n_197)
);

INVxp33_ASAP7_75t_SL g198 ( 
.A(n_21),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_3),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_139),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_0),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_0),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_1),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_132),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_3),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_133),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_136),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_138),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_134),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_143),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_144),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_130),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_140),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_149),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

AND2x4_ASAP7_75t_L g225 ( 
.A(n_169),
.B(n_181),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_153),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_155),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_128),
.B(n_162),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_156),
.A2(n_7),
.B(n_8),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_158),
.Y(n_234)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

NAND2x1p5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_220),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

AND2x4_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_127),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_188),
.Y(n_247)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_179),
.C(n_162),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_200),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_159),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_141),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_160),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_127),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_216),
.B(n_167),
.Y(n_257)
);

AND2x4_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_142),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_215),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_202),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_210),
.B(n_161),
.Y(n_261)
);

NAND2x1p5_ASAP7_75t_L g262 ( 
.A(n_203),
.B(n_166),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_214),
.B(n_168),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_218),
.B(n_170),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_211),
.B(n_186),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g270 ( 
.A(n_223),
.B(n_142),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_217),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_219),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_242),
.A2(n_233),
.B1(n_211),
.B2(n_206),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_237),
.Y(n_274)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_235),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

AND2x6_ASAP7_75t_SL g277 ( 
.A(n_254),
.B(n_204),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_257),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_239),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_244),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_259),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_259),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_247),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_249),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

AND2x4_ASAP7_75t_L g293 ( 
.A(n_242),
.B(n_180),
.Y(n_293)
);

AND3x1_ASAP7_75t_SL g294 ( 
.A(n_265),
.B(n_221),
.C(n_172),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_247),
.A2(n_198),
.B1(n_135),
.B2(n_178),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_256),
.B(n_253),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_197),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_258),
.B(n_270),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_251),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_255),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_253),
.B(n_226),
.Y(n_304)
);

BUFx4f_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_248),
.A2(n_177),
.B1(n_175),
.B2(n_148),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

BUFx12f_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_267),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_276),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_280),
.Y(n_312)
);

AOI221xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_248),
.B1(n_221),
.B2(n_263),
.C(n_266),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_308),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_288),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_262),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

NOR3xp33_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_261),
.C(n_128),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_285),
.Y(n_320)
);

HAxp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_8),
.CON(n_321),
.SN(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_299),
.B(n_137),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_253),
.Y(n_323)
);

AND2x6_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_174),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_274),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_276),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_309),
.Y(n_327)
);

OR2x6_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_230),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_L g329 ( 
.A(n_272),
.B(n_145),
.C(n_146),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_309),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_284),
.B(n_236),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_303),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_292),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_310),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_301),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_279),
.Y(n_337)
);

AND3x1_ASAP7_75t_SL g338 ( 
.A(n_277),
.B(n_189),
.C(n_182),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_303),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_281),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_298),
.Y(n_341)
);

OAI33xp33_ASAP7_75t_L g342 ( 
.A1(n_278),
.A2(n_250),
.A3(n_236),
.B1(n_234),
.B2(n_231),
.B3(n_224),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_273),
.A2(n_197),
.B1(n_176),
.B2(n_183),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_282),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_303),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

INVx3_ASAP7_75t_SL g348 ( 
.A(n_316),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_313),
.A2(n_233),
.B1(n_253),
.B2(n_304),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_327),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_290),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_330),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_305),
.Y(n_353)
);

NAND2x1p5_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_286),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_343),
.A2(n_195),
.B1(n_192),
.B2(n_190),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_320),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_330),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_315),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_319),
.A2(n_324),
.B1(n_334),
.B2(n_332),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_341),
.Y(n_361)
);

BUFx8_ASAP7_75t_L g362 ( 
.A(n_314),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_321),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_342),
.A2(n_229),
.B1(n_295),
.B2(n_250),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_332),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_324),
.A2(n_271),
.B1(n_291),
.B2(n_287),
.Y(n_367)
);

OA21x2_ASAP7_75t_L g368 ( 
.A1(n_323),
.A2(n_271),
.B(n_163),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_338),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_317),
.B(n_264),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_346),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_325),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_347),
.Y(n_373)
);

AOI221xp5_ASAP7_75t_L g374 ( 
.A1(n_363),
.A2(n_322),
.B1(n_336),
.B2(n_329),
.C(n_311),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_371),
.A2(n_346),
.B(n_333),
.Y(n_375)
);

AO221x2_ASAP7_75t_L g376 ( 
.A1(n_363),
.A2(n_9),
.B1(n_331),
.B2(n_345),
.C(n_344),
.Y(n_376)
);

OAI211xp5_ASAP7_75t_L g377 ( 
.A1(n_361),
.A2(n_337),
.B(n_340),
.C(n_325),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_371),
.A2(n_339),
.B1(n_328),
.B2(n_311),
.Y(n_378)
);

AO21x2_ASAP7_75t_L g379 ( 
.A1(n_350),
.A2(n_324),
.B(n_340),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_349),
.A2(n_339),
.B(n_307),
.Y(n_380)
);

AOI221xp5_ASAP7_75t_L g381 ( 
.A1(n_355),
.A2(n_318),
.B1(n_164),
.B2(n_196),
.C(n_165),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_349),
.A2(n_318),
.B1(n_287),
.B2(n_286),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_355),
.A2(n_365),
.B1(n_366),
.B2(n_358),
.Y(n_383)
);

CKINVDCx6p67_ASAP7_75t_R g384 ( 
.A(n_348),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_352),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_359),
.A2(n_291),
.B1(n_286),
.B2(n_307),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_353),
.A2(n_324),
.B1(n_291),
.B2(n_275),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_372),
.A2(n_275),
.B1(n_14),
.B2(n_15),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_348),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_373),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_376),
.A2(n_369),
.B1(n_362),
.B2(n_370),
.Y(n_393)
);

OAI222xp33_ASAP7_75t_L g394 ( 
.A1(n_383),
.A2(n_367),
.B1(n_364),
.B2(n_372),
.C1(n_351),
.C2(n_360),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_386),
.A2(n_367),
.B1(n_354),
.B2(n_351),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_385),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_384),
.Y(n_397)
);

OAI221xp5_ASAP7_75t_L g398 ( 
.A1(n_374),
.A2(n_364),
.B1(n_368),
.B2(n_362),
.C(n_20),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_10),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_389),
.B(n_381),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_379),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_25),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_382),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_403)
);

AOI221xp5_ASAP7_75t_L g404 ( 
.A1(n_390),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.C(n_38),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_379),
.A2(n_39),
.B1(n_40),
.B2(n_45),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_400),
.A2(n_388),
.B1(n_377),
.B2(n_375),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_392),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_401),
.Y(n_408)
);

AOI33xp33_ASAP7_75t_L g409 ( 
.A1(n_393),
.A2(n_46),
.A3(n_47),
.B1(n_48),
.B2(n_51),
.B3(n_55),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_396),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_397),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_391),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_395),
.Y(n_413)
);

A2O1A1Ixp33_ASAP7_75t_L g414 ( 
.A1(n_398),
.A2(n_60),
.B(n_63),
.C(n_64),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_399),
.Y(n_415)
);

OAI211xp5_ASAP7_75t_L g416 ( 
.A1(n_404),
.A2(n_405),
.B(n_402),
.C(n_403),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_392),
.Y(n_418)
);

OAI31xp33_ASAP7_75t_L g419 ( 
.A1(n_400),
.A2(n_65),
.A3(n_67),
.B(n_72),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_73),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_74),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_415),
.B(n_75),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_76),
.Y(n_423)
);

OAI33xp33_ASAP7_75t_L g424 ( 
.A1(n_413),
.A2(n_79),
.A3(n_80),
.B1(n_84),
.B2(n_87),
.B3(n_88),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_418),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_408),
.Y(n_426)
);

NOR2x1_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_94),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_95),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_100),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_411),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_101),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_102),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_409),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_425),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_426),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_409),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_428),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_422),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_422),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_431),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_429),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_SL g442 ( 
.A(n_436),
.B(n_433),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_434),
.Y(n_443)
);

AOI322xp5_ASAP7_75t_L g444 ( 
.A1(n_442),
.A2(n_438),
.A3(n_432),
.B1(n_439),
.B2(n_427),
.C1(n_435),
.C2(n_414),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_443),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_441),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_444),
.A2(n_414),
.B(n_423),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_447),
.A2(n_437),
.B1(n_424),
.B2(n_419),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_446),
.Y(n_449)
);

NAND4xp25_ASAP7_75t_L g450 ( 
.A(n_448),
.B(n_421),
.C(n_420),
.D(n_435),
.Y(n_450)
);

AO22x2_ASAP7_75t_L g451 ( 
.A1(n_449),
.A2(n_416),
.B1(n_106),
.B2(n_107),
.Y(n_451)
);

AND3x1_ASAP7_75t_L g452 ( 
.A(n_450),
.B(n_112),
.C(n_113),
.Y(n_452)
);

OA22x2_ASAP7_75t_L g453 ( 
.A1(n_452),
.A2(n_451),
.B1(n_116),
.B2(n_119),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_452),
.B(n_114),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_454),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_455),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_456),
.B(n_453),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_457),
.A2(n_124),
.B(n_120),
.Y(n_458)
);


endmodule