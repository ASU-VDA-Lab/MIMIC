module real_jpeg_30266_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g159 ( 
.A(n_0),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_0),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g333 ( 
.A(n_0),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_0),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_0),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_1),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_1),
.B(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_1),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_1),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_1),
.B(n_90),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g462 ( 
.A(n_1),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_1),
.B(n_489),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_2),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_2),
.B(n_327),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_2),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_2),
.B(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_2),
.B(n_498),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_2),
.B(n_503),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_2),
.B(n_508),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_3),
.B(n_533),
.Y(n_532)
);

CKINVDCx11_ASAP7_75t_R g537 ( 
.A(n_3),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_5),
.Y(n_295)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_6),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_6),
.Y(n_193)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_6),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_7),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_7),
.B(n_45),
.Y(n_44)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_7),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_7),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_7),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_7),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_7),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_8),
.B(n_37),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_8),
.B(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_8),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_8),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_8),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_8),
.B(n_485),
.Y(n_484)
);

AND2x2_ASAP7_75t_SL g495 ( 
.A(n_8),
.B(n_248),
.Y(n_495)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_9),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_9),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_9),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_10),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_11),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_11),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_SL g264 ( 
.A(n_11),
.B(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_11),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_11),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_11),
.B(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_11),
.B(n_437),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_11),
.B(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_12),
.Y(n_146)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_12),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_13),
.B(n_62),
.Y(n_61)
);

AND2x6_ASAP7_75t_SL g71 ( 
.A(n_13),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_13),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_13),
.B(n_141),
.Y(n_140)
);

NAND2x1_ASAP7_75t_L g199 ( 
.A(n_13),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g270 ( 
.A(n_13),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_13),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_13),
.B(n_360),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_14),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_15),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_16),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_16),
.B(n_68),
.Y(n_67)
);

NAND2x1_ASAP7_75t_L g89 ( 
.A(n_16),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_16),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_16),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_16),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_16),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_17),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_17),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_17),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_17),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_17),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_17),
.B(n_333),
.Y(n_332)
);

OAI311xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_167),
.A3(n_532),
.B1(n_534),
.C1(n_536),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_20),
.B(n_532),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_165),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_103),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_22),
.B(n_103),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_50),
.C(n_65),
.Y(n_23)
);

XNOR2x1_ASAP7_75t_L g104 ( 
.A(n_24),
.B(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_39),
.B1(n_48),
.B2(n_49),
.Y(n_24)
);

INVxp67_ASAP7_75t_SL g48 ( 
.A(n_25),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_R g25 ( 
.A(n_26),
.B(n_31),
.C(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_26),
.A2(n_31),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_26),
.Y(n_132)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_31),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_31),
.B(n_199),
.C(n_202),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_31),
.A2(n_133),
.B1(n_202),
.B2(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_32),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_33),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_33),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_33),
.Y(n_310)
);

XOR2x2_ASAP7_75t_L g130 ( 
.A(n_34),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_38),
.Y(n_189)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

MAJx2_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_47),
.C(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_43),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_43),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_43),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_44),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_44),
.A2(n_47),
.B1(n_163),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_44),
.A2(n_47),
.B1(n_204),
.B2(n_253),
.Y(n_252)
);

INVx8_ASAP7_75t_L g314 ( 
.A(n_45),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_47),
.B(n_156),
.C(n_163),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_47),
.B(n_198),
.C(n_204),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2x1_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_65),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_56),
.C(n_61),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_R g108 ( 
.A1(n_52),
.A2(n_56),
.B1(n_57),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_52),
.B(n_120),
.C(n_125),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_52),
.B(n_291),
.C(n_297),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_52),
.B(n_291),
.Y(n_303)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_55),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_57),
.B1(n_67),
.B2(n_70),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_92),
.C(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_56),
.B(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_56),
.B(n_143),
.C(n_337),
.Y(n_363)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_58),
.Y(n_307)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_108),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_82),
.B1(n_83),
.B2(n_91),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_67),
.A2(n_70),
.B1(n_232),
.B2(n_366),
.Y(n_365)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_70),
.B(n_138),
.C(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_75),
.Y(n_205)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_75),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_93),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_111),
.C(n_114),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_88),
.B(n_240),
.C(n_246),
.Y(n_239)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2x1_ASAP7_75t_L g379 ( 
.A(n_89),
.B(n_247),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.C(n_129),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_104),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_119),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_107),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_120),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_110),
.B(n_119),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_114),
.B1(n_115),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_111),
.A2(n_138),
.B1(n_365),
.B2(n_367),
.Y(n_364)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_112),
.Y(n_499)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_123),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_124),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_126),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_157),
.C(n_160),
.Y(n_156)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_126),
.B(n_160),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_126),
.B(n_244),
.Y(n_430)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_128),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_129),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_531)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.C(n_155),
.Y(n_129)
);

XNOR2x1_ASAP7_75t_SL g215 ( 
.A(n_130),
.B(n_155),
.Y(n_215)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_135),
.B(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.C(n_152),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_136),
.B(n_139),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_147),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_140),
.A2(n_147),
.B1(n_148),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_144),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_143),
.A2(n_144),
.B1(n_337),
.B2(n_340),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_146),
.Y(n_434)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_152),
.Y(n_223)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_156),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_191),
.Y(n_194)
);

XOR2x2_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_196),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g236 ( 
.A(n_157),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_157),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_157),
.A2(n_436),
.B1(n_438),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_159),
.Y(n_245)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_167),
.B(n_535),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_256),
.B(n_527),
.Y(n_167)
);

NAND2x1_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_216),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_170),
.A2(n_529),
.B(n_530),
.Y(n_528)
);

AOI21x1_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_174),
.B(n_177),
.Y(n_170)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_177),
.B(n_531),
.Y(n_530)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_210),
.C(n_213),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_179),
.B(n_255),
.Y(n_254)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_197),
.C(n_206),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_186),
.C(n_195),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_182),
.B(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_186),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_190),
.B(n_194),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_191),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_191),
.B(n_284),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_191),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_192),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_193),
.Y(n_464)
);

INVx6_ASAP7_75t_L g487 ( 
.A(n_193),
.Y(n_487)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_194),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_194),
.A2(n_321),
.B1(n_440),
.B2(n_441),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_195),
.B(n_405),
.Y(n_404)
);

XNOR2x1_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_207),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_198),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_201),
.Y(n_299)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_203),
.Y(n_328)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_214),
.Y(n_255)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_254),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_217),
.B(n_254),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.C(n_225),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_219),
.B(n_222),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_225),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_239),
.C(n_250),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_226),
.A2(n_227),
.B1(n_400),
.B2(n_401),
.Y(n_399)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.C(n_236),
.Y(n_227)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_228),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_231),
.B(n_236),
.Y(n_384)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_232),
.Y(n_366)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_239),
.A2(n_250),
.B1(n_251),
.B2(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_239),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_240),
.B(n_379),
.Y(n_378)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.C(n_244),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_241),
.B(n_243),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_244),
.B(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_419),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_388),
.B1(n_413),
.B2(n_418),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_368),
.B(n_385),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_341),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_260),
.B(n_341),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_301),
.C(n_318),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_261),
.B(n_319),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_281),
.B2(n_300),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_262),
.B(n_282),
.C(n_290),
.Y(n_350)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g348 ( 
.A(n_264),
.B(n_270),
.C(n_275),
.Y(n_348)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_275),
.B2(n_276),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_289),
.B2(n_290),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_284),
.A2(n_285),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_288),
.Y(n_466)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_296),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_296),
.B(n_459),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_297),
.B(n_303),
.Y(n_302)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_301),
.B(n_425),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.C(n_315),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_302),
.B(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_304),
.B(n_315),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_308),
.C(n_311),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_305),
.B(n_474),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_309),
.B(n_312),
.Y(n_474)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_310),
.Y(n_456)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_329),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_320),
.B(n_330),
.C(n_335),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.C(n_325),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_322),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.Y(n_440)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.Y(n_329)
);

OA21x2_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B(n_334),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_332),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_334),
.B(n_348),
.Y(n_347)
);

MAJx2_ASAP7_75t_L g376 ( 
.A(n_334),
.B(n_345),
.C(n_348),
.Y(n_376)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_337),
.Y(n_340)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_349),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

MAJx2_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_344),
.C(n_349),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_352),
.C(n_364),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_364),
.Y(n_351)
);

XNOR2x2_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_362),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_359),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_359),
.C(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_363),
.Y(n_381)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_365),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

AOI21x1_ASAP7_75t_L g385 ( 
.A1(n_369),
.A2(n_386),
.B(n_387),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_373),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_391),
.C(n_392),
.Y(n_390)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_374),
.Y(n_386)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_382),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_375),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_378),
.C(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_380),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_380),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_382),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_408),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_394),
.Y(n_389)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_398),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_396),
.B(n_399),
.C(n_403),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_403),
.B1(n_404),
.B2(n_407),
.Y(n_398)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_399),
.Y(n_407)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_408),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_409),
.Y(n_415)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_410),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

NAND3xp33_ASAP7_75t_L g419 ( 
.A(n_413),
.B(n_420),
.C(n_422),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_442),
.B(n_526),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_426),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_424),
.B(n_426),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_429),
.C(n_439),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_427),
.B(n_524),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_429),
.B(n_439),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.C(n_435),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_430),
.A2(n_431),
.B1(n_432),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_434),
.Y(n_460)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_434),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_435),
.B(n_478),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_438),
.Y(n_435)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_436),
.Y(n_469)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_440),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_520),
.B(n_525),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_444),
.A2(n_480),
.B(n_519),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_470),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_445),
.B(n_470),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_461),
.C(n_467),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_446),
.A2(n_447),
.B1(n_515),
.B2(n_517),
.Y(n_514)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_458),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_450),
.B1(n_454),
.B2(n_457),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_449),
.B(n_457),
.C(n_458),
.Y(n_472)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_454),
.Y(n_457)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_461),
.A2(n_467),
.B1(n_468),
.B2(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_461),
.Y(n_516)
);

NAND2x1_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_465),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_465),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_477),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_473),
.B1(n_475),
.B2(n_476),
.Y(n_471)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_472),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_473),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_473),
.B(n_475),
.C(n_522),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_477),
.Y(n_522)
);

AOI21x1_ASAP7_75t_SL g480 ( 
.A1(n_481),
.A2(n_512),
.B(n_518),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_482),
.A2(n_500),
.B(n_511),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_491),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_483),
.B(n_491),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_488),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_488),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_484),
.B(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

BUFx4f_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_492),
.B(n_495),
.C(n_496),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_494),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_506),
.B(n_510),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_505),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_505),
.Y(n_510)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_514),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_SL g518 ( 
.A(n_513),
.B(n_514),
.Y(n_518)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_515),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_523),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_523),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_532),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_538),
.Y(n_536)
);


endmodule