module fake_jpeg_17049_n_195 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_195);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_26),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_33),
.Y(n_55)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_38),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_25),
.B1(n_17),
.B2(n_16),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_30),
.B1(n_27),
.B2(n_16),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_16),
.B1(n_17),
.B2(n_33),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_43),
.B1(n_31),
.B2(n_22),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_22),
.Y(n_66)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_16),
.B1(n_27),
.B2(n_30),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_60),
.A2(n_59),
.B1(n_80),
.B2(n_21),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_62),
.B(n_67),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_20),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_59),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_34),
.B1(n_18),
.B2(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_72),
.A2(n_84),
.B1(n_45),
.B2(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_2),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_19),
.B(n_26),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_20),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_79),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_26),
.B(n_19),
.C(n_36),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_32),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_83),
.Y(n_105)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_19),
.B1(n_21),
.B2(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_40),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_98),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_87),
.A2(n_102),
.B1(n_103),
.B2(n_77),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_82),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_15),
.C(n_13),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_96),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_106),
.B(n_74),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_45),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_71),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_63),
.B(n_71),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_103),
.B(n_86),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_81),
.B1(n_64),
.B2(n_83),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_85),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_89),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_97),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_41),
.B(n_36),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_98),
.B(n_41),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_3),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_61),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_127),
.B(n_103),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_123),
.B1(n_110),
.B2(n_118),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_106),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_132),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_92),
.B(n_103),
.C(n_104),
.D(n_95),
.Y(n_131)
);

XOR2x2_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_141),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_101),
.C(n_40),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_70),
.C(n_29),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_135),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_70),
.C(n_103),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_29),
.C(n_41),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_110),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_3),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_142),
.B(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_142),
.B(n_129),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_116),
.B(n_115),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_158),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_155),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_143),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_144),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_159),
.C(n_117),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_138),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_166),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_137),
.C(n_131),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_157),
.C(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_169),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_154),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_168),
.A2(n_147),
.B1(n_148),
.B2(n_157),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_147),
.A2(n_113),
.B(n_4),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_153),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_3),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_162),
.Y(n_178)
);

OAI21x1_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_9),
.B(n_12),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_176),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_6),
.C(n_10),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_182),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_161),
.B1(n_165),
.B2(n_167),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_181),
.B1(n_176),
.B2(n_174),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_6),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_187),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_179),
.A2(n_172),
.B(n_177),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_188),
.B(n_178),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_12),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_177),
.B(n_5),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_189),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_188),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_191),
.A2(n_13),
.B(n_4),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_190),
.C(n_5),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_193),
.Y(n_195)
);


endmodule