module fake_aes_6756_n_809 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_96, n_39, n_809);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_96;
input n_39;
output n_809;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_808;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_223;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_40), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_6), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_77), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_87), .Y(n_101) );
CKINVDCx14_ASAP7_75t_R g102 ( .A(n_5), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_10), .Y(n_103) );
INVxp33_ASAP7_75t_L g104 ( .A(n_38), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_34), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_26), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_96), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_10), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_71), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_45), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_84), .Y(n_111) );
INVx2_ASAP7_75t_SL g112 ( .A(n_37), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_80), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_26), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_51), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_3), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_33), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_20), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_86), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_23), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_89), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_15), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_58), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_61), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_85), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_29), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_42), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_46), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_25), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_70), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_41), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_44), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_48), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_35), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_14), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_19), .Y(n_137) );
BUFx10_ASAP7_75t_L g138 ( .A(n_93), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_56), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_90), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_91), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_137), .Y(n_142) );
BUFx12f_ASAP7_75t_L g143 ( .A(n_138), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_104), .B(n_0), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_132), .Y(n_145) );
INVxp67_ASAP7_75t_L g146 ( .A(n_105), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_105), .B(n_0), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_137), .B(n_1), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_138), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_137), .B(n_1), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_132), .Y(n_151) );
BUFx2_ASAP7_75t_L g152 ( .A(n_102), .Y(n_152) );
INVx5_ASAP7_75t_L g153 ( .A(n_132), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_138), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_138), .B(n_2), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_113), .B(n_2), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_113), .B(n_39), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_112), .B(n_3), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_116), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_126), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_112), .B(n_4), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_132), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_116), .B(n_4), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_117), .B(n_5), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g165 ( .A1(n_146), .A2(n_98), .B1(n_140), .B2(n_119), .Y(n_165) );
OA22x2_ASAP7_75t_L g166 ( .A1(n_146), .A2(n_117), .B1(n_114), .B2(n_136), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_149), .B(n_126), .Y(n_167) );
OAI22x1_ASAP7_75t_L g168 ( .A1(n_146), .A2(n_114), .B1(n_130), .B2(n_135), .Y(n_168) );
AO22x2_ASAP7_75t_L g169 ( .A1(n_156), .A2(n_131), .B1(n_101), .B2(n_8), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_155), .A2(n_99), .B1(n_127), .B2(n_103), .Y(n_170) );
OAI22xp33_ASAP7_75t_L g171 ( .A1(n_163), .A2(n_106), .B1(n_108), .B2(n_118), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_155), .A2(n_120), .B1(n_122), .B2(n_131), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_152), .B(n_101), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_155), .A2(n_141), .B1(n_139), .B2(n_134), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_148), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_153), .Y(n_176) );
OA22x2_ASAP7_75t_L g177 ( .A1(n_159), .A2(n_133), .B1(n_129), .B2(n_128), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_152), .B(n_100), .Y(n_178) );
OA22x2_ASAP7_75t_L g179 ( .A1(n_159), .A2(n_107), .B1(n_109), .B2(n_110), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_153), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
OAI22xp33_ASAP7_75t_R g183 ( .A1(n_158), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_155), .A2(n_125), .B1(n_124), .B2(n_123), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_152), .A2(n_121), .B1(n_115), .B2(n_111), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_152), .B(n_159), .Y(n_186) );
OAI22xp33_ASAP7_75t_SL g187 ( .A1(n_164), .A2(n_7), .B1(n_9), .B2(n_11), .Y(n_187) );
OAI22xp33_ASAP7_75t_L g188 ( .A1(n_163), .A2(n_132), .B1(n_11), .B2(n_12), .Y(n_188) );
AO22x2_ASAP7_75t_L g189 ( .A1(n_156), .A2(n_9), .B1(n_12), .B2(n_13), .Y(n_189) );
OAI22xp33_ASAP7_75t_SL g190 ( .A1(n_164), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_190) );
INVx8_ASAP7_75t_L g191 ( .A(n_143), .Y(n_191) );
OAI22xp33_ASAP7_75t_L g192 ( .A1(n_163), .A2(n_132), .B1(n_17), .B2(n_18), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
OAI22xp33_ASAP7_75t_SL g194 ( .A1(n_164), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_148), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_153), .Y(n_196) );
OAI22xp33_ASAP7_75t_R g197 ( .A1(n_158), .A2(n_16), .B1(n_19), .B2(n_20), .Y(n_197) );
OR2x2_ASAP7_75t_L g198 ( .A(n_147), .B(n_21), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_147), .A2(n_21), .B1(n_22), .B2(n_23), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_153), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_148), .Y(n_201) );
BUFx10_ASAP7_75t_L g202 ( .A(n_156), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_149), .A2(n_22), .B1(n_24), .B2(n_25), .Y(n_203) );
AO22x2_ASAP7_75t_L g204 ( .A1(n_156), .A2(n_24), .B1(n_27), .B2(n_28), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_148), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_148), .Y(n_206) );
AO22x2_ASAP7_75t_L g207 ( .A1(n_156), .A2(n_27), .B1(n_28), .B2(n_29), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_149), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_153), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_147), .B(n_143), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_165), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_191), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_201), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_201), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_201), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_186), .B(n_147), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_206), .Y(n_217) );
XNOR2x2_ASAP7_75t_L g218 ( .A(n_169), .B(n_189), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_206), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_191), .B(n_210), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_173), .B(n_143), .Y(n_221) );
INVxp67_ASAP7_75t_L g222 ( .A(n_178), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_191), .B(n_149), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_206), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_175), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_185), .B(n_143), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_180), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_195), .Y(n_228) );
NAND2x1p5_ASAP7_75t_L g229 ( .A(n_205), .B(n_156), .Y(n_229) );
NOR2xp33_ASAP7_75t_SL g230 ( .A(n_202), .B(n_143), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_202), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_202), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_198), .B(n_149), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_170), .Y(n_234) );
NAND2x1p5_ASAP7_75t_L g235 ( .A(n_199), .B(n_156), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_167), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_167), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_189), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_189), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_204), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_204), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_174), .Y(n_242) );
NAND2xp33_ASAP7_75t_SL g243 ( .A(n_168), .B(n_149), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_204), .Y(n_244) );
XNOR2xp5_ASAP7_75t_L g245 ( .A(n_177), .B(n_149), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_184), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_172), .B(n_154), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_207), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_207), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_171), .B(n_154), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_171), .A2(n_156), .B(n_157), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_176), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_207), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_169), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_169), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_177), .B(n_154), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_179), .B(n_154), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_168), .B(n_154), .Y(n_258) );
CKINVDCx14_ASAP7_75t_R g259 ( .A(n_203), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_166), .B(n_154), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_179), .B(n_154), .Y(n_261) );
INVxp67_ASAP7_75t_SL g262 ( .A(n_188), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_188), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_166), .B(n_148), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_187), .B(n_144), .Y(n_265) );
AOI21x1_ASAP7_75t_L g266 ( .A1(n_176), .A2(n_157), .B(n_160), .Y(n_266) );
INVx1_ASAP7_75t_SL g267 ( .A(n_208), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_192), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_183), .Y(n_269) );
INVxp33_ASAP7_75t_L g270 ( .A(n_197), .Y(n_270) );
XOR2x2_ASAP7_75t_L g271 ( .A(n_190), .B(n_144), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_181), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_219), .Y(n_273) );
INVx4_ASAP7_75t_L g274 ( .A(n_212), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_219), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_219), .Y(n_276) );
AND2x4_ASAP7_75t_SL g277 ( .A(n_212), .B(n_148), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_212), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_252), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_252), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_221), .B(n_150), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_221), .B(n_150), .Y(n_282) );
INVx6_ASAP7_75t_L g283 ( .A(n_212), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_252), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_216), .B(n_150), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_229), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_216), .B(n_150), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_213), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_235), .B(n_150), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_213), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_214), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_231), .Y(n_292) );
OAI21xp5_ASAP7_75t_L g293 ( .A1(n_251), .A2(n_157), .B(n_161), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_235), .B(n_247), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_236), .B(n_160), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_231), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_235), .B(n_150), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_236), .B(n_160), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_237), .B(n_192), .Y(n_299) );
INVx2_ASAP7_75t_SL g300 ( .A(n_232), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_237), .B(n_144), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_265), .B(n_150), .Y(n_302) );
OAI21xp5_ASAP7_75t_L g303 ( .A1(n_251), .A2(n_158), .B(n_161), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_232), .Y(n_304) );
INVx2_ASAP7_75t_SL g305 ( .A(n_229), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_247), .B(n_150), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_225), .B(n_194), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_222), .B(n_161), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_225), .B(n_142), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_227), .B(n_142), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_229), .Y(n_311) );
AND2x2_ASAP7_75t_SL g312 ( .A(n_238), .B(n_142), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_214), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_215), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_233), .B(n_181), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_238), .B(n_30), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_256), .B(n_209), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_218), .Y(n_318) );
INVx4_ASAP7_75t_L g319 ( .A(n_233), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_267), .B(n_209), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_215), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_227), .B(n_200), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_211), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_294), .B(n_267), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_286), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_294), .B(n_264), .Y(n_326) );
AND2x6_ASAP7_75t_L g327 ( .A(n_278), .B(n_286), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_290), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_274), .B(n_239), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_290), .Y(n_330) );
OR2x6_ASAP7_75t_L g331 ( .A(n_274), .B(n_239), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_290), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_274), .B(n_228), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_294), .B(n_264), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_302), .B(n_228), .Y(n_335) );
AND2x2_ASAP7_75t_SL g336 ( .A(n_318), .B(n_254), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_294), .B(n_262), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_286), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_289), .B(n_240), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_274), .Y(n_340) );
NOR2xp33_ASAP7_75t_SL g341 ( .A(n_274), .B(n_230), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_308), .B(n_234), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_302), .B(n_263), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_319), .B(n_270), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_319), .B(n_271), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_289), .B(n_240), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_289), .B(n_241), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_290), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_274), .B(n_217), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_286), .Y(n_350) );
OR2x4_ASAP7_75t_L g351 ( .A(n_286), .B(n_226), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_274), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_278), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_302), .B(n_263), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_306), .B(n_268), .Y(n_355) );
OR2x6_ASAP7_75t_SL g356 ( .A(n_345), .B(n_254), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_327), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_325), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_328), .Y(n_359) );
BUFx12f_ASAP7_75t_L g360 ( .A(n_327), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_325), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_327), .Y(n_362) );
BUFx12f_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_327), .Y(n_365) );
BUFx12f_ASAP7_75t_SL g366 ( .A(n_329), .Y(n_366) );
INVx3_ASAP7_75t_SL g367 ( .A(n_352), .Y(n_367) );
BUFx5_ASAP7_75t_L g368 ( .A(n_327), .Y(n_368) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_327), .Y(n_369) );
INVx5_ASAP7_75t_SL g370 ( .A(n_329), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_330), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_327), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_330), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_337), .B(n_289), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_332), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_332), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_348), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_348), .Y(n_378) );
INVx5_ASAP7_75t_L g379 ( .A(n_327), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g380 ( .A(n_338), .B(n_286), .Y(n_380) );
INVx4_ASAP7_75t_L g381 ( .A(n_340), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_338), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_340), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_339), .Y(n_384) );
BUFx12f_ASAP7_75t_L g385 ( .A(n_360), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_364), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_360), .Y(n_387) );
AOI22xp5_ASAP7_75t_SL g388 ( .A1(n_365), .A2(n_269), .B1(n_246), .B2(n_259), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_367), .A2(n_345), .B1(n_351), .B2(n_318), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_364), .Y(n_390) );
CKINVDCx6p67_ASAP7_75t_R g391 ( .A(n_367), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_366), .A2(n_342), .B1(n_243), .B2(n_344), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_364), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_360), .Y(n_394) );
OAI21xp5_ASAP7_75t_SL g395 ( .A1(n_357), .A2(n_245), .B(n_297), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_364), .Y(n_396) );
INVx4_ASAP7_75t_SL g397 ( .A(n_360), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_359), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_367), .Y(n_399) );
BUFx2_ASAP7_75t_L g400 ( .A(n_366), .Y(n_400) );
INVx5_ASAP7_75t_L g401 ( .A(n_363), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_366), .A2(n_344), .B1(n_318), .B2(n_271), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_366), .A2(n_218), .B1(n_337), .B2(n_336), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_371), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_359), .Y(n_405) );
BUFx12f_ASAP7_75t_L g406 ( .A(n_363), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_371), .Y(n_407) );
CKINVDCx11_ASAP7_75t_R g408 ( .A(n_367), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_384), .A2(n_337), .B1(n_336), .B2(n_245), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_384), .A2(n_336), .B1(n_297), .B2(n_324), .Y(n_410) );
INVx6_ASAP7_75t_L g411 ( .A(n_363), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_384), .B(n_307), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_379), .Y(n_413) );
INVx5_ASAP7_75t_L g414 ( .A(n_363), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g415 ( .A1(n_383), .A2(n_299), .B(n_343), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_367), .A2(n_297), .B1(n_324), .B2(n_346), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_371), .B(n_339), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_371), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_374), .A2(n_242), .B1(n_308), .B2(n_333), .Y(n_419) );
INVx6_ASAP7_75t_SL g420 ( .A(n_379), .Y(n_420) );
INVx5_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_373), .Y(n_422) );
BUFx2_ASAP7_75t_R g423 ( .A(n_356), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_356), .A2(n_351), .B1(n_341), .B2(n_340), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_370), .A2(n_341), .B1(n_340), .B2(n_353), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_375), .Y(n_426) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_370), .A2(n_353), .B1(n_316), .B2(n_241), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_389), .A2(n_374), .B1(n_370), .B2(n_334), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_423), .A2(n_351), .B1(n_370), .B2(n_356), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_407), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g431 ( .A1(n_401), .A2(n_351), .B1(n_356), .B2(n_379), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_386), .B(n_375), .Y(n_432) );
AOI211xp5_ASAP7_75t_L g433 ( .A1(n_424), .A2(n_257), .B(n_260), .C(n_308), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_386), .B(n_375), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_398), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_425), .B(n_379), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_405), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_403), .A2(n_374), .B1(n_370), .B2(n_334), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_401), .Y(n_439) );
INVx11_ASAP7_75t_L g440 ( .A(n_385), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_407), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_408), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_402), .A2(n_374), .B1(n_370), .B2(n_334), .Y(n_443) );
AOI222xp33_ASAP7_75t_L g444 ( .A1(n_409), .A2(n_244), .B1(n_253), .B2(n_249), .C1(n_248), .C2(n_297), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_416), .A2(n_370), .B1(n_379), .B2(n_357), .Y(n_445) );
OAI21xp5_ASAP7_75t_SL g446 ( .A1(n_400), .A2(n_357), .B(n_258), .Y(n_446) );
BUFx4f_ASAP7_75t_SL g447 ( .A(n_399), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_422), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_417), .B(n_373), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_408), .A2(n_370), .B1(n_326), .B2(n_333), .Y(n_450) );
OAI22xp33_ASAP7_75t_L g451 ( .A1(n_401), .A2(n_379), .B1(n_381), .B2(n_365), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_390), .Y(n_452) );
BUFx4f_ASAP7_75t_SL g453 ( .A(n_399), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_410), .A2(n_379), .B1(n_329), .B2(n_331), .Y(n_454) );
AOI22xp33_ASAP7_75t_SL g455 ( .A1(n_400), .A2(n_365), .B1(n_379), .B2(n_368), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_392), .A2(n_326), .B1(n_333), .B2(n_339), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_390), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_385), .A2(n_326), .B1(n_333), .B2(n_346), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_426), .Y(n_459) );
BUFx6f_ASAP7_75t_SL g460 ( .A(n_413), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_395), .A2(n_305), .B1(n_311), .B2(n_319), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_406), .A2(n_347), .B1(n_346), .B2(n_253), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_406), .A2(n_347), .B1(n_248), .B2(n_244), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_426), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_417), .A2(n_347), .B1(n_249), .B2(n_258), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g466 ( .A1(n_411), .A2(n_365), .B1(n_379), .B2(n_368), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_420), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_421), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_393), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_396), .B(n_375), .Y(n_470) );
OAI21xp5_ASAP7_75t_SL g471 ( .A1(n_387), .A2(n_362), .B(n_303), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_391), .A2(n_381), .B1(n_303), .B2(n_331), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_391), .A2(n_381), .B1(n_303), .B2(n_331), .Y(n_473) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_421), .Y(n_474) );
OAI222xp33_ASAP7_75t_L g475 ( .A1(n_388), .A2(n_381), .B1(n_373), .B2(n_378), .C1(n_377), .C2(n_376), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_412), .B(n_376), .Y(n_476) );
AOI211xp5_ASAP7_75t_L g477 ( .A1(n_415), .A2(n_260), .B(n_307), .C(n_323), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_397), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_396), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_419), .A2(n_381), .B1(n_331), .B2(n_329), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_427), .A2(n_331), .B1(n_329), .B2(n_377), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_404), .Y(n_482) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_421), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_404), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_418), .B(n_376), .Y(n_485) );
OAI222xp33_ASAP7_75t_L g486 ( .A1(n_401), .A2(n_381), .B1(n_377), .B2(n_378), .C1(n_255), .C2(n_362), .Y(n_486) );
INVx5_ASAP7_75t_SL g487 ( .A(n_397), .Y(n_487) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_401), .A2(n_331), .B1(n_329), .B2(n_372), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_411), .A2(n_305), .B1(n_311), .B2(n_319), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_411), .A2(n_316), .B1(n_268), .B2(n_343), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_418), .B(n_378), .Y(n_491) );
AOI22xp33_ASAP7_75t_SL g492 ( .A1(n_411), .A2(n_368), .B1(n_362), .B2(n_372), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_414), .A2(n_383), .B1(n_255), .B2(n_316), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g494 ( .A1(n_414), .A2(n_323), .B1(n_316), .B2(n_369), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_414), .A2(n_383), .B1(n_316), .B2(n_362), .Y(n_495) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_414), .A2(n_368), .B1(n_362), .B2(n_369), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_387), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_387), .B(n_307), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_479), .Y(n_499) );
OAI22xp33_ASAP7_75t_SL g500 ( .A1(n_439), .A2(n_394), .B1(n_414), .B2(n_413), .Y(n_500) );
INVxp67_ASAP7_75t_SL g501 ( .A(n_469), .Y(n_501) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_429), .A2(n_394), .B1(n_368), .B2(n_369), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_477), .A2(n_394), .B1(n_421), .B2(n_420), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_491), .B(n_358), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_435), .B(n_361), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_480), .A2(n_421), .B1(n_420), .B2(n_362), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_479), .B(n_361), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_482), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_481), .A2(n_354), .B1(n_355), .B2(n_316), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_438), .A2(n_316), .B1(n_368), .B2(n_383), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_428), .A2(n_316), .B1(n_368), .B2(n_372), .Y(n_511) );
OAI21xp33_ASAP7_75t_SL g512 ( .A1(n_436), .A2(n_361), .B(n_382), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g513 ( .A1(n_478), .A2(n_368), .B1(n_372), .B2(n_369), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_458), .A2(n_369), .B1(n_372), .B2(n_380), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_452), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_437), .B(n_380), .Y(n_516) );
OAI22xp5_ASAP7_75t_SL g517 ( .A1(n_442), .A2(n_397), .B1(n_372), .B2(n_369), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_443), .A2(n_368), .B1(n_372), .B2(n_369), .Y(n_518) );
OAI22xp33_ASAP7_75t_L g519 ( .A1(n_461), .A2(n_369), .B1(n_372), .B2(n_380), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_454), .A2(n_368), .B1(n_372), .B2(n_369), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_445), .A2(n_368), .B1(n_354), .B2(n_355), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_456), .A2(n_368), .B1(n_312), .B2(n_293), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_431), .A2(n_498), .B1(n_447), .B2(n_453), .Y(n_523) );
OAI221xp5_ASAP7_75t_L g524 ( .A1(n_498), .A2(n_301), .B1(n_293), .B2(n_261), .C(n_299), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_432), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_432), .Y(n_526) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_489), .A2(n_380), .B1(n_382), .B2(n_350), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_472), .A2(n_473), .B1(n_450), .B2(n_478), .Y(n_528) );
OAI221xp5_ASAP7_75t_L g529 ( .A1(n_433), .A2(n_301), .B1(n_293), .B2(n_299), .C(n_250), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_434), .B(n_382), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_457), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_471), .B(n_151), .C(n_145), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_494), .A2(n_444), .B1(n_490), .B2(n_462), .Y(n_533) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_436), .A2(n_486), .B(n_485), .Y(n_534) );
AOI221xp5_ASAP7_75t_L g535 ( .A1(n_475), .A2(n_301), .B1(n_281), .B2(n_285), .C(n_287), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_497), .A2(n_368), .B1(n_312), .B2(n_397), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_434), .B(n_382), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_460), .A2(n_368), .B1(n_312), .B2(n_281), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_460), .A2(n_368), .B1(n_312), .B2(n_281), .Y(n_539) );
OAI221xp5_ASAP7_75t_SL g540 ( .A1(n_446), .A2(n_463), .B1(n_465), .B2(n_488), .C(n_449), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_448), .B(n_312), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_484), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_470), .B(n_338), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_470), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_460), .A2(n_281), .B1(n_349), .B2(n_335), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_495), .A2(n_281), .B1(n_349), .B2(n_335), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_476), .B(n_320), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_430), .B(n_338), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_487), .A2(n_350), .B1(n_338), .B2(n_281), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_487), .A2(n_350), .B1(n_295), .B2(n_298), .Y(n_550) );
OAI221xp5_ASAP7_75t_SL g551 ( .A1(n_439), .A2(n_306), .B1(n_287), .B2(n_285), .C(n_282), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_493), .A2(n_281), .B1(n_349), .B2(n_306), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_430), .B(n_350), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_467), .A2(n_442), .B1(n_455), .B2(n_466), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_468), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_467), .A2(n_281), .B1(n_349), .B2(n_306), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_468), .A2(n_350), .B1(n_320), .B2(n_282), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_468), .A2(n_320), .B1(n_282), .B2(n_317), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_468), .A2(n_320), .B1(n_282), .B2(n_317), .Y(n_559) );
NAND4xp25_ASAP7_75t_L g560 ( .A(n_492), .B(n_285), .C(n_287), .D(n_317), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_441), .B(n_151), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_440), .A2(n_295), .B1(n_298), .B2(n_311), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_474), .A2(n_319), .B1(n_277), .B2(n_287), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_474), .B(n_230), .Y(n_564) );
OAI222xp33_ASAP7_75t_L g565 ( .A1(n_496), .A2(n_319), .B1(n_305), .B2(n_298), .C1(n_295), .C2(n_309), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_459), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_474), .A2(n_319), .B1(n_277), .B2(n_285), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_440), .A2(n_305), .B1(n_309), .B2(n_310), .Y(n_568) );
OAI222xp33_ASAP7_75t_L g569 ( .A1(n_451), .A2(n_305), .B1(n_309), .B2(n_310), .C1(n_292), .C2(n_278), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_459), .B(n_31), .Y(n_570) );
AOI21xp33_ASAP7_75t_L g571 ( .A1(n_474), .A2(n_310), .B(n_151), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_483), .A2(n_277), .B1(n_286), .B2(n_290), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_483), .A2(n_277), .B1(n_286), .B2(n_291), .Y(n_573) );
NOR3xp33_ASAP7_75t_L g574 ( .A(n_464), .B(n_151), .C(n_266), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_483), .A2(n_277), .B1(n_292), .B2(n_313), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_483), .A2(n_292), .B1(n_286), .B2(n_278), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_464), .A2(n_286), .B1(n_321), .B2(n_291), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_491), .B(n_32), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_479), .B(n_151), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_479), .Y(n_580) );
AOI222xp33_ASAP7_75t_L g581 ( .A1(n_475), .A2(n_313), .B1(n_288), .B2(n_314), .C1(n_315), .C2(n_273), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_477), .A2(n_273), .B1(n_296), .B2(n_304), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_479), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_479), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_481), .A2(n_321), .B1(n_291), .B2(n_288), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_469), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_481), .A2(n_321), .B1(n_291), .B2(n_288), .Y(n_587) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_429), .A2(n_283), .B1(n_296), .B2(n_304), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_477), .B(n_145), .C(n_162), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_479), .B(n_153), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_481), .A2(n_291), .B1(n_321), .B2(n_313), .Y(n_591) );
OAI21xp33_ASAP7_75t_L g592 ( .A1(n_540), .A2(n_145), .B(n_162), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_526), .B(n_33), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_526), .B(n_34), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_560), .A2(n_314), .B1(n_321), .B2(n_315), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_544), .B(n_145), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_526), .B(n_35), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_544), .B(n_145), .Y(n_598) );
NAND3xp33_ASAP7_75t_L g599 ( .A(n_532), .B(n_145), .C(n_162), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_515), .B(n_36), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_531), .Y(n_601) );
OAI21xp5_ASAP7_75t_SL g602 ( .A1(n_554), .A2(n_162), .B(n_145), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_530), .B(n_145), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_530), .B(n_145), .Y(n_604) );
OA211x2_ASAP7_75t_L g605 ( .A1(n_586), .A2(n_220), .B(n_322), .C(n_43), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_537), .B(n_145), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_533), .A2(n_283), .B1(n_279), .B2(n_284), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_565), .A2(n_145), .B(n_162), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_534), .B(n_162), .C(n_153), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_542), .B(n_162), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_542), .B(n_162), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_501), .B(n_162), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_525), .B(n_162), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_523), .A2(n_314), .B1(n_153), .B2(n_322), .C(n_315), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_525), .B(n_153), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_499), .B(n_153), .Y(n_616) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_589), .B(n_266), .C(n_322), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_562), .A2(n_315), .B1(n_275), .B2(n_276), .Y(n_618) );
OAI21xp33_ASAP7_75t_L g619 ( .A1(n_512), .A2(n_280), .B(n_279), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_499), .B(n_284), .Y(n_620) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_578), .B(n_300), .C(n_275), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_508), .B(n_580), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_508), .B(n_284), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_534), .A2(n_283), .B1(n_304), .B2(n_296), .Y(n_624) );
OAI21xp33_ASAP7_75t_SL g625 ( .A1(n_581), .A2(n_300), .B(n_284), .Y(n_625) );
OAI21xp5_ASAP7_75t_SL g626 ( .A1(n_549), .A2(n_280), .B(n_279), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g627 ( .A1(n_528), .A2(n_283), .B1(n_300), .B2(n_296), .C(n_304), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_583), .B(n_47), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_504), .B(n_280), .Y(n_629) );
OAI21xp5_ASAP7_75t_SL g630 ( .A1(n_569), .A2(n_279), .B(n_300), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_551), .A2(n_224), .B1(n_217), .B2(n_275), .C(n_276), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_583), .B(n_49), .Y(n_632) );
OAI221xp5_ASAP7_75t_L g633 ( .A1(n_585), .A2(n_283), .B1(n_300), .B2(n_296), .C(n_304), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_584), .B(n_50), .Y(n_634) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_534), .A2(n_283), .B1(n_279), .B2(n_276), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_534), .B(n_276), .C(n_275), .Y(n_636) );
NOR3xp33_ASAP7_75t_L g637 ( .A(n_570), .B(n_276), .C(n_275), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_505), .B(n_52), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_568), .B(n_53), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_587), .A2(n_224), .B1(n_283), .B2(n_272), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_507), .B(n_54), .Y(n_641) );
NAND4xp25_ASAP7_75t_L g642 ( .A(n_591), .B(n_223), .C(n_196), .D(n_193), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_516), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_509), .A2(n_283), .B1(n_272), .B2(n_193), .C(n_182), .Y(n_644) );
OA21x2_ASAP7_75t_L g645 ( .A1(n_520), .A2(n_182), .B(n_57), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_507), .B(n_55), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_588), .B(n_59), .C(n_60), .Y(n_647) );
OAI22xp5_ASAP7_75t_SL g648 ( .A1(n_517), .A2(n_283), .B1(n_63), .B2(n_64), .Y(n_648) );
OAI21xp33_ASAP7_75t_L g649 ( .A1(n_509), .A2(n_62), .B(n_65), .Y(n_649) );
OAI21xp33_ASAP7_75t_L g650 ( .A1(n_500), .A2(n_66), .B(n_67), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_556), .A2(n_68), .B1(n_69), .B2(n_72), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_543), .B(n_73), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_566), .B(n_74), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_541), .B(n_75), .Y(n_654) );
AOI211xp5_ASAP7_75t_SL g655 ( .A1(n_503), .A2(n_76), .B(n_79), .C(n_81), .Y(n_655) );
NOR2xp33_ASAP7_75t_R g656 ( .A(n_555), .B(n_82), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g657 ( .A(n_550), .B(n_83), .C(n_88), .Y(n_657) );
NOR3xp33_ASAP7_75t_SL g658 ( .A(n_529), .B(n_92), .C(n_94), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_548), .B(n_553), .Y(n_659) );
OA21x2_ASAP7_75t_L g660 ( .A1(n_521), .A2(n_95), .B(n_97), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g661 ( .A(n_502), .B(n_536), .C(n_579), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_579), .B(n_547), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_590), .B(n_518), .C(n_575), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_553), .B(n_561), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_561), .B(n_590), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_555), .B(n_514), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_527), .B(n_522), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_506), .B(n_546), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_575), .B(n_519), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_577), .B(n_510), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_513), .B(n_511), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g672 ( .A1(n_582), .A2(n_545), .B(n_564), .Y(n_672) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_538), .A2(n_539), .B(n_573), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_557), .B(n_558), .Y(n_674) );
OA21x2_ASAP7_75t_L g675 ( .A1(n_574), .A2(n_571), .B(n_572), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_559), .B(n_552), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_535), .B(n_524), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_643), .B(n_576), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_592), .A2(n_563), .B1(n_567), .B2(n_625), .Y(n_679) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_635), .B(n_636), .C(n_609), .Y(n_680) );
NAND4xp75_ASAP7_75t_L g681 ( .A(n_605), .B(n_671), .C(n_672), .D(n_673), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_659), .B(n_664), .Y(n_682) );
OAI211xp5_ASAP7_75t_SL g683 ( .A1(n_602), .A2(n_608), .B(n_595), .C(n_624), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_664), .B(n_603), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_661), .B(n_667), .C(n_663), .Y(n_685) );
OA21x2_ASAP7_75t_L g686 ( .A1(n_622), .A2(n_669), .B(n_666), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_604), .B(n_606), .Y(n_687) );
OAI21xp5_ASAP7_75t_L g688 ( .A1(n_630), .A2(n_650), .B(n_626), .Y(n_688) );
AO21x2_ASAP7_75t_L g689 ( .A1(n_593), .A2(n_597), .B(n_613), .Y(n_689) );
AOI211xp5_ASAP7_75t_L g690 ( .A1(n_648), .A2(n_607), .B(n_671), .C(n_656), .Y(n_690) );
AOI211x1_ASAP7_75t_L g691 ( .A1(n_614), .A2(n_668), .B(n_627), .C(n_677), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_662), .B(n_665), .Y(n_692) );
OR2x2_ASAP7_75t_L g693 ( .A(n_615), .B(n_629), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_596), .B(n_598), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_595), .A2(n_618), .B1(n_674), .B2(n_619), .Y(n_695) );
OAI21xp5_ASAP7_75t_L g696 ( .A1(n_655), .A2(n_658), .B(n_649), .Y(n_696) );
XNOR2xp5_ASAP7_75t_L g697 ( .A(n_594), .B(n_676), .Y(n_697) );
NAND4xp25_ASAP7_75t_L g698 ( .A(n_618), .B(n_676), .C(n_616), .D(n_639), .Y(n_698) );
INVx2_ASAP7_75t_SL g699 ( .A(n_656), .Y(n_699) );
NOR3xp33_ASAP7_75t_SL g700 ( .A(n_639), .B(n_647), .C(n_657), .Y(n_700) );
INVxp67_ASAP7_75t_SL g701 ( .A(n_600), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_670), .A2(n_621), .B1(n_637), .B2(n_631), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_620), .B(n_623), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_641), .B(n_652), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_660), .A2(n_675), .B1(n_652), .B2(n_644), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_651), .B(n_638), .C(n_599), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_651), .B(n_617), .C(n_646), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_628), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_628), .B(n_632), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_654), .A2(n_642), .B1(n_640), .B2(n_633), .C(n_653), .Y(n_710) );
AND2x2_ASAP7_75t_SL g711 ( .A(n_645), .B(n_634), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_645), .B(n_640), .Y(n_712) );
AND2x2_ASAP7_75t_SL g713 ( .A(n_666), .B(n_534), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_592), .B(n_635), .C(n_636), .Y(n_714) );
NOR3xp33_ASAP7_75t_SL g715 ( .A(n_592), .B(n_442), .C(n_602), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_601), .Y(n_716) );
XNOR2xp5_ASAP7_75t_SL g717 ( .A(n_648), .B(n_442), .Y(n_717) );
OAI211xp5_ASAP7_75t_L g718 ( .A1(n_625), .A2(n_602), .B(n_608), .C(n_630), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_643), .B(n_601), .Y(n_719) );
AOI22xp33_ASAP7_75t_SL g720 ( .A1(n_671), .A2(n_534), .B1(n_636), .B2(n_625), .Y(n_720) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_671), .A2(n_534), .B1(n_636), .B2(n_625), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_592), .A2(n_625), .B1(n_671), .B2(n_607), .Y(n_722) );
OA211x2_ASAP7_75t_L g723 ( .A1(n_650), .A2(n_554), .B(n_649), .C(n_619), .Y(n_723) );
OAI21xp33_ASAP7_75t_L g724 ( .A1(n_592), .A2(n_635), .B(n_624), .Y(n_724) );
BUFx2_ASAP7_75t_L g725 ( .A(n_656), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_592), .B(n_442), .Y(n_726) );
NOR3xp33_ASAP7_75t_L g727 ( .A(n_592), .B(n_608), .C(n_602), .Y(n_727) );
NAND4xp75_ASAP7_75t_L g728 ( .A(n_625), .B(n_605), .C(n_671), .D(n_534), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_659), .B(n_664), .Y(n_729) );
INVx5_ASAP7_75t_L g730 ( .A(n_603), .Y(n_730) );
AO21x2_ASAP7_75t_L g731 ( .A1(n_612), .A2(n_611), .B(n_610), .Y(n_731) );
NAND3xp33_ASAP7_75t_L g732 ( .A(n_685), .B(n_720), .C(n_721), .Y(n_732) );
NAND4xp75_ASAP7_75t_L g733 ( .A(n_723), .B(n_688), .C(n_699), .D(n_691), .Y(n_733) );
OA22x2_ASAP7_75t_L g734 ( .A1(n_725), .A2(n_697), .B1(n_688), .B2(n_701), .Y(n_734) );
XOR2x2_ASAP7_75t_L g735 ( .A(n_717), .B(n_681), .Y(n_735) );
XOR2x2_ASAP7_75t_L g736 ( .A(n_690), .B(n_728), .Y(n_736) );
NAND4xp75_ASAP7_75t_L g737 ( .A(n_713), .B(n_696), .C(n_715), .D(n_700), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_718), .A2(n_695), .B1(n_683), .B2(n_722), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_686), .B(n_682), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_716), .Y(n_740) );
INVx3_ASAP7_75t_L g741 ( .A(n_730), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_720), .B(n_721), .C(n_705), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_686), .B(n_729), .Y(n_743) );
INVxp67_ASAP7_75t_L g744 ( .A(n_726), .Y(n_744) );
OR2x2_ASAP7_75t_L g745 ( .A(n_692), .B(n_719), .Y(n_745) );
AND2x4_ASAP7_75t_SL g746 ( .A(n_687), .B(n_684), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_695), .A2(n_698), .B1(n_702), .B2(n_727), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_678), .Y(n_748) );
XNOR2x2_ASAP7_75t_L g749 ( .A(n_707), .B(n_712), .Y(n_749) );
XOR2xp5_ASAP7_75t_L g750 ( .A(n_693), .B(n_702), .Y(n_750) );
XOR2x2_ASAP7_75t_L g751 ( .A(n_727), .B(n_711), .Y(n_751) );
XNOR2xp5_ASAP7_75t_L g752 ( .A(n_704), .B(n_679), .Y(n_752) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_748), .Y(n_753) );
INVx1_ASAP7_75t_SL g754 ( .A(n_746), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_740), .Y(n_755) );
XOR2xp5_ASAP7_75t_L g756 ( .A(n_735), .B(n_703), .Y(n_756) );
XOR2x2_ASAP7_75t_L g757 ( .A(n_736), .B(n_714), .Y(n_757) );
INVx1_ASAP7_75t_SL g758 ( .A(n_746), .Y(n_758) );
INVxp67_ASAP7_75t_L g759 ( .A(n_733), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_739), .B(n_689), .Y(n_760) );
AO22x2_ASAP7_75t_L g761 ( .A1(n_732), .A2(n_680), .B1(n_694), .B2(n_708), .Y(n_761) );
XNOR2x1_ASAP7_75t_L g762 ( .A(n_736), .B(n_706), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_745), .Y(n_763) );
AO22x2_ASAP7_75t_L g764 ( .A1(n_742), .A2(n_694), .B1(n_709), .B2(n_705), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_738), .A2(n_724), .B1(n_710), .B2(n_731), .Y(n_765) );
INVxp67_ASAP7_75t_L g766 ( .A(n_733), .Y(n_766) );
XNOR2xp5_ASAP7_75t_L g767 ( .A(n_738), .B(n_710), .Y(n_767) );
XOR2x2_ASAP7_75t_L g768 ( .A(n_757), .B(n_751), .Y(n_768) );
OA22x2_ASAP7_75t_L g769 ( .A1(n_765), .A2(n_747), .B1(n_750), .B2(n_752), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_763), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_762), .A2(n_747), .B1(n_734), .B2(n_737), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_753), .Y(n_772) );
OA22x2_ASAP7_75t_L g773 ( .A1(n_756), .A2(n_749), .B1(n_744), .B2(n_743), .Y(n_773) );
INVx2_ASAP7_75t_SL g774 ( .A(n_754), .Y(n_774) );
AOI22x1_ASAP7_75t_L g775 ( .A1(n_761), .A2(n_741), .B1(n_743), .B2(n_739), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_755), .Y(n_776) );
AOI22x1_ASAP7_75t_L g777 ( .A1(n_767), .A2(n_759), .B1(n_766), .B2(n_764), .Y(n_777) );
INVx4_ASAP7_75t_L g778 ( .A(n_757), .Y(n_778) );
INVx1_ASAP7_75t_SL g779 ( .A(n_774), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_774), .Y(n_780) );
INVx1_ASAP7_75t_SL g781 ( .A(n_768), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_772), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_770), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_776), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_776), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_775), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_780), .Y(n_787) );
INVx1_ASAP7_75t_SL g788 ( .A(n_779), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_782), .Y(n_789) );
OA22x2_ASAP7_75t_L g790 ( .A1(n_781), .A2(n_771), .B1(n_778), .B2(n_767), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_782), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_788), .B(n_778), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_790), .A2(n_769), .B1(n_768), .B2(n_778), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_788), .Y(n_794) );
NOR2x1_ASAP7_75t_L g795 ( .A(n_794), .B(n_787), .Y(n_795) );
INVxp67_ASAP7_75t_L g796 ( .A(n_792), .Y(n_796) );
NOR2xp67_ASAP7_75t_L g797 ( .A(n_796), .B(n_793), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_795), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_798), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_797), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_800), .A2(n_769), .B1(n_762), .B2(n_773), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_801), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_802), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_803), .A2(n_799), .B1(n_789), .B2(n_791), .Y(n_804) );
INVxp67_ASAP7_75t_SL g805 ( .A(n_804), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_805), .A2(n_786), .B1(n_777), .B2(n_783), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_806), .Y(n_807) );
AOI221xp5_ASAP7_75t_L g808 ( .A1(n_807), .A2(n_786), .B1(n_785), .B2(n_784), .C(n_758), .Y(n_808) );
AOI211xp5_ASAP7_75t_L g809 ( .A1(n_808), .A2(n_785), .B(n_784), .C(n_760), .Y(n_809) );
endmodule