module real_jpeg_11391_n_19 (n_17, n_8, n_116, n_0, n_2, n_10, n_114, n_9, n_12, n_6, n_121, n_11, n_14, n_120, n_7, n_117, n_18, n_3, n_119, n_5, n_4, n_115, n_122, n_1, n_118, n_16, n_15, n_13, n_113, n_19);

input n_17;
input n_8;
input n_116;
input n_0;
input n_2;
input n_10;
input n_114;
input n_9;
input n_12;
input n_6;
input n_121;
input n_11;
input n_14;
input n_120;
input n_7;
input n_117;
input n_18;
input n_3;
input n_119;
input n_5;
input n_4;
input n_115;
input n_122;
input n_1;
input n_118;
input n_16;
input n_15;
input n_13;
input n_113;

output n_19;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_1),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_1),
.B(n_47),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_2),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_2),
.B(n_80),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_3),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_3),
.B(n_89),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_4),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_5),
.Y(n_82)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_5),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_7),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_7),
.B(n_86),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_9),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_9),
.B(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_10),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_10),
.B(n_97),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_12),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_12),
.B(n_65),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_14),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_15),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_15),
.B(n_57),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_17),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_17),
.B(n_53),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_23),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_54),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_28),
.B(n_102),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_35),
.B(n_37),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_111),
.Y(n_38)
);

NAND3xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_105),
.C(n_110),
.Y(n_39)
);

NAND4xp25_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_46),
.C(n_51),
.D(n_55),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_41),
.A2(n_46),
.B(n_106),
.C(n_109),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_42),
.B(n_43),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_49),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_52),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_100),
.B(n_104),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_96),
.B(n_99),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_84),
.B(n_93),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_79),
.B(n_83),
.Y(n_62)
);

OA21x2_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_68),
.B(n_78),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B(n_77),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_103),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_113),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_114),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_115),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_116),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_117),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_118),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_119),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_120),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_121),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_122),
.Y(n_102)
);


endmodule