module fake_jpeg_22989_n_277 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_8),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_25),
.B1(n_32),
.B2(n_29),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_27),
.B1(n_22),
.B2(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_25),
.B1(n_33),
.B2(n_32),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_49),
.A2(n_56),
.B(n_38),
.Y(n_98)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_50),
.B(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_28),
.Y(n_64)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_55),
.B(n_9),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_18),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_24),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_27),
.B1(n_29),
.B2(n_33),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_22),
.B1(n_20),
.B2(n_26),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_95),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_65),
.A2(n_74),
.B1(n_98),
.B2(n_5),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_76),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_67),
.B(n_69),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_56),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_68),
.A2(n_88),
.B(n_6),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_72),
.B(n_75),
.Y(n_118)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_77),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_17),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_78),
.B(n_81),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_63),
.B1(n_43),
.B2(n_60),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_79),
.A2(n_85),
.B1(n_99),
.B2(n_5),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_16),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_43),
.B(n_26),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_82),
.B(n_91),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_31),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_31),
.B1(n_16),
.B2(n_15),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_89),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_19),
.B1(n_24),
.B2(n_2),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_10),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_97),
.Y(n_128)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_15),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_51),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_47),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_0),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_95),
.Y(n_125)
);

NAND2x1_ASAP7_75t_SL g105 ( 
.A(n_68),
.B(n_0),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_105),
.A2(n_129),
.B(n_8),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_115),
.Y(n_135)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_0),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_64),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_121),
.Y(n_140)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_3),
.C(n_4),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_101),
.C(n_93),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_126),
.B1(n_99),
.B2(n_75),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_66),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_70),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_130),
.A2(n_134),
.B(n_154),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_83),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_97),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_132),
.B(n_143),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_138),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_80),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_141),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_68),
.C(n_72),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_83),
.C(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_76),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_153),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_86),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_65),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_155),
.B1(n_112),
.B2(n_85),
.Y(n_160)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_149),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_100),
.C(n_84),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_124),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_74),
.Y(n_151)
);

AO22x1_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_88),
.B1(n_79),
.B2(n_84),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_105),
.B(n_119),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_88),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_77),
.B1(n_81),
.B2(n_78),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_91),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_160),
.A2(n_180),
.B1(n_182),
.B2(n_147),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_164),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_156),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_165),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_140),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_166),
.B(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_122),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_144),
.Y(n_187)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_183),
.Y(n_191)
);

AOI211xp5_ASAP7_75t_SL g199 ( 
.A1(n_174),
.A2(n_159),
.B(n_180),
.C(n_162),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_153),
.A2(n_112),
.B1(n_105),
.B2(n_120),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_176),
.B1(n_133),
.B2(n_130),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_117),
.B1(n_125),
.B2(n_113),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_119),
.B(n_108),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_152),
.A2(n_117),
.B(n_113),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_104),
.B(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_146),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_137),
.C(n_131),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_187),
.Y(n_211)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_172),
.A2(n_104),
.B1(n_142),
.B2(n_141),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_190),
.A2(n_166),
.B1(n_184),
.B2(n_178),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_177),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_157),
.Y(n_193)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_196),
.Y(n_210)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_201),
.Y(n_209)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_174),
.B(n_170),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_175),
.B1(n_176),
.B2(n_174),
.Y(n_218)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_207),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_148),
.B1(n_89),
.B2(n_87),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_206),
.Y(n_208)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_165),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_217),
.Y(n_240)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_187),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_161),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_218),
.A2(n_219),
.B(n_189),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_197),
.A2(n_160),
.B1(n_170),
.B2(n_179),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_224),
.B1(n_196),
.B2(n_203),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_161),
.B1(n_168),
.B2(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_168),
.B1(n_171),
.B2(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_205),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_218),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_207),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_237),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_186),
.C(n_192),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_231),
.C(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_193),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_199),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_235),
.C(n_221),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_201),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_236),
.B(n_222),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_109),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_188),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_238),
.A2(n_239),
.B(n_221),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_210),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_241),
.B(n_234),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_220),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_246),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_248),
.C(n_250),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_249),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_216),
.Y(n_249)
);

INVxp33_ASAP7_75t_SL g250 ( 
.A(n_240),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_233),
.C(n_232),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_254),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_230),
.C(n_236),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_219),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_244),
.B(n_211),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_256),
.A2(n_257),
.B1(n_242),
.B2(n_214),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_243),
.B(n_230),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_259),
.B(n_251),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_262),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_208),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_194),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_258),
.B(n_209),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

AOI31xp33_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_245),
.A3(n_194),
.B(n_227),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_268),
.A3(n_269),
.B1(n_194),
.B2(n_109),
.C1(n_11),
.C2(n_13),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_266),
.A2(n_265),
.B(n_263),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_11),
.C(n_14),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_272),
.B1(n_10),
.B2(n_11),
.Y(n_273)
);

AOI21x1_ASAP7_75t_L g272 ( 
.A1(n_269),
.A2(n_9),
.B(n_10),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_274),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_14),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_276),
.Y(n_277)
);


endmodule