module fake_ariane_2903_n_932 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_932);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_932;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_283;
wire n_919;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_731;
wire n_336;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_928;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_365;
wire n_455;
wire n_238;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_861;
wire n_780;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_856;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_54),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_75),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_145),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_85),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_43),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_89),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_92),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_176),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_53),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_109),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_104),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_73),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_25),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_125),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_27),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_87),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_159),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_184),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_91),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_30),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_77),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_114),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_11),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_41),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g218 ( 
.A(n_122),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_106),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_115),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_76),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_8),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_172),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_160),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_19),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_0),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_56),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_2),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_146),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_97),
.Y(n_232)
);

BUFx2_ASAP7_75t_SL g233 ( 
.A(n_182),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_46),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_94),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_44),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_173),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_110),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_139),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_103),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_27),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_67),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_14),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_80),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_118),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_3),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_64),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_50),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_142),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_121),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_131),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_130),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_63),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_116),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_132),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_55),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_141),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_72),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_171),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_29),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_29),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_136),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_90),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_13),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_0),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_124),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_23),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_38),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_1),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_69),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_128),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_28),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_58),
.Y(n_273)
);

BUFx8_ASAP7_75t_SL g274 ( 
.A(n_40),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_150),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_157),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_86),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_16),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_18),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_25),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_51),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_144),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_2),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_225),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_226),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_269),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_279),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_243),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_243),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_274),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_194),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g295 ( 
.A(n_203),
.B(n_1),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_274),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_209),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_210),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_206),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_243),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_202),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_258),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_269),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_263),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_266),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_188),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_216),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_186),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_190),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_212),
.B(n_3),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_222),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_191),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_201),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_241),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_208),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_246),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_261),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_214),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_248),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_264),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_265),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_267),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_231),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_272),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_232),
.B(n_4),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_278),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_280),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_213),
.B(n_4),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_248),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_185),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_188),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_240),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_187),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_239),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_247),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_250),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_253),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_239),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_256),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_257),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_192),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_259),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_193),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_281),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_195),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_213),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_196),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_305),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_337),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_284),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_R g354 ( 
.A(n_293),
.B(n_197),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_327),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_307),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_285),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_344),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_286),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_344),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_290),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_308),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_322),
.B(n_270),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_270),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_346),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_308),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_349),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_296),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_333),
.B(n_189),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_336),
.B(n_204),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_308),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_327),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_309),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_346),
.Y(n_376)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_347),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_198),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_291),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_329),
.B(n_199),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_292),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_287),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_301),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_348),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_302),
.A2(n_221),
.B1(n_255),
.B2(n_233),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_303),
.B(n_200),
.Y(n_389)
);

AND2x2_ASAP7_75t_SL g390 ( 
.A(n_313),
.B(n_229),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_312),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_316),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_287),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_326),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_314),
.B(n_205),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_348),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_335),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_338),
.B(n_207),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_288),
.B(n_211),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_317),
.B(n_215),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_332),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_339),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_289),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_289),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_408),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_352),
.B(n_304),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_408),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_390),
.B(n_319),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_408),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_320),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_L g415 ( 
.A(n_370),
.B(n_323),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_408),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_355),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_375),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_385),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_397),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_364),
.B(n_306),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_390),
.B(n_342),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_324),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_372),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_385),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_353),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_379),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_351),
.B(n_300),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_383),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_389),
.B(n_325),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

BUFx4f_ASAP7_75t_L g434 ( 
.A(n_364),
.Y(n_434)
);

BUFx10_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_379),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_364),
.B(n_343),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_356),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_383),
.Y(n_440)
);

AND2x6_ASAP7_75t_L g441 ( 
.A(n_397),
.B(n_229),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_398),
.B(n_345),
.Y(n_443)
);

INVx5_ASAP7_75t_L g444 ( 
.A(n_372),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_359),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_356),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_397),
.B(n_334),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_403),
.B(n_330),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_229),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_358),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_381),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_361),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_393),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_405),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_393),
.A2(n_328),
.B1(n_331),
.B2(n_310),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_358),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_374),
.Y(n_458)
);

AND2x6_ASAP7_75t_L g459 ( 
.A(n_405),
.B(n_332),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

INVxp33_ASAP7_75t_L g461 ( 
.A(n_354),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_371),
.B(n_334),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_383),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_378),
.B(n_295),
.C(n_219),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_360),
.Y(n_465)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_395),
.B(n_400),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_377),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_387),
.B(n_298),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_395),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_384),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_400),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_404),
.B(n_360),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_391),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_365),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_377),
.Y(n_475)
);

OR2x6_ASAP7_75t_L g476 ( 
.A(n_363),
.B(n_294),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_382),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_392),
.B(n_217),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_362),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_431),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_388),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_420),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_443),
.B(n_380),
.Y(n_483)
);

A2O1A1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_424),
.A2(n_394),
.B(n_367),
.C(n_365),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_420),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_L g486 ( 
.A(n_448),
.B(n_218),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_409),
.Y(n_487)
);

OAI22x1_ASAP7_75t_L g488 ( 
.A1(n_450),
.A2(n_386),
.B1(n_376),
.B2(n_399),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_431),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_412),
.A2(n_376),
.B1(n_386),
.B2(n_399),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_424),
.B(n_377),
.Y(n_491)
);

AND3x1_ASAP7_75t_L g492 ( 
.A(n_414),
.B(n_404),
.C(n_396),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_434),
.A2(n_421),
.B1(n_455),
.B2(n_432),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_426),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_423),
.B(n_377),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_418),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_434),
.B(n_410),
.Y(n_497)
);

NAND2xp33_ASAP7_75t_L g498 ( 
.A(n_461),
.B(n_218),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_410),
.B(n_377),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_297),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_466),
.A2(n_362),
.B1(n_366),
.B2(n_373),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_426),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_461),
.B(n_220),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_462),
.A2(n_252),
.B1(n_223),
.B2(n_224),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_421),
.B(n_5),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_455),
.B(n_227),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_422),
.A2(n_262),
.B1(n_230),
.B2(n_234),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_470),
.A2(n_407),
.B1(n_406),
.B2(n_396),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_438),
.B(n_235),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_428),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_422),
.A2(n_271),
.B1(n_236),
.B2(n_237),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_430),
.B(n_384),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_447),
.B(n_238),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_427),
.B(n_242),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_442),
.B(n_244),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_447),
.B(n_406),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_478),
.B(n_446),
.Y(n_517)
);

O2A1O1Ixp33_ASAP7_75t_L g518 ( 
.A1(n_445),
.A2(n_366),
.B(n_373),
.C(n_7),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_468),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_476),
.B(n_407),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_452),
.A2(n_473),
.B1(n_478),
.B2(n_464),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_428),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_429),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_453),
.B(n_245),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_469),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_435),
.B(n_249),
.Y(n_526)
);

NAND2x1_ASAP7_75t_L g527 ( 
.A(n_466),
.B(n_372),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_L g528 ( 
.A(n_459),
.B(n_466),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_457),
.Y(n_529)
);

NOR2x1p5_ASAP7_75t_L g530 ( 
.A(n_465),
.B(n_251),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_456),
.A2(n_277),
.B1(n_276),
.B2(n_275),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_411),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_L g533 ( 
.A(n_459),
.B(n_218),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_471),
.B(n_254),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_458),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_429),
.Y(n_536)
);

OAI22xp33_ASAP7_75t_L g537 ( 
.A1(n_437),
.A2(n_439),
.B1(n_476),
.B2(n_458),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_466),
.A2(n_218),
.B1(n_273),
.B2(n_268),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_436),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_417),
.B(n_5),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_437),
.Y(n_541)
);

NOR3x1_ASAP7_75t_L g542 ( 
.A(n_472),
.B(n_6),
.C(n_7),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_440),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_435),
.B(n_282),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_463),
.B(n_218),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_477),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_439),
.B(n_218),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_466),
.A2(n_218),
.B1(n_8),
.B2(n_9),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_416),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_436),
.Y(n_550)
);

NOR3xp33_ASAP7_75t_SL g551 ( 
.A(n_517),
.B(n_474),
.C(n_419),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_535),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_523),
.Y(n_553)
);

NOR3xp33_ASAP7_75t_SL g554 ( 
.A(n_484),
.B(n_474),
.C(n_415),
.Y(n_554)
);

BUFx12f_ASAP7_75t_L g555 ( 
.A(n_520),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_487),
.Y(n_556)
);

O2A1O1Ixp33_ASAP7_75t_L g557 ( 
.A1(n_541),
.A2(n_456),
.B(n_411),
.C(n_468),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_536),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_497),
.B(n_459),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_493),
.B(n_417),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_487),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_481),
.B(n_459),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_520),
.B(n_476),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_487),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_539),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_496),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_541),
.B(n_409),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_549),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_481),
.B(n_459),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_527),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_R g571 ( 
.A(n_529),
.B(n_409),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_500),
.B(n_451),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_516),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_483),
.B(n_451),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_504),
.B(n_454),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_550),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_519),
.B(n_409),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_502),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_535),
.B(n_454),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_516),
.B(n_460),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_532),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_532),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_510),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_537),
.B(n_513),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_512),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_530),
.B(n_413),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_520),
.B(n_492),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_537),
.B(n_480),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_R g589 ( 
.A(n_533),
.B(n_528),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_508),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_505),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_489),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_482),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_522),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_490),
.B(n_488),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_547),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_521),
.B(n_413),
.Y(n_597)
);

BUFx4f_ASAP7_75t_L g598 ( 
.A(n_525),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_509),
.B(n_505),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_507),
.B(n_460),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_485),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_494),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_514),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_546),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_540),
.Y(n_605)
);

AND2x6_ASAP7_75t_SL g606 ( 
.A(n_540),
.B(n_6),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_515),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_543),
.B(n_413),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_R g609 ( 
.A(n_498),
.B(n_413),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_552),
.B(n_542),
.Y(n_610)
);

OAI21x1_ASAP7_75t_L g611 ( 
.A1(n_560),
.A2(n_545),
.B(n_495),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_572),
.B(n_499),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_560),
.A2(n_491),
.B(n_501),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_599),
.B(n_538),
.Y(n_614)
);

NOR2x1_ASAP7_75t_SL g615 ( 
.A(n_582),
.B(n_526),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_562),
.A2(n_534),
.B(n_524),
.Y(n_616)
);

AO21x1_ASAP7_75t_L g617 ( 
.A1(n_569),
.A2(n_486),
.B(n_518),
.Y(n_617)
);

NAND2x1p5_ASAP7_75t_L g618 ( 
.A(n_598),
.B(n_544),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_561),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_559),
.A2(n_506),
.B(n_503),
.Y(n_620)
);

BUFx4f_ASAP7_75t_L g621 ( 
.A(n_555),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_597),
.B(n_548),
.Y(n_622)
);

OAI21x1_ASAP7_75t_L g623 ( 
.A1(n_570),
.A2(n_501),
.B(n_479),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_568),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_588),
.B(n_538),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_571),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_607),
.B(n_511),
.Y(n_627)
);

AND2x6_ASAP7_75t_SL g628 ( 
.A(n_587),
.B(n_548),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_570),
.A2(n_479),
.B(n_518),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_605),
.A2(n_531),
.B1(n_433),
.B2(n_425),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_598),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_597),
.A2(n_603),
.B(n_567),
.Y(n_632)
);

OA21x2_ASAP7_75t_L g633 ( 
.A1(n_574),
.A2(n_433),
.B(n_425),
.Y(n_633)
);

OAI21xp33_ASAP7_75t_L g634 ( 
.A1(n_591),
.A2(n_9),
.B(n_10),
.Y(n_634)
);

AOI31xp67_ASAP7_75t_L g635 ( 
.A1(n_601),
.A2(n_433),
.A3(n_425),
.B(n_449),
.Y(n_635)
);

AOI221x1_ASAP7_75t_L g636 ( 
.A1(n_584),
.A2(n_433),
.B1(n_425),
.B2(n_475),
.C(n_467),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_590),
.B(n_10),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_570),
.A2(n_444),
.B(n_449),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_573),
.B(n_11),
.Y(n_639)
);

AOI21xp33_ASAP7_75t_L g640 ( 
.A1(n_584),
.A2(n_444),
.B(n_13),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_566),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_571),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_567),
.A2(n_475),
.B(n_467),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_588),
.B(n_441),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_601),
.A2(n_444),
.B(n_449),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_551),
.B(n_444),
.Y(n_646)
);

O2A1O1Ixp5_ASAP7_75t_L g647 ( 
.A1(n_575),
.A2(n_449),
.B(n_441),
.C(n_15),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_585),
.B(n_12),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_564),
.Y(n_649)
);

OAI21x1_ASAP7_75t_L g650 ( 
.A1(n_608),
.A2(n_449),
.B(n_441),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_579),
.B(n_441),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_593),
.Y(n_652)
);

OA22x2_ASAP7_75t_L g653 ( 
.A1(n_563),
.A2(n_441),
.B1(n_14),
.B2(n_15),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_L g654 ( 
.A1(n_600),
.A2(n_12),
.B(n_16),
.Y(n_654)
);

AO31x2_ASAP7_75t_L g655 ( 
.A1(n_553),
.A2(n_102),
.A3(n_178),
.B(n_177),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_L g656 ( 
.A(n_622),
.B(n_554),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_652),
.Y(n_657)
);

O2A1O1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_634),
.A2(n_595),
.B(n_557),
.C(n_596),
.Y(n_658)
);

NAND2x1p5_ASAP7_75t_L g659 ( 
.A(n_631),
.B(n_582),
.Y(n_659)
);

O2A1O1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_634),
.A2(n_596),
.B(n_592),
.C(n_586),
.Y(n_660)
);

OAI21x1_ASAP7_75t_L g661 ( 
.A1(n_611),
.A2(n_578),
.B(n_583),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_641),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_624),
.Y(n_663)
);

NAND2x1p5_ASAP7_75t_L g664 ( 
.A(n_631),
.B(n_582),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_649),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_632),
.A2(n_592),
.B(n_586),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_645),
.A2(n_578),
.B(n_583),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_613),
.A2(n_594),
.B(n_556),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_648),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_614),
.A2(n_586),
.B(n_580),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_629),
.A2(n_594),
.B(n_556),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_649),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_653),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_654),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_654),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_616),
.A2(n_556),
.B(n_553),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_650),
.A2(n_558),
.B(n_565),
.Y(n_677)
);

AND2x6_ASAP7_75t_L g678 ( 
.A(n_625),
.B(n_602),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_627),
.B(n_563),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_614),
.A2(n_604),
.B(n_587),
.C(n_602),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_642),
.B(n_577),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_626),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_639),
.Y(n_683)
);

CKINVDCx11_ASAP7_75t_R g684 ( 
.A(n_649),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_621),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_620),
.A2(n_558),
.B(n_565),
.Y(n_686)
);

OAI21x1_ASAP7_75t_SL g687 ( 
.A1(n_615),
.A2(n_561),
.B(n_576),
.Y(n_687)
);

OAI21xp33_ASAP7_75t_SL g688 ( 
.A1(n_625),
.A2(n_561),
.B(n_576),
.Y(n_688)
);

O2A1O1Ixp33_ASAP7_75t_SL g689 ( 
.A1(n_640),
.A2(n_589),
.B(n_606),
.C(n_582),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_621),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_622),
.B(n_563),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_623),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_622),
.B(n_563),
.Y(n_693)
);

A2O1A1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_640),
.A2(n_587),
.B(n_602),
.C(n_577),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_618),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_618),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_638),
.A2(n_589),
.B(n_609),
.Y(n_697)
);

NAND2x1_ASAP7_75t_L g698 ( 
.A(n_687),
.B(n_619),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_682),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_SL g700 ( 
.A(n_674),
.B(n_630),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_691),
.B(n_619),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_683),
.B(n_637),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_669),
.B(n_610),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_692),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_661),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_SL g706 ( 
.A(n_675),
.B(n_630),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_665),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_656),
.A2(n_622),
.B1(n_555),
.B2(n_612),
.Y(n_708)
);

AOI221xp5_ASAP7_75t_L g709 ( 
.A1(n_689),
.A2(n_612),
.B1(n_617),
.B2(n_647),
.C(n_644),
.Y(n_709)
);

OA21x2_ASAP7_75t_L g710 ( 
.A1(n_668),
.A2(n_636),
.B(n_644),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_691),
.A2(n_602),
.B1(n_577),
.B2(n_628),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_662),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_657),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_684),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_676),
.Y(n_715)
);

AOI221xp5_ASAP7_75t_L g716 ( 
.A1(n_689),
.A2(n_651),
.B1(n_646),
.B2(n_628),
.C(n_581),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_669),
.A2(n_582),
.B1(n_651),
.B2(n_581),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_679),
.B(n_17),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_665),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_688),
.A2(n_643),
.B(n_633),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_680),
.B(n_635),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_686),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_SL g723 ( 
.A(n_682),
.B(n_609),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_685),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_663),
.Y(n_725)
);

CKINVDCx16_ASAP7_75t_R g726 ( 
.A(n_690),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_SL g727 ( 
.A1(n_693),
.A2(n_633),
.B1(n_581),
.B2(n_655),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_673),
.A2(n_581),
.B1(n_564),
.B2(n_655),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_665),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_679),
.B(n_564),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_693),
.B(n_655),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_670),
.A2(n_564),
.B1(n_18),
.B2(n_19),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_694),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_665),
.Y(n_734)
);

CKINVDCx11_ASAP7_75t_R g735 ( 
.A(n_695),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_694),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_696),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_658),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_678),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_SL g740 ( 
.A1(n_680),
.A2(n_24),
.B(n_26),
.C(n_28),
.Y(n_740)
);

OAI211xp5_ASAP7_75t_L g741 ( 
.A1(n_658),
.A2(n_26),
.B(n_30),
.C(n_179),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_678),
.A2(n_681),
.B1(n_666),
.B2(n_677),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_681),
.B(n_31),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_667),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_671),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_672),
.B(n_32),
.Y(n_746)
);

AO21x2_ASAP7_75t_L g747 ( 
.A1(n_728),
.A2(n_660),
.B(n_697),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_733),
.A2(n_678),
.B1(n_672),
.B2(n_664),
.Y(n_748)
);

OAI211xp5_ASAP7_75t_L g749 ( 
.A1(n_741),
.A2(n_660),
.B(n_678),
.C(n_664),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_732),
.A2(n_659),
.B1(n_678),
.B2(n_35),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_700),
.A2(n_659),
.B(n_34),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_708),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_718),
.B(n_39),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_699),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_736),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_755)
);

OAI21x1_ASAP7_75t_L g756 ( 
.A1(n_720),
.A2(n_48),
.B(n_49),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_734),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_731),
.B(n_52),
.Y(n_758)
);

OA21x2_ASAP7_75t_L g759 ( 
.A1(n_744),
.A2(n_745),
.B(n_705),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_738),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_730),
.B(n_61),
.Y(n_761)
);

OAI21x1_ASAP7_75t_L g762 ( 
.A1(n_744),
.A2(n_62),
.B(n_65),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_731),
.A2(n_66),
.B1(n_68),
.B2(n_70),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_739),
.B(n_71),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_739),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_714),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_702),
.B(n_74),
.Y(n_767)
);

AO221x1_ASAP7_75t_L g768 ( 
.A1(n_739),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.C(n_82),
.Y(n_768)
);

AO21x1_ASAP7_75t_SL g769 ( 
.A1(n_742),
.A2(n_83),
.B(n_84),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_SL g770 ( 
.A1(n_724),
.A2(n_88),
.B(n_93),
.C(n_95),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_703),
.B(n_96),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_700),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_706),
.A2(n_101),
.B1(n_105),
.B2(n_107),
.Y(n_773)
);

OAI22xp33_ASAP7_75t_L g774 ( 
.A1(n_714),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_713),
.B(n_725),
.Y(n_775)
);

AO21x2_ASAP7_75t_L g776 ( 
.A1(n_705),
.A2(n_117),
.B(n_119),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_737),
.B(n_120),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_706),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_711),
.A2(n_129),
.B1(n_133),
.B2(n_134),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_716),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_780)
);

OA21x2_ASAP7_75t_L g781 ( 
.A1(n_745),
.A2(n_140),
.B(n_143),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_717),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_704),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_701),
.B(n_151),
.Y(n_784)
);

OAI221xp5_ASAP7_75t_L g785 ( 
.A1(n_773),
.A2(n_740),
.B1(n_712),
.B2(n_709),
.C(n_723),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_765),
.B(n_721),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_783),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_783),
.Y(n_788)
);

NOR2x1_ASAP7_75t_L g789 ( 
.A(n_766),
.B(n_729),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_775),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_768),
.A2(n_701),
.B1(n_735),
.B2(n_721),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_754),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_765),
.B(n_721),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_759),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_758),
.B(n_721),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_758),
.B(n_710),
.Y(n_796)
);

AND2x4_ASAP7_75t_SL g797 ( 
.A(n_757),
.B(n_701),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_757),
.B(n_715),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_766),
.B(n_710),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_759),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_759),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_757),
.B(n_710),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_759),
.B(n_704),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_757),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_757),
.B(n_715),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_747),
.B(n_722),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_781),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_781),
.Y(n_808)
);

NAND2x1_ASAP7_75t_L g809 ( 
.A(n_768),
.B(n_734),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_767),
.B(n_771),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_747),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_747),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_794),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_792),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_799),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_SL g816 ( 
.A1(n_785),
.A2(n_773),
.B(n_784),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_790),
.Y(n_817)
);

CKINVDCx8_ASAP7_75t_R g818 ( 
.A(n_798),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_790),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_788),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_L g821 ( 
.A(n_811),
.B(n_740),
.C(n_760),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_804),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_787),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_787),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_799),
.Y(n_825)
);

AOI211xp5_ASAP7_75t_L g826 ( 
.A1(n_810),
.A2(n_770),
.B(n_774),
.C(n_750),
.Y(n_826)
);

AOI221xp5_ASAP7_75t_L g827 ( 
.A1(n_811),
.A2(n_767),
.B1(n_753),
.B2(n_771),
.C(n_752),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_796),
.B(n_729),
.Y(n_828)
);

OR2x6_ASAP7_75t_L g829 ( 
.A(n_809),
.B(n_784),
.Y(n_829)
);

AOI222xp33_ASAP7_75t_L g830 ( 
.A1(n_796),
.A2(n_749),
.B1(n_763),
.B2(n_755),
.C1(n_761),
.C2(n_772),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_795),
.B(n_714),
.Y(n_831)
);

AND2x2_ASAP7_75t_SL g832 ( 
.A(n_831),
.B(n_795),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_829),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_815),
.B(n_786),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_815),
.B(n_786),
.Y(n_835)
);

OR2x2_ASAP7_75t_L g836 ( 
.A(n_825),
.B(n_788),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_814),
.B(n_802),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_814),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_825),
.B(n_793),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_822),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_822),
.B(n_793),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_822),
.B(n_802),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_828),
.B(n_805),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_836),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_833),
.B(n_789),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_838),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_841),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_837),
.B(n_817),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_836),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_846),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_847),
.B(n_834),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_845),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_845),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_845),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_844),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_855),
.A2(n_827),
.B1(n_826),
.B2(n_833),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_850),
.Y(n_857)
);

OAI322xp33_ASAP7_75t_L g858 ( 
.A1(n_852),
.A2(n_844),
.A3(n_849),
.B1(n_848),
.B2(n_816),
.C1(n_819),
.C2(n_833),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_851),
.Y(n_859)
);

OAI221xp5_ASAP7_75t_L g860 ( 
.A1(n_853),
.A2(n_791),
.B1(n_812),
.B2(n_821),
.C(n_829),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_SL g861 ( 
.A1(n_860),
.A2(n_854),
.B1(n_855),
.B2(n_851),
.Y(n_861)
);

OAI21xp33_ASAP7_75t_SL g862 ( 
.A1(n_859),
.A2(n_854),
.B(n_835),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_857),
.Y(n_863)
);

OAI31xp33_ASAP7_75t_L g864 ( 
.A1(n_858),
.A2(n_812),
.A3(n_807),
.B(n_808),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_863),
.B(n_856),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_862),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_861),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_864),
.B(n_835),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_863),
.B(n_843),
.Y(n_869)
);

NAND4xp75_ASAP7_75t_L g870 ( 
.A(n_865),
.B(n_714),
.C(n_832),
.D(n_751),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_869),
.Y(n_871)
);

NAND4xp25_ASAP7_75t_L g872 ( 
.A(n_866),
.B(n_830),
.C(n_834),
.D(n_839),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_865),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_867),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_868),
.A2(n_724),
.B(n_809),
.C(n_808),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_865),
.B(n_726),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_865),
.B(n_840),
.Y(n_877)
);

AOI21xp33_ASAP7_75t_L g878 ( 
.A1(n_874),
.A2(n_777),
.B(n_806),
.Y(n_878)
);

OAI211xp5_ASAP7_75t_L g879 ( 
.A1(n_873),
.A2(n_871),
.B(n_876),
.C(n_877),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_872),
.Y(n_880)
);

AOI221x1_ASAP7_75t_L g881 ( 
.A1(n_875),
.A2(n_764),
.B1(n_784),
.B2(n_723),
.C(n_746),
.Y(n_881)
);

NAND2xp33_ASAP7_75t_R g882 ( 
.A(n_870),
.B(n_829),
.Y(n_882)
);

AOI32xp33_ASAP7_75t_L g883 ( 
.A1(n_874),
.A2(n_842),
.A3(n_839),
.B1(n_834),
.B2(n_841),
.Y(n_883)
);

AOI221xp5_ASAP7_75t_L g884 ( 
.A1(n_874),
.A2(n_807),
.B1(n_778),
.B2(n_820),
.C(n_839),
.Y(n_884)
);

AOI211xp5_ASAP7_75t_L g885 ( 
.A1(n_876),
.A2(n_842),
.B(n_840),
.C(n_822),
.Y(n_885)
);

NAND3xp33_ASAP7_75t_SL g886 ( 
.A(n_873),
.B(n_780),
.C(n_779),
.Y(n_886)
);

OAI21xp33_ASAP7_75t_SL g887 ( 
.A1(n_874),
.A2(n_832),
.B(n_789),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_879),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_R g889 ( 
.A(n_880),
.B(n_735),
.Y(n_889)
);

AOI221xp5_ASAP7_75t_L g890 ( 
.A1(n_878),
.A2(n_887),
.B1(n_886),
.B2(n_884),
.C(n_885),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_883),
.B(n_824),
.Y(n_891)
);

NOR2x1p5_ASAP7_75t_L g892 ( 
.A(n_882),
.B(n_804),
.Y(n_892)
);

OAI22xp33_ASAP7_75t_L g893 ( 
.A1(n_881),
.A2(n_806),
.B1(n_813),
.B2(n_818),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_880),
.Y(n_894)
);

XNOR2x2_ASAP7_75t_SL g895 ( 
.A(n_880),
.B(n_743),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_R g896 ( 
.A(n_880),
.B(n_746),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_888),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_894),
.B(n_804),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_889),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_895),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_892),
.B(n_797),
.Y(n_901)
);

OAI321xp33_ASAP7_75t_L g902 ( 
.A1(n_890),
.A2(n_782),
.A3(n_748),
.B1(n_801),
.B2(n_813),
.C(n_707),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_896),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_893),
.A2(n_769),
.B1(n_764),
.B2(n_781),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_897),
.Y(n_905)
);

OAI221xp5_ASAP7_75t_L g906 ( 
.A1(n_899),
.A2(n_891),
.B1(n_781),
.B2(n_727),
.C(n_698),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_L g907 ( 
.A(n_900),
.B(n_762),
.C(n_764),
.Y(n_907)
);

AND3x1_ASAP7_75t_L g908 ( 
.A(n_898),
.B(n_707),
.C(n_719),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_903),
.A2(n_776),
.B1(n_805),
.B2(n_798),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_SL g910 ( 
.A1(n_901),
.A2(n_734),
.B1(n_719),
.B2(n_769),
.Y(n_910)
);

NOR4xp25_ASAP7_75t_L g911 ( 
.A(n_902),
.B(n_801),
.C(n_823),
.D(n_794),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_L g912 ( 
.A(n_901),
.B(n_152),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_905),
.Y(n_913)
);

OAI221xp5_ASAP7_75t_L g914 ( 
.A1(n_907),
.A2(n_904),
.B1(n_800),
.B2(n_734),
.C(n_803),
.Y(n_914)
);

XNOR2xp5_ASAP7_75t_L g915 ( 
.A(n_912),
.B(n_756),
.Y(n_915)
);

XOR2xp5_ASAP7_75t_L g916 ( 
.A(n_908),
.B(n_153),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_909),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_913),
.Y(n_918)
);

AOI22x1_ASAP7_75t_L g919 ( 
.A1(n_916),
.A2(n_910),
.B1(n_911),
.B2(n_906),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_917),
.B(n_756),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_918),
.A2(n_915),
.B(n_914),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_919),
.A2(n_798),
.B1(n_800),
.B2(n_797),
.Y(n_922)
);

OR3x1_ASAP7_75t_L g923 ( 
.A(n_921),
.B(n_920),
.C(n_922),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_921),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_924),
.Y(n_925)
);

NOR2x1_ASAP7_75t_L g926 ( 
.A(n_923),
.B(n_776),
.Y(n_926)
);

AO22x2_ASAP7_75t_L g927 ( 
.A1(n_924),
.A2(n_798),
.B1(n_776),
.B2(n_762),
.Y(n_927)
);

AOI221xp5_ASAP7_75t_L g928 ( 
.A1(n_925),
.A2(n_797),
.B1(n_803),
.B2(n_722),
.C(n_162),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_926),
.A2(n_154),
.B1(n_156),
.B2(n_161),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_929),
.Y(n_930)
);

OAI221xp5_ASAP7_75t_R g931 ( 
.A1(n_930),
.A2(n_928),
.B1(n_927),
.B2(n_166),
.C(n_167),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_SL g932 ( 
.A1(n_931),
.A2(n_163),
.B1(n_164),
.B2(n_170),
.Y(n_932)
);


endmodule