module fake_jpeg_431_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_2),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_5),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_0),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_20),
.C(n_21),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g16 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_7),
.A2(n_4),
.B1(n_6),
.B2(n_3),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_18),
.B(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_10),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_20),
.B1(n_21),
.B2(n_15),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_21),
.B1(n_14),
.B2(n_22),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_21),
.B1(n_14),
.B2(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_41),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_29),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.C(n_27),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_47),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_46),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_12),
.C(n_9),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_39),
.B(n_40),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_11),
.B(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_50),
.B(n_14),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_53),
.B(n_54),
.Y(n_55)
);

NAND4xp25_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_11),
.C(n_3),
.D(n_9),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_55),
.B(n_49),
.Y(n_56)
);


endmodule