module fake_jpeg_11287_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_7),
.B(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_62),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_3),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_65),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_3),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_19),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_63),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_4),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_49),
.B1(n_41),
.B2(n_51),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_71),
.B1(n_77),
.B2(n_56),
.Y(n_83)
);

NOR4xp25_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_27),
.C(n_40),
.D(n_38),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_23),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_49),
.B1(n_41),
.B2(n_45),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_54),
.C(n_52),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_53),
.C(n_10),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_63),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_54),
.B1(n_52),
.B2(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_87),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_84),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_16),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_55),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_53),
.B1(n_6),
.B2(n_7),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_86),
.B1(n_11),
.B2(n_12),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_53),
.B1(n_6),
.B2(n_8),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_5),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_93),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_9),
.Y(n_92)
);

XNOR2x1_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_94),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_100),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_70),
.B(n_9),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_107),
.B(n_109),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_13),
.C(n_14),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_107),
.C(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_15),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_34),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_104),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_17),
.B(n_21),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_36),
.B(n_24),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_114),
.Y(n_120)
);

XNOR2x1_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_116),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_22),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_25),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_118),
.A2(n_119),
.B1(n_99),
.B2(n_101),
.Y(n_122)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_110),
.B1(n_97),
.B2(n_120),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_126),
.C(n_123),
.Y(n_128)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_105),
.B(n_113),
.C(n_112),
.D(n_111),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_127),
.A2(n_128),
.B(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_114),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_102),
.B1(n_104),
.B2(n_119),
.Y(n_131)
);

AOI211xp5_ASAP7_75t_SL g132 ( 
.A1(n_131),
.A2(n_29),
.B(n_30),
.C(n_32),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_33),
.Y(n_133)
);


endmodule