module real_jpeg_371_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_2),
.A2(n_21),
.B1(n_22),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_2),
.A2(n_24),
.B1(n_30),
.B2(n_63),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_35),
.B1(n_42),
.B2(n_63),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_4),
.A2(n_21),
.B1(n_22),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_4),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_4),
.A2(n_24),
.B1(n_30),
.B2(n_66),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_4),
.A2(n_35),
.B1(n_42),
.B2(n_66),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_5),
.B(n_70),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_5),
.A2(n_21),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_5),
.B(n_60),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_5),
.B(n_35),
.C(n_52),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_5),
.A2(n_24),
.B1(n_28),
.B2(n_30),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_5),
.B(n_38),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_5),
.B(n_56),
.Y(n_119)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_8),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_8),
.A2(n_24),
.B1(n_30),
.B2(n_41),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_9),
.A2(n_35),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_11),
.A2(n_35),
.B1(n_42),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_11),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_12),
.A2(n_24),
.B1(n_30),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_12),
.A2(n_35),
.B1(n_42),
.B2(n_49),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_90),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_88),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_79),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_17),
.B(n_79),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_57),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_32),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.A3(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_21),
.A2(n_22),
.B1(n_26),
.B2(n_31),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_21),
.A2(n_22),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_24),
.A2(n_30),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

AO22x2_ASAP7_75t_SL g60 ( 
.A1(n_24),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_24),
.B(n_105),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_28),
.A2(n_34),
.B1(n_38),
.B2(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_37),
.B1(n_39),
.B2(n_43),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_33),
.A2(n_37),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_34),
.A2(n_38),
.B1(n_44),
.B2(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_34),
.A2(n_38),
.B1(n_40),
.B2(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_34),
.A2(n_38),
.B1(n_117),
.B2(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_42),
.B1(n_52),
.B2(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_35),
.B(n_115),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_54),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_50),
.A2(n_56),
.B1(n_87),
.B2(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_50),
.A2(n_56),
.B1(n_94),
.B2(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_67),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_62),
.B1(n_64),
.B2(n_82),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_75),
.B2(n_78),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.C(n_84),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_84),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_100),
.B(n_130),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_98),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.C(n_96),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_95),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_111),
.B(n_129),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_109),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_123),
.B(n_128),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_118),
.B(n_122),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_120),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_127),
.Y(n_128)
);


endmodule