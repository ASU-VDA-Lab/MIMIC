module fake_jpeg_12670_n_517 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVxp33_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_56),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_23),
.B(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_18),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_68),
.Y(n_160)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_72),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_90),
.Y(n_124)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_34),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_28),
.B(n_15),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_99),
.Y(n_129)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_93),
.Y(n_103)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_25),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_56),
.B(n_28),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_108),
.B(n_119),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_65),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_113),
.B(n_118),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_50),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_92),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_58),
.B(n_21),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_74),
.A2(n_21),
.B(n_47),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_156),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_88),
.A2(n_44),
.B1(n_50),
.B2(n_38),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_132),
.A2(n_54),
.B1(n_86),
.B2(n_99),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_87),
.B(n_0),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_140),
.C(n_29),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_82),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_32),
.C(n_46),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_54),
.A2(n_47),
.B(n_26),
.Y(n_156)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_162),
.Y(n_247)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx3_ASAP7_75t_SL g248 ( 
.A(n_164),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_75),
.B1(n_57),
.B2(n_60),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_169),
.A2(n_207),
.B1(n_19),
.B2(n_1),
.Y(n_258)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_171),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_172),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_73),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_173),
.B(n_185),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_176),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_114),
.A2(n_102),
.B1(n_101),
.B2(n_96),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_178),
.A2(n_214),
.B1(n_120),
.B2(n_134),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_210),
.Y(n_224)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_181),
.Y(n_249)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_115),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_183),
.B(n_186),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_197),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_122),
.B(n_73),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_112),
.B(n_35),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_105),
.B(n_27),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_188),
.B(n_190),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_189),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_105),
.B(n_27),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_112),
.A2(n_81),
.B1(n_80),
.B2(n_67),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_194),
.A2(n_134),
.B1(n_110),
.B2(n_158),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_32),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_195),
.B(n_201),
.Y(n_259)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_144),
.Y(n_196)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_124),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_130),
.A2(n_38),
.B1(n_46),
.B2(n_53),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_198),
.A2(n_200),
.B1(n_209),
.B2(n_211),
.Y(n_227)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_35),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_126),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_204),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_106),
.B(n_29),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_206),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_143),
.A2(n_37),
.B1(n_26),
.B2(n_45),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_208),
.B(n_212),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_130),
.A2(n_99),
.B1(n_86),
.B2(n_45),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_131),
.A2(n_43),
.B1(n_37),
.B2(n_36),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_129),
.B(n_43),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_137),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_132),
.A2(n_36),
.B1(n_19),
.B2(n_15),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_153),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_215),
.A2(n_142),
.B1(n_155),
.B2(n_145),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_149),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_216),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_103),
.B(n_14),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_217),
.Y(n_228)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_103),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_218),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_221),
.B(n_167),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_163),
.B(n_133),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_222),
.B(n_210),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_223),
.A2(n_239),
.B1(n_245),
.B2(n_263),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_168),
.A2(n_116),
.B(n_127),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_229),
.A2(n_256),
.B(n_215),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_168),
.A2(n_157),
.B1(n_120),
.B2(n_148),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_243),
.A2(n_181),
.B1(n_196),
.B2(n_176),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_184),
.A2(n_121),
.B1(n_125),
.B2(n_152),
.Y(n_245)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_111),
.B(n_146),
.C(n_154),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_251),
.A2(n_264),
.B(n_198),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_180),
.B(n_155),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_209),
.Y(n_283)
);

AO22x1_ASAP7_75t_L g256 ( 
.A1(n_187),
.A2(n_111),
.B1(n_19),
.B2(n_2),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_258),
.A2(n_174),
.B1(n_172),
.B2(n_8),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_175),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_204),
.A2(n_3),
.B(n_5),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_266),
.B(n_274),
.Y(n_343)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_267),
.Y(n_315)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_270),
.A2(n_256),
.B(n_264),
.Y(n_319)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_272),
.Y(n_333)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_226),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_273),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_225),
.B(n_193),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_165),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_235),
.A2(n_202),
.B1(n_164),
.B2(n_177),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_277),
.Y(n_340)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_278),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_289),
.Y(n_308)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_280),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_228),
.B(n_162),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_281),
.B(n_296),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_235),
.A2(n_206),
.B1(n_205),
.B2(n_191),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_L g317 ( 
.A1(n_282),
.A2(n_293),
.B1(n_302),
.B2(n_256),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_242),
.Y(n_331)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_286),
.Y(n_328)
);

BUFx12f_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_285),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_255),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_287),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_288),
.A2(n_263),
.B(n_245),
.Y(n_324)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_294),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_223),
.A2(n_199),
.B1(n_212),
.B2(n_200),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_268),
.B1(n_248),
.B2(n_258),
.Y(n_310)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_226),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_292),
.Y(n_336)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_257),
.Y(n_294)
);

AO22x2_ASAP7_75t_L g295 ( 
.A1(n_229),
.A2(n_192),
.B1(n_189),
.B2(n_179),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_301),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_259),
.B(n_13),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_232),
.B(n_216),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_297),
.B(n_298),
.Y(n_330)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_237),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_299),
.B(n_300),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_233),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_234),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_236),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_303),
.B(n_305),
.Y(n_345)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_306),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_259),
.B(n_13),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_247),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_244),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_220),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_253),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_309),
.B(n_322),
.C(n_278),
.Y(n_355)
);

OA22x2_ASAP7_75t_L g369 ( 
.A1(n_310),
.A2(n_238),
.B1(n_261),
.B2(n_219),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_288),
.A2(n_227),
.B1(n_239),
.B2(n_222),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_312),
.A2(n_326),
.B1(n_335),
.B2(n_248),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_317),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_319),
.A2(n_273),
.B(n_166),
.Y(n_373)
);

OA21x2_ASAP7_75t_L g320 ( 
.A1(n_293),
.A2(n_251),
.B(n_224),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_320),
.B(n_326),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_268),
.A2(n_291),
.B1(n_224),
.B2(n_276),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_321),
.A2(n_246),
.B1(n_290),
.B2(n_249),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_279),
.B(n_224),
.C(n_221),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_324),
.A2(n_325),
.B(n_339),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_271),
.A2(n_244),
.B(n_231),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_270),
.A2(n_271),
.B1(n_295),
.B2(n_267),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_295),
.A2(n_233),
.B1(n_249),
.B2(n_234),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_327),
.A2(n_284),
.B1(n_269),
.B2(n_294),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_331),
.B(n_166),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_295),
.A2(n_248),
.B1(n_261),
.B2(n_238),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_295),
.A2(n_307),
.B(n_306),
.Y(n_339)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_344),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_346),
.A2(n_359),
.B1(n_362),
.B2(n_323),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_343),
.B(n_304),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_347),
.B(n_349),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_348),
.A2(n_321),
.B1(n_316),
.B2(n_324),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_343),
.B(n_240),
.Y(n_349)
);

INVx13_ASAP7_75t_L g350 ( 
.A(n_341),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_350),
.Y(n_401)
);

INVx13_ASAP7_75t_L g351 ( 
.A(n_341),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_351),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_345),
.B(n_231),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_352),
.B(n_353),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_334),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_332),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_356),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_357),
.C(n_367),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_332),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_280),
.C(n_299),
.Y(n_357)
);

OAI21xp33_ASAP7_75t_L g359 ( 
.A1(n_330),
.A2(n_298),
.B(n_301),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_314),
.B(n_289),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_360),
.B(n_365),
.Y(n_405)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_337),
.Y(n_363)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_363),
.Y(n_382)
);

NAND3xp33_ASAP7_75t_L g365 ( 
.A(n_313),
.B(n_334),
.C(n_330),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_331),
.B(n_220),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_315),
.Y(n_368)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_368),
.Y(n_387)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_370),
.B(n_328),
.Y(n_407)
);

AOI22x1_ASAP7_75t_L g403 ( 
.A1(n_371),
.A2(n_338),
.B1(n_328),
.B2(n_336),
.Y(n_403)
);

OA21x2_ASAP7_75t_L g372 ( 
.A1(n_316),
.A2(n_246),
.B(n_292),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_336),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_373),
.A2(n_377),
.B(n_325),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_313),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_378),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_SL g375 ( 
.A(n_322),
.B(n_241),
.C(n_272),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_375),
.B(n_320),
.C(n_344),
.Y(n_392)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_323),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_318),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_319),
.A2(n_286),
.B(n_285),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_308),
.Y(n_378)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_380),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_348),
.A2(n_339),
.B1(n_310),
.B2(n_312),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_396),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_308),
.Y(n_384)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_385),
.A2(n_408),
.B(n_361),
.Y(n_416)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_388),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_318),
.Y(n_389)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_389),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_320),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_390),
.B(n_373),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_392),
.B(n_398),
.C(n_370),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_393),
.A2(n_399),
.B1(n_362),
.B2(n_366),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_356),
.B(n_311),
.Y(n_394)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_394),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_358),
.B(n_329),
.Y(n_395)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_395),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_311),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_357),
.B(n_320),
.C(n_329),
.Y(n_398)
);

AOI22x1_ASAP7_75t_SL g399 ( 
.A1(n_364),
.A2(n_340),
.B1(n_335),
.B2(n_342),
.Y(n_399)
);

AND2x2_ASAP7_75t_SL g402 ( 
.A(n_364),
.B(n_342),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_403),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_407),
.B(n_372),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_367),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_409),
.B(n_412),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_379),
.C(n_375),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_415),
.C(n_425),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_377),
.C(n_361),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_416),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_418),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_384),
.A2(n_372),
.B1(n_376),
.B2(n_368),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_420),
.A2(n_424),
.B1(n_402),
.B2(n_408),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_346),
.C(n_338),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_404),
.B(n_333),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_426),
.Y(n_449)
);

XNOR2x1_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_383),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_380),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_389),
.B(n_328),
.Y(n_428)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_428),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_391),
.B(n_363),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_433),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_405),
.A2(n_369),
.B1(n_337),
.B2(n_350),
.Y(n_432)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_432),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_381),
.B(n_369),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_R g434 ( 
.A(n_411),
.B(n_406),
.Y(n_434)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_434),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_422),
.A2(n_393),
.B1(n_397),
.B2(n_384),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_435),
.B(n_447),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_438),
.B(n_446),
.Y(n_465)
);

AOI21x1_ASAP7_75t_L g440 ( 
.A1(n_431),
.A2(n_381),
.B(n_385),
.Y(n_440)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_440),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_429),
.A2(n_397),
.B1(n_399),
.B2(n_400),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_443),
.B(n_452),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_445),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_409),
.B(n_402),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_413),
.A2(n_388),
.B(n_401),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_403),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_448),
.B(n_454),
.C(n_416),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_422),
.A2(n_395),
.B1(n_394),
.B2(n_396),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_450),
.B(n_453),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_410),
.A2(n_403),
.B1(n_400),
.B2(n_401),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_412),
.B(n_387),
.C(n_386),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_387),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_458),
.B(n_448),
.Y(n_480)
);

OAI322xp33_ASAP7_75t_L g459 ( 
.A1(n_434),
.A2(n_428),
.A3(n_414),
.B1(n_423),
.B2(n_421),
.C1(n_431),
.C2(n_417),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_470),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_453),
.B(n_451),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_463),
.Y(n_473)
);

BUFx12_ASAP7_75t_L g463 ( 
.A(n_439),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_425),
.C(n_415),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_466),
.B(n_467),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_441),
.B(n_382),
.Y(n_467)
);

BUFx12_ASAP7_75t_L g468 ( 
.A(n_439),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_469),
.Y(n_484)
);

AOI322xp5_ASAP7_75t_SL g469 ( 
.A1(n_449),
.A2(n_436),
.A3(n_433),
.B1(n_421),
.B2(n_452),
.C1(n_420),
.C2(n_451),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_382),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_466),
.B(n_460),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_471),
.B(n_474),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_454),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_456),
.A2(n_442),
.B1(n_423),
.B2(n_419),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_475),
.A2(n_171),
.B1(n_6),
.B2(n_8),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_456),
.A2(n_445),
.B1(n_419),
.B2(n_386),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_476),
.A2(n_457),
.B1(n_462),
.B2(n_463),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_455),
.B(n_446),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_478),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_438),
.C(n_437),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_437),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_480),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_369),
.C(n_285),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_483),
.C(n_468),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_285),
.C(n_351),
.Y(n_483)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_486),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_462),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_491),
.Y(n_497)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_473),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_492),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_457),
.Y(n_491)
);

FAx1_ASAP7_75t_SL g492 ( 
.A(n_478),
.B(n_468),
.CI(n_463),
.CON(n_492),
.SN(n_492)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_493),
.B(n_171),
.C(n_6),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_494),
.B(n_493),
.C(n_482),
.Y(n_501)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_484),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_495),
.A2(n_481),
.B(n_472),
.Y(n_496)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_496),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_489),
.A2(n_471),
.B(n_483),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_500),
.B(n_501),
.C(n_502),
.Y(n_505)
);

AOI322xp5_ASAP7_75t_L g503 ( 
.A1(n_498),
.A2(n_492),
.A3(n_489),
.B1(n_491),
.B2(n_487),
.C1(n_485),
.C2(n_490),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_506),
.Y(n_509)
);

AOI322xp5_ASAP7_75t_L g506 ( 
.A1(n_499),
.A2(n_490),
.A3(n_6),
.B1(n_9),
.B2(n_10),
.C1(n_12),
.C2(n_5),
.Y(n_506)
);

AND2x4_ASAP7_75t_SL g507 ( 
.A(n_497),
.B(n_5),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_507),
.A2(n_502),
.B(n_9),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_504),
.B(n_497),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_508),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_510),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_511),
.B(n_509),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_505),
.C(n_512),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_514),
.A2(n_6),
.B(n_10),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_12),
.C(n_300),
.Y(n_516)
);

BUFx24_ASAP7_75t_SL g517 ( 
.A(n_516),
.Y(n_517)
);


endmodule