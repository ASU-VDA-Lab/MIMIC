module real_aes_2871_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_41;
wire n_34;
wire n_12;
wire n_19;
wire n_40;
wire n_25;
wire n_43;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
INVx1_ASAP7_75t_L g28 ( .A(n_0), .Y(n_28) );
NOR2xp33_ASAP7_75t_L g13 ( .A(n_1), .B(n_5), .Y(n_13) );
CKINVDCx16_ASAP7_75t_R g23 ( .A(n_2), .Y(n_23) );
INVx3_ASAP7_75t_L g26 ( .A(n_3), .Y(n_26) );
AOI221xp5_ASAP7_75t_SL g10 ( .A1(n_4), .A2(n_11), .B1(n_29), .B2(n_32), .C(n_38), .Y(n_10) );
INVx1_ASAP7_75t_L g40 ( .A(n_4), .Y(n_40) );
INVx1_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_6), .B(n_17), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_6), .B(n_20), .Y(n_19) );
NOR2xp33_ASAP7_75t_L g21 ( .A(n_6), .B(n_22), .Y(n_21) );
AND2x4_ASAP7_75t_L g45 ( .A(n_6), .B(n_28), .Y(n_45) );
BUFx2_ASAP7_75t_L g31 ( .A(n_7), .Y(n_31) );
INVx2_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
INVxp67_ASAP7_75t_L g20 ( .A(n_9), .Y(n_20) );
OAI21xp33_ASAP7_75t_SL g11 ( .A1(n_12), .A2(n_13), .B(n_14), .Y(n_11) );
CKINVDCx14_ASAP7_75t_R g37 ( .A(n_12), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_13), .B(n_40), .Y(n_39) );
NOR4xp25_ASAP7_75t_L g14 ( .A(n_15), .B(n_18), .C(n_21), .D(n_27), .Y(n_14) );
INVxp67_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
NOR2xp33_ASAP7_75t_L g43 ( .A(n_17), .B(n_20), .Y(n_43) );
INVx1_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
INVx1_ASAP7_75t_L g36 ( .A(n_22), .Y(n_36) );
NOR2xp33_ASAP7_75t_L g22 ( .A(n_23), .B(n_24), .Y(n_22) );
INVx2_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_26), .Y(n_25) );
INVx1_ASAP7_75t_L g34 ( .A(n_27), .Y(n_34) );
INVx1_ASAP7_75t_L g27 ( .A(n_28), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_30), .Y(n_29) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_31), .Y(n_30) );
CKINVDCx14_ASAP7_75t_R g32 ( .A(n_33), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_34), .B(n_35), .Y(n_33) );
NOR2xp33_ASAP7_75t_L g35 ( .A(n_36), .B(n_37), .Y(n_35) );
NOR2xp33_ASAP7_75t_L g38 ( .A(n_39), .B(n_41), .Y(n_38) );
OR2x2_ASAP7_75t_L g41 ( .A(n_42), .B(n_44), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_43), .Y(n_42) );
INVxp67_ASAP7_75t_L g44 ( .A(n_45), .Y(n_44) );
endmodule