module real_jpeg_25265_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_0),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_0),
.A2(n_36),
.B1(n_56),
.B2(n_57),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_0),
.A2(n_36),
.B1(n_68),
.B2(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_0),
.A2(n_22),
.B1(n_26),
.B2(n_36),
.Y(n_158)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_22),
.B1(n_26),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_2),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_2),
.A2(n_68),
.B1(n_70),
.B2(n_97),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_2),
.A2(n_30),
.B1(n_42),
.B2(n_97),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_2),
.A2(n_56),
.B1(n_57),
.B2(n_97),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_7),
.A2(n_22),
.B1(n_26),
.B2(n_87),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_7),
.A2(n_68),
.B1(n_70),
.B2(n_87),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_7),
.A2(n_56),
.B1(n_57),
.B2(n_87),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_8),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_8),
.A2(n_22),
.B1(n_26),
.B2(n_170),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_8),
.A2(n_68),
.B1(n_70),
.B2(n_170),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_8),
.A2(n_56),
.B1(n_57),
.B2(n_170),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_9),
.A2(n_31),
.B1(n_37),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_9),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_9),
.A2(n_22),
.B1(n_26),
.B2(n_119),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_9),
.A2(n_68),
.B1(n_70),
.B2(n_119),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_9),
.A2(n_56),
.B1(n_57),
.B2(n_119),
.Y(n_281)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_10),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_11),
.A2(n_33),
.B1(n_37),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_11),
.A2(n_22),
.B1(n_26),
.B2(n_83),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_11),
.A2(n_68),
.B1(n_70),
.B2(n_83),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_11),
.A2(n_56),
.B1(n_57),
.B2(n_83),
.Y(n_232)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_13),
.B(n_30),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_13),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_13),
.B(n_21),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_13),
.B(n_68),
.C(n_93),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_13),
.A2(n_22),
.B1(n_26),
.B2(n_223),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_13),
.B(n_134),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_13),
.A2(n_68),
.B1(n_70),
.B2(n_223),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_13),
.B(n_56),
.C(n_73),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_13),
.A2(n_55),
.B(n_282),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_14),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_14),
.A2(n_22),
.B1(n_26),
.B2(n_67),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_14),
.A2(n_33),
.B1(n_67),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_14),
.A2(n_56),
.B1(n_57),
.B2(n_67),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_15),
.A2(n_41),
.B1(n_68),
.B2(n_70),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_15),
.A2(n_41),
.B1(n_56),
.B2(n_57),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_15),
.A2(n_22),
.B1(n_26),
.B2(n_41),
.Y(n_136)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_16),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_16),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_47),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_45),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_28),
.B(n_35),
.Y(n_20)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_21),
.A2(n_28),
.B1(n_35),
.B2(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_21),
.A2(n_28),
.B1(n_118),
.B2(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_21),
.A2(n_28),
.B1(n_40),
.B2(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_22),
.A2(n_26),
.B1(n_93),
.B2(n_94),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_22),
.B(n_27),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_22),
.B(n_248),
.Y(n_247)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_27),
.B1(n_30),
.B2(n_33),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_24),
.A2(n_26),
.A3(n_31),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_28),
.B(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_28),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_28),
.A2(n_122),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_32),
.Y(n_154)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_33),
.A2(n_223),
.B(n_224),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_34),
.A2(n_82),
.B(n_84),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_34),
.B(n_86),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_34),
.A2(n_82),
.B1(n_120),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_34),
.A2(n_120),
.B1(n_142),
.B2(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_34),
.A2(n_84),
.B(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_39),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_39),
.B(n_357),
.Y(n_358)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_356),
.B(n_358),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_344),
.B(n_355),
.Y(n_48)
);

OAI31xp33_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_144),
.A3(n_160),
.B(n_341),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_123),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_51),
.B(n_123),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_88),
.C(n_104),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_52),
.A2(n_88),
.B1(n_89),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_52),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_78),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_53),
.A2(n_54),
.B(n_80),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_64),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_54),
.A2(n_64),
.B1(n_65),
.B2(n_79),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B(n_63),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_55),
.A2(n_60),
.B1(n_63),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_55),
.A2(n_109),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_55),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_55),
.A2(n_199),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_55),
.B(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_55),
.A2(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_57),
.B1(n_73),
.B2(n_74),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_57),
.B(n_307),
.Y(n_306)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_59),
.Y(n_180)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_59),
.Y(n_309)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_66),
.A2(n_71),
.B1(n_77),
.B2(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_SL g70 ( 
.A(n_68),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_70),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_68),
.B(n_289),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_71),
.A2(n_77),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_71),
.B(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_71),
.A2(n_77),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_75),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_75),
.A2(n_100),
.B1(n_113),
.B2(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_75),
.A2(n_182),
.B(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_75),
.A2(n_219),
.B(n_255),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_75),
.B(n_223),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_77),
.B(n_220),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_99),
.B(n_103),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_99),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_98),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_91),
.A2(n_92),
.B1(n_136),
.B2(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_91),
.A2(n_189),
.B(n_191),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_91),
.A2(n_191),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_92),
.A2(n_115),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_92),
.A2(n_173),
.B(n_228),
.Y(n_227)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_98),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_100),
.A2(n_269),
.B(n_270),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_100),
.A2(n_270),
.B(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_102),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_104),
.A2(n_105),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_114),
.C(n_116),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_106),
.A2(n_107),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_184),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_108),
.Y(n_184)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_114),
.B(n_116),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_120),
.B(n_121),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_126),
.C(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_141),
.B2(n_143),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_137),
.B1(n_138),
.B2(n_140),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_138),
.C(n_141),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_133),
.A2(n_134),
.B1(n_190),
.B2(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_133),
.A2(n_134),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_134),
.B(n_174),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_138),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_138),
.B(n_151),
.C(n_157),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_141),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_143),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_141),
.B(n_147),
.C(n_150),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_145),
.A2(n_342),
.B(n_343),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_159),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_146),
.B(n_159),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_152),
.Y(n_351)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_158),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_334),
.B(n_340),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_208),
.B(n_333),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_201),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_163),
.B(n_201),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_183),
.C(n_185),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_164),
.A2(n_165),
.B1(n_183),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_175),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_171),
.C(n_175),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_181),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_176),
.B(n_181),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_196)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_180),
.A2(n_250),
.B(n_251),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_183),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_185),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_192),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_188),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_192),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_196),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_197),
.A2(n_293),
.B1(n_295),
.B2(n_297),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_203),
.B(n_204),
.C(n_207),
.Y(n_339)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_240),
.B(n_327),
.C(n_332),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_234),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_234),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_225),
.C(n_226),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_211),
.A2(n_212),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_221),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_217),
.C(n_221),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_223),
.B(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_225),
.B(n_226),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_231),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_233),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_235),
.B(n_238),
.C(n_239),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_321),
.B(n_326),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_271),
.B(n_320),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_260),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_245),
.B(n_260),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.C(n_257),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_246),
.B(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_253),
.A2(n_257),
.B1(n_258),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_253),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_265),
.B2(n_266),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_261),
.B(n_267),
.C(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_314),
.B(n_319),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_290),
.B(n_313),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_284),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_284),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_280),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_276),
.B(n_279),
.C(n_280),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_300),
.B(n_312),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_298),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_298),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_296),
.B(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_305),
.B(n_311),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_303),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_310),
.Y(n_305)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_318),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_325),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_325),
.Y(n_326)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_339),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_339),
.Y(n_340)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_336),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_345),
.B(n_346),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_354),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_350),
.B1(n_352),
.B2(n_353),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_348),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_350),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_352),
.C(n_354),
.Y(n_357)
);


endmodule