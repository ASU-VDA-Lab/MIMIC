module real_jpeg_5321_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_0),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_0),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_0),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_0),
.B(n_79),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_0),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_0),
.B(n_147),
.Y(n_146)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_2),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_2),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_2),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_2),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_2),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_2),
.B(n_40),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_2),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_3),
.B(n_79),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_3),
.B(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_3),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_3),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_3),
.B(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_3),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_3),
.B(n_241),
.Y(n_449)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_4),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_4),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_4),
.Y(n_301)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_6),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_6),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_6),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_6),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_6),
.B(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_6),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_6),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_6),
.B(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_7),
.Y(n_147)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_7),
.Y(n_231)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_7),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_7),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_7),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_7),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_8),
.Y(n_508)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_9),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_9),
.Y(n_423)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_11),
.Y(n_505)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_12),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_12),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_13),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_13),
.B(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_13),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_13),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_13),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_13),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_13),
.B(n_363),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_13),
.A2(n_418),
.B(n_423),
.Y(n_422)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_14),
.Y(n_151)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_14),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_14),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_15),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_15),
.B(n_155),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_15),
.B(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_15),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_15),
.B(n_272),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_15),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_15),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_15),
.B(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_16),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_16),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_16),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_16),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_16),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_16),
.B(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_16),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_17),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_17),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_17),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_17),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_17),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_17),
.B(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_17),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_17),
.B(n_332),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_503),
.B(n_506),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_69),
.B(n_102),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_21),
.B(n_69),
.Y(n_102)
);

BUFx24_ASAP7_75t_SL g510 ( 
.A(n_21),
.Y(n_510)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_57),
.CI(n_58),
.CON(n_21),
.SN(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_42),
.C(n_46),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_23),
.A2(n_24),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_47),
.C(n_52),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_27),
.A2(n_28),
.B1(n_47),
.B2(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_27),
.A2(n_28),
.B1(n_458),
.B2(n_459),
.Y(n_457)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_28),
.B(n_33),
.C(n_39),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_28),
.B(n_226),
.C(n_232),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g374 ( 
.A(n_30),
.Y(n_374)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_32),
.Y(n_132)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_32),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_32),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_33),
.A2(n_34),
.B1(n_61),
.B2(n_65),
.Y(n_60)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_34),
.B(n_179),
.C(n_182),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_34),
.B(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g363 ( 
.A(n_36),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_37),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_38),
.A2(n_39),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_39),
.B(n_133),
.C(n_137),
.Y(n_161)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_46),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_66),
.C(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_47),
.A2(n_96),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_47),
.A2(n_96),
.B1(n_404),
.B2(n_408),
.Y(n_403)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_50),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_50),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_50),
.Y(n_340)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_51),
.Y(n_136)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_51),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_51),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_53),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_52),
.A2(n_53),
.B1(n_122),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_120),
.C(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_66),
.B2(n_68),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_61),
.B(n_190),
.C(n_194),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_61),
.A2(n_65),
.B1(n_154),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_61),
.A2(n_65),
.B1(n_194),
.B2(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_65),
.B(n_144),
.C(n_154),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_66),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_66),
.A2(n_68),
.B1(n_73),
.B2(n_74),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_97),
.C(n_98),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_70),
.B(n_501),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_83),
.C(n_93),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_71),
.B(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_78),
.C(n_81),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_73),
.A2(n_74),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_73),
.B(n_113),
.C(n_120),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_73),
.A2(n_74),
.B1(n_371),
.B2(n_375),
.Y(n_370)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_74),
.B(n_371),
.C(n_376),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_81),
.B2(n_82),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_77),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_83),
.B(n_93),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.C(n_90),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_84),
.A2(n_87),
.B1(n_88),
.B2(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_84),
.Y(n_141)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_86),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_87),
.A2(n_88),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_88),
.B(n_146),
.C(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_92),
.B(n_285),
.Y(n_417)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_96),
.B(n_397),
.C(n_408),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_97),
.B(n_98),
.Y(n_501)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AO21x1_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_498),
.B(n_502),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_247),
.B(n_495),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_202),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_SL g495 ( 
.A1(n_106),
.A2(n_496),
.B(n_497),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_168),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_107),
.B(n_168),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_159),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_108),
.B(n_160),
.C(n_166),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_139),
.C(n_142),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_109),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_121),
.C(n_126),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_110),
.B(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_119),
.B2(n_120),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_114),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_114),
.A2(n_120),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_114),
.A2(n_120),
.B1(n_226),
.B2(n_227),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_114),
.B(n_227),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_118),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_118),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_121),
.B(n_126),
.Y(n_207)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_128)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_131),
.Y(n_266)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_132),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_133),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_133),
.B(n_216),
.Y(n_442)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_138),
.B(n_215),
.C(n_217),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_144),
.A2(n_145),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_152),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_152),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_146),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_146),
.A2(n_185),
.B1(n_191),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_146),
.A2(n_185),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_146),
.B(n_281),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_148),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_148),
.A2(n_187),
.B1(n_426),
.B2(n_427),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_148),
.B(n_427),
.C(n_430),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_150),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_151),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_158),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_169),
.C(n_172),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_160),
.B(n_169),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.CI(n_163),
.CON(n_160),
.SN(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_172),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_189),
.C(n_198),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.C(n_183),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_174),
.B(n_178),
.Y(n_466)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_182),
.Y(n_223)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_183),
.B(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_198),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_191),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_191),
.A2(n_213),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_191),
.B(n_383),
.Y(n_411)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_194),
.Y(n_244)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_245),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_203),
.B(n_245),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.C(n_208),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_204),
.B(n_206),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_208),
.B(n_472),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_224),
.C(n_242),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g467 ( 
.A(n_209),
.B(n_468),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.C(n_222),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_210),
.B(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_214),
.B(n_222),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_217),
.B(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g468 ( 
.A(n_224),
.B(n_242),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_234),
.C(n_237),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_225),
.B(n_451),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_226),
.A2(n_227),
.B1(n_232),
.B2(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_231),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_232),
.Y(n_460)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_233),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_234),
.A2(n_237),
.B1(n_238),
.B2(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_234),
.Y(n_452)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI221xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_435),
.B1(n_488),
.B2(n_493),
.C(n_494),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_390),
.B(n_434),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_351),
.B(n_389),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_326),
.B(n_350),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_293),
.B(n_325),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_282),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_253),
.B(n_282),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_267),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_254),
.B(n_268),
.C(n_279),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_259),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_255),
.B(n_260),
.C(n_264),
.Y(n_336)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_279),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_274),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_274),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_270),
.B(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_273),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.C(n_289),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_283),
.B(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_284),
.A2(n_289),
.B1(n_290),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_319),
.B(n_324),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_309),
.B(n_318),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_306),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_306),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_302),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_302),
.Y(n_320)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_314),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_321),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_328),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_335),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_329),
.B(n_336),
.C(n_337),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_334),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_333),
.C(n_334),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_341),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_338),
.B(n_342),
.C(n_349),
.Y(n_385)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_345),
.B2(n_349),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_345),
.Y(n_349)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_388),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_352),
.B(n_388),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_368),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_354),
.B(n_357),
.C(n_368),
.Y(n_391)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_365),
.B1(n_366),
.B2(n_367),
.Y(n_357)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_358),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_362),
.B2(n_364),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_359),
.B(n_364),
.C(n_365),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_362),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_381),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_369),
.B(n_385),
.C(n_387),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_376),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_371),
.Y(n_375)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_385),
.B1(n_386),
.B2(n_387),
.Y(n_381)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_382),
.Y(n_387)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_385),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_392),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_414),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_394),
.B(n_395),
.C(n_414),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_409),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_396),
.B(n_410),
.C(n_413),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_403),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_404),
.Y(n_408)
);

INVx6_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_411),
.B1(n_412),
.B2(n_413),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_433),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_424),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_416),
.B(n_424),
.C(n_433),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_418),
.B(n_422),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_422),
.B(n_448),
.C(n_449),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_422),
.B(n_462),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_430),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

NOR3xp33_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_470),
.C(n_474),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_436),
.A2(n_489),
.B(n_492),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_463),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_437),
.B(n_463),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_453),
.C(n_455),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_438),
.B(n_453),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_446),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_447),
.C(n_450),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_443),
.C(n_444),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_441),
.B(n_445),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_443),
.B(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_450),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_448),
.B(n_449),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_483),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.C(n_461),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_456),
.B(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_461),
.Y(n_478)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_469),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_467),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_465),
.B(n_467),
.C(n_469),
.Y(n_473)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_470),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_473),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_484),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_475),
.A2(n_490),
.B(n_491),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_482),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_482),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_479),
.C(n_480),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_477),
.B(n_487),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_480),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_486),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_499),
.B(n_500),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g507 ( 
.A(n_504),
.Y(n_507)
);

INVx13_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);


endmodule