module fake_jpeg_30227_n_490 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_490);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_490;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_2),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_24),
.B(n_16),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_71),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_70),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_24),
.B(n_15),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_55),
.B(n_68),
.Y(n_108)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_63),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_28),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_27),
.B(n_15),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_27),
.B(n_1),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_83),
.Y(n_124)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_30),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_87),
.Y(n_126)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

BUFx4f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_1),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_18),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_85),
.A2(n_38),
.B1(n_47),
.B2(n_43),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_34),
.B(n_2),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_86),
.B(n_88),
.Y(n_158)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_18),
.B(n_25),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_34),
.B(n_5),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_89),
.B(n_97),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_40),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_45),
.Y(n_128)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_45),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_100),
.B(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_37),
.B(n_6),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_51),
.B1(n_49),
.B2(n_46),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_109),
.A2(n_119),
.B1(n_135),
.B2(n_136),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_64),
.A2(n_51),
.B1(n_49),
.B2(n_46),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_128),
.B(n_143),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_84),
.A2(n_20),
.B1(n_19),
.B2(n_46),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_132),
.A2(n_148),
.B1(n_50),
.B2(n_37),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_19),
.B1(n_20),
.B2(n_44),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_66),
.A2(n_49),
.B1(n_20),
.B2(n_36),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_137),
.A2(n_141),
.B1(n_156),
.B2(n_36),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_57),
.A2(n_99),
.B1(n_62),
.B2(n_69),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_85),
.A2(n_41),
.B1(n_33),
.B2(n_26),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_60),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_146),
.B(n_76),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_88),
.A2(n_50),
.B1(n_47),
.B2(n_43),
.Y(n_148)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_72),
.A2(n_32),
.B1(n_36),
.B2(n_41),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_77),
.B(n_38),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_159),
.B(n_33),
.Y(n_201)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_56),
.Y(n_160)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_165),
.Y(n_225)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_107),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_169),
.B(n_171),
.Y(n_226)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_88),
.Y(n_171)
);

BUFx2_ASAP7_75t_SL g172 ( 
.A(n_105),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_172),
.Y(n_251)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_124),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_204),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_106),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_176),
.B(n_182),
.Y(n_231)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_140),
.Y(n_180)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_180),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_60),
.C(n_70),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_181),
.B(n_122),
.C(n_113),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_108),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_183),
.A2(n_185),
.B1(n_188),
.B2(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_189),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_120),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_112),
.B(n_91),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_187),
.Y(n_241)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx11_ASAP7_75t_L g189 ( 
.A(n_134),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_190),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_114),
.B(n_87),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_191),
.B(n_197),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_96),
.B1(n_95),
.B2(n_90),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_133),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

BUFx12f_ASAP7_75t_SL g196 ( 
.A(n_108),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_196),
.A2(n_206),
.B1(n_209),
.B2(n_214),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_162),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_212),
.B1(n_135),
.B2(n_109),
.Y(n_216)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_200),
.B(n_201),
.Y(n_232)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_202),
.B(n_205),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_143),
.B(n_82),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_116),
.Y(n_205)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_97),
.B1(n_127),
.B2(n_138),
.Y(n_242)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_115),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_211),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_59),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_126),
.Y(n_236)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_143),
.A2(n_79),
.B1(n_90),
.B2(n_80),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_137),
.A2(n_81),
.B1(n_75),
.B2(n_32),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_132),
.A2(n_80),
.B1(n_91),
.B2(n_87),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_215),
.A2(n_210),
.B(n_196),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_216),
.A2(n_221),
.B1(n_222),
.B2(n_229),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_204),
.A2(n_198),
.B1(n_199),
.B2(n_177),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_119),
.B1(n_149),
.B2(n_130),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_199),
.A2(n_141),
.B1(n_131),
.B2(n_149),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_230),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_175),
.A2(n_121),
.B1(n_127),
.B2(n_130),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_233),
.A2(n_246),
.B1(n_180),
.B2(n_176),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_237),
.B(n_193),
.C(n_202),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_181),
.B(n_117),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_249),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_252),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_138),
.B1(n_123),
.B2(n_145),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_211),
.A2(n_139),
.B1(n_153),
.B2(n_42),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_166),
.A2(n_150),
.B1(n_144),
.B2(n_116),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_144),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_179),
.A2(n_42),
.B1(n_129),
.B2(n_98),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_170),
.B(n_150),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_238),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_223),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_262),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_260),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_178),
.Y(n_260)
);

OAI32xp33_ASAP7_75t_L g262 ( 
.A1(n_220),
.A2(n_173),
.A3(n_208),
.B1(n_213),
.B2(n_195),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_263),
.A2(n_267),
.B1(n_277),
.B2(n_279),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_248),
.A2(n_190),
.B1(n_188),
.B2(n_180),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_223),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_265),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_254),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_266),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_221),
.A2(n_213),
.B1(n_167),
.B2(n_203),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_217),
.Y(n_268)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_225),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_174),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_273),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_231),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_271),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g272 ( 
.A(n_220),
.B(n_167),
.CI(n_203),
.CON(n_272),
.SN(n_272)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_272),
.B(n_284),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_195),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_237),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_275),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_222),
.B(n_249),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_236),
.C(n_247),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_216),
.A2(n_229),
.B1(n_233),
.B2(n_242),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_217),
.Y(n_278)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_278),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_231),
.A2(n_209),
.B1(n_165),
.B2(n_183),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_200),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_283),
.Y(n_304)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_224),
.Y(n_282)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_232),
.B(n_184),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_232),
.B(n_168),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_250),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_224),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_286),
.B(n_245),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_235),
.A2(n_185),
.B1(n_194),
.B2(n_189),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_288),
.A2(n_228),
.B1(n_244),
.B2(n_252),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_235),
.B(n_241),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_291),
.A2(n_315),
.B(n_292),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_292),
.B(n_309),
.Y(n_322)
);

XOR2x2_ASAP7_75t_SL g293 ( 
.A(n_281),
.B(n_272),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_293),
.B(n_313),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_246),
.B1(n_230),
.B2(n_245),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_308),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_256),
.A2(n_277),
.B1(n_265),
.B2(n_257),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_234),
.B1(n_243),
.B2(n_247),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_300),
.B(n_261),
.C(n_283),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_234),
.B1(n_219),
.B2(n_236),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_250),
.B1(n_227),
.B2(n_225),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_310),
.A2(n_311),
.B1(n_279),
.B2(n_280),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_256),
.A2(n_267),
.B1(n_274),
.B2(n_263),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_271),
.A2(n_228),
.B(n_251),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_258),
.A2(n_228),
.B1(n_227),
.B2(n_225),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_318),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_258),
.A2(n_218),
.B1(n_239),
.B2(n_253),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_276),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_336),
.C(n_346),
.Y(n_356)
);

OAI21xp33_ASAP7_75t_SL g320 ( 
.A1(n_290),
.A2(n_259),
.B(n_285),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_320),
.A2(n_332),
.B1(n_206),
.B2(n_42),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_302),
.A2(n_261),
.B(n_270),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_321),
.A2(n_307),
.B(n_309),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_291),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_323),
.B(n_262),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_289),
.B(n_260),
.Y(n_324)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_290),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_326),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_297),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_331),
.Y(n_349)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_329),
.Y(n_351)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_306),
.Y(n_330)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_330),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_314),
.B(n_266),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_306),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_339),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_301),
.A2(n_303),
.B(n_302),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_335),
.A2(n_298),
.B(n_311),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_337),
.B(n_344),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_272),
.Y(n_338)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_272),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_289),
.B(n_273),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_340),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_268),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_341),
.A2(n_343),
.B1(n_345),
.B2(n_317),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_299),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_342),
.Y(n_369)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_293),
.B(n_282),
.C(n_278),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_293),
.B(n_288),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_299),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_347),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_295),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_348),
.B(n_358),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_335),
.A2(n_298),
.B(n_308),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_354),
.B(n_367),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_336),
.Y(n_358)
);

NOR3xp33_ASAP7_75t_SL g359 ( 
.A(n_331),
.B(n_304),
.C(n_317),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_359),
.B(n_326),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_322),
.A2(n_294),
.B1(n_310),
.B2(n_296),
.Y(n_360)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_361),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_344),
.C(n_313),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_365),
.C(n_373),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_322),
.A2(n_304),
.B1(n_315),
.B2(n_307),
.Y(n_364)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_364),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_316),
.C(n_318),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_368),
.B(n_376),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_339),
.A2(n_286),
.B1(n_269),
.B2(n_251),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_370),
.A2(n_374),
.B1(n_333),
.B2(n_334),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_321),
.A2(n_218),
.B(n_269),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_342),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_337),
.B(n_239),
.C(n_129),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_161),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_377),
.A2(n_350),
.B1(n_375),
.B2(n_359),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_366),
.A2(n_338),
.B1(n_333),
.B2(n_325),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_378),
.A2(n_384),
.B1(n_388),
.B2(n_360),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_341),
.Y(n_381)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_381),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_328),
.Y(n_382)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_382),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_325),
.C(n_332),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_356),
.C(n_358),
.Y(n_412)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_387),
.Y(n_409)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_351),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_366),
.A2(n_345),
.B1(n_343),
.B2(n_330),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_352),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_390),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_372),
.B(n_329),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_352),
.Y(n_391)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_391),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_392),
.Y(n_402)
);

XOR2x2_ASAP7_75t_L g395 ( 
.A(n_348),
.B(n_347),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_395),
.B(n_376),
.Y(n_407)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_397),
.Y(n_405)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_357),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_399),
.B(n_401),
.Y(n_403)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_367),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_401),
.B(n_373),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_382),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_412),
.Y(n_425)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_410),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_393),
.B(n_365),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_420),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_386),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_415),
.B(n_369),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_371),
.C(n_362),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_416),
.B(n_417),
.C(n_400),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_383),
.B(n_368),
.C(n_355),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_379),
.A2(n_374),
.B(n_354),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_418),
.A2(n_406),
.B(n_421),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_355),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_419),
.B(n_421),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_353),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_422),
.B(n_363),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_423),
.B(n_428),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_402),
.A2(n_396),
.B1(n_380),
.B2(n_394),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_424),
.A2(n_405),
.B1(n_408),
.B2(n_369),
.Y(n_446)
);

O2A1O1Ixp33_ASAP7_75t_SL g426 ( 
.A1(n_403),
.A2(n_398),
.B(n_381),
.C(n_378),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_426),
.A2(n_437),
.B(n_418),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_385),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_398),
.C(n_400),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_438),
.C(n_419),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_407),
.B(n_380),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_432),
.B(n_433),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_416),
.Y(n_433)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_434),
.Y(n_439)
);

OA21x2_ASAP7_75t_SL g435 ( 
.A1(n_411),
.A2(n_399),
.B(n_397),
.Y(n_435)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_435),
.Y(n_442)
);

AOI21xp33_ASAP7_75t_L g436 ( 
.A1(n_409),
.A2(n_391),
.B(n_389),
.Y(n_436)
);

NOR3xp33_ASAP7_75t_L g445 ( 
.A(n_436),
.B(n_404),
.C(n_414),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_388),
.C(n_387),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_441),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_446),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_415),
.Y(n_444)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_444),
.Y(n_456)
);

AOI21xp33_ASAP7_75t_L g459 ( 
.A1(n_445),
.A2(n_432),
.B(n_427),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_447),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_428),
.B(n_438),
.C(n_425),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_448),
.B(n_453),
.C(n_427),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_426),
.A2(n_363),
.B1(n_8),
.B2(n_9),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_449),
.A2(n_63),
.B1(n_8),
.B2(n_9),
.Y(n_460)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_431),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_450),
.B(n_452),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_6),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_430),
.C(n_423),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g457 ( 
.A(n_441),
.B(n_442),
.Y(n_457)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_457),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_458),
.B(n_461),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_459),
.A2(n_460),
.B1(n_9),
.B2(n_10),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_22),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_444),
.A2(n_6),
.B(n_8),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_462),
.B(n_449),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_439),
.A2(n_9),
.B(n_10),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_462),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_451),
.B(n_22),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_443),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_468),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_465),
.B(n_448),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_473),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_455),
.B(n_453),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_470),
.B(n_465),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_471),
.B(n_475),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_440),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_474),
.A2(n_455),
.B1(n_464),
.B2(n_463),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_479),
.B(n_480),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_472),
.B(n_454),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_481),
.A2(n_469),
.B(n_475),
.Y(n_483)
);

OAI31xp33_ASAP7_75t_SL g487 ( 
.A1(n_483),
.A2(n_485),
.A3(n_10),
.B(n_12),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_478),
.B(n_467),
.C(n_456),
.Y(n_484)
);

O2A1O1Ixp33_ASAP7_75t_SL g486 ( 
.A1(n_484),
.A2(n_476),
.B(n_477),
.C(n_13),
.Y(n_486)
);

OAI311xp33_ASAP7_75t_L g485 ( 
.A1(n_478),
.A2(n_460),
.A3(n_12),
.B1(n_13),
.C1(n_14),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_486),
.B(n_487),
.C(n_482),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_488),
.B(n_12),
.C(n_14),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_489),
.A2(n_22),
.B(n_476),
.Y(n_490)
);


endmodule