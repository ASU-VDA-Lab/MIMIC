module real_jpeg_16935_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_16),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_0),
.B(n_17),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_26),
.Y(n_25)
);

AND2x4_ASAP7_75t_SL g29 ( 
.A(n_1),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

NAND2x1p5_ASAP7_75t_L g66 ( 
.A(n_1),
.B(n_46),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_1),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_1),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_1),
.B(n_60),
.Y(n_100)
);

AND2x4_ASAP7_75t_L g127 ( 
.A(n_1),
.B(n_128),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_2),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_3),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_3),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_4),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_4),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_4),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_4),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_4),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_4),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_4),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_4),
.B(n_236),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_5),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_5),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_6),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_6),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_6),
.B(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_6),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_6),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_6),
.B(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_7),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_9),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_9),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_9),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_9),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g277 ( 
.A(n_9),
.B(n_278),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_9),
.B(n_283),
.Y(n_282)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_11),
.Y(n_96)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g140 ( 
.A(n_12),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_13),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_71),
.B(n_219),
.C(n_326),
.D(n_343),
.Y(n_17)
);

NOR3xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_174),
.C(n_198),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_150),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_20),
.B(n_150),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_89),
.C(n_114),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_21),
.B(n_90),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_61),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_22),
.B(n_62),
.C(n_72),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_47),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_23),
.B(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_23)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B(n_31),
.Y(n_24)
);

NAND2x1p5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_29),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_25),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_25),
.A2(n_64),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_25),
.B(n_93),
.C(n_99),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_25),
.A2(n_64),
.B1(n_141),
.B2(n_232),
.Y(n_316)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_29),
.A2(n_41),
.B(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_32),
.C(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_29),
.A2(n_41),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_29),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_31),
.B(n_32),
.C(n_248),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_32),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_32),
.A2(n_38),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_32),
.A2(n_38),
.B1(n_67),
.B2(n_68),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_36),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_36),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_38),
.B(n_75),
.C(n_106),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_SL g343 ( 
.A(n_38),
.B(n_68),
.C(n_211),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_39),
.B(n_47),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_40),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_41),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_41),
.B(n_79),
.C(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_41),
.A2(n_79),
.B1(n_120),
.B2(n_134),
.Y(n_272)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XNOR2x1_ASAP7_75t_L g117 ( 
.A(n_45),
.B(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_45),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_45),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_45),
.A2(n_211),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_46),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_57),
.Y(n_47)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_49),
.A2(n_50),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_49),
.A2(n_50),
.B1(n_99),
.B2(n_100),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_50),
.B(n_52),
.C(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_50),
.B(n_66),
.C(n_158),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_50),
.A2(n_100),
.B(n_277),
.C(n_281),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_51),
.Y(n_244)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_57),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_57),
.A2(n_113),
.B1(n_247),
.B2(n_248),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_94),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_58),
.B(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_72),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_63),
.B(n_66),
.C(n_68),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_66),
.A2(n_71),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_66),
.B(n_100),
.C(n_127),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_66),
.A2(n_71),
.B1(n_172),
.B2(n_173),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_73),
.C(n_86),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_67),
.A2(n_68),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_67),
.A2(n_68),
.B1(n_144),
.B2(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_68),
.B(n_136),
.C(n_144),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_68),
.B(n_86),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_68),
.B(n_75),
.C(n_242),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_68),
.B(n_124),
.C(n_133),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_73),
.A2(n_74),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.C(n_83),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_75),
.Y(n_105)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_79),
.A2(n_83),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AO21x1_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_122),
.B(n_130),
.Y(n_121)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_83),
.A2(n_126),
.B1(n_127),
.B2(n_133),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_83),
.B(n_123),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_86),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_137),
.C(n_141),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_101),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_91),
.B(n_102),
.C(n_112),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_97),
.B2(n_98),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_92),
.A2(n_93),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_93),
.B(n_182),
.C(n_185),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_93),
.B(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_93),
.A2(n_234),
.B(n_235),
.Y(n_303)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_95),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_99),
.B(n_127),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_99),
.A2(n_122),
.B(n_130),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_112),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_113),
.B(n_246),
.C(n_247),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_114),
.B(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_135),
.C(n_146),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_115),
.B(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.C(n_131),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_121),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_123),
.A2(n_124),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_127),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_126),
.A2(n_127),
.B1(n_215),
.B2(n_216),
.Y(n_287)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_127),
.B(n_133),
.C(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_127),
.B(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2x2_ASAP7_75t_L g288 ( 
.A(n_131),
.B(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_135),
.A2(n_146),
.B1(n_147),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_135),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_136),
.B(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_137),
.A2(n_141),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_137),
.Y(n_231)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_141),
.Y(n_232)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_144),
.Y(n_255)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_153),
.C(n_165),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_165),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_164),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_163),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_163),
.C(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_171),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_170),
.C(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_175),
.A2(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_197),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_176),
.B(n_197),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_196),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_196),
.C(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_190),
.B1(n_191),
.B2(n_195),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_194),
.C(n_195),
.Y(n_218)
);

OAI211xp5_ASAP7_75t_L g326 ( 
.A1(n_198),
.A2(n_327),
.B(n_330),
.C(n_331),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NAND2x1_ASAP7_75t_SL g330 ( 
.A(n_199),
.B(n_201),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_218),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_217),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_203),
.B(n_217),
.C(n_218),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_213),
.B2(n_214),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_205)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_334)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_215),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_260),
.B(n_325),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_258),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_222),
.B(n_258),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.C(n_256),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_256),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_245),
.C(n_252),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.C(n_241),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_229),
.B(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_233),
.A2(n_234),
.B1(n_241),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_241),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_242),
.A2(n_243),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_252),
.B1(n_253),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

XNOR2x2_ASAP7_75t_L g284 ( 
.A(n_246),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

AOI31xp67_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_291),
.A3(n_323),
.B(n_324),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_262),
.B(n_264),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.C(n_288),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_265),
.A2(n_266),
.B1(n_288),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_284),
.C(n_286),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.C(n_275),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_271),
.B(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_276),
.Y(n_320)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_277),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_286),
.B1(n_287),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_307),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_304),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_304),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.C(n_300),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_322),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_300),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.C(n_303),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_303),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_321),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.C(n_319),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.C(n_317),
.Y(n_311)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_341),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_342),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_340),
.B2(n_341),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_340),
.Y(n_341)
);


endmodule