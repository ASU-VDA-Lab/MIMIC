module fake_netlist_6_1275_n_1800 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1800);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1800;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_79),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_93),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_6),
.Y(n_174)
);

BUFx10_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_14),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_113),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_110),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_70),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_21),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_116),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_46),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_123),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_33),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_62),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_74),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_122),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_80),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_17),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_85),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_139),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_33),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_138),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_48),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_75),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_111),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_86),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_40),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_36),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_28),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_24),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_169),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_42),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_92),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_130),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_160),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_144),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_126),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_95),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_26),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_142),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_106),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_56),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_5),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_82),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_100),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_46),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_99),
.Y(n_230)
);

INVxp33_ASAP7_75t_SL g231 ( 
.A(n_148),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_6),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_65),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_149),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_112),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_66),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_4),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_60),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_119),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_16),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_8),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_103),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_81),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_21),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_23),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_146),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_38),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_3),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_97),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_167),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_159),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_41),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_109),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_11),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_56),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_28),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_162),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_24),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_87),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_150),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_152),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_83),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_76),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_101),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_22),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_0),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_43),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_63),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_37),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_105),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_120),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_131),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_90),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_17),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_32),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_31),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_78),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_11),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_132),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_25),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_32),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_145),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_36),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_41),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_38),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_64),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_115),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_102),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_57),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_5),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_40),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_73),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_89),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_161),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_30),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_88),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_67),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_27),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_134),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_20),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_50),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_15),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_54),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_158),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_117),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_94),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_72),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_170),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_133),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_61),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_137),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_20),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_107),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_0),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_3),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_59),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_57),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_77),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_127),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_22),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_27),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_42),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_8),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_128),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_23),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_13),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_19),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_18),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_155),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_9),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_53),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_135),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_25),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_154),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_71),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_52),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_98),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_143),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_13),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_69),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_118),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_26),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_12),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_52),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_91),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_129),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_15),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_68),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_241),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_241),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_331),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_241),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_241),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_241),
.B(n_299),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_314),
.B(n_1),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_207),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_231),
.B(n_1),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_208),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_241),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_241),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_241),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_248),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_314),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_224),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_178),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_187),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_299),
.B(n_2),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_172),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_196),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_226),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_196),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_282),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_221),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_232),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_237),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_187),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_305),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_316),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_221),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_281),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_340),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_240),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_281),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_245),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_247),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_181),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_303),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_252),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_209),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_231),
.B(n_2),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_255),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_256),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_258),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_209),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_209),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_197),
.B(n_4),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_197),
.B(n_7),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_261),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_265),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_278),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_209),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_300),
.B(n_7),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_209),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_174),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_266),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_177),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_263),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_215),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_267),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_232),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_232),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_269),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_189),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_184),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_210),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_274),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_205),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_206),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_212),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_216),
.Y(n_421)
);

NOR2xp67_ASAP7_75t_L g422 ( 
.A(n_300),
.B(n_9),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_229),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_193),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_219),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_222),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_193),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_275),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_244),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_290),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_276),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_295),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_280),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_223),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_227),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_284),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_298),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_285),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_225),
.B(n_10),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_233),
.Y(n_440)
);

INVx6_ASAP7_75t_L g441 ( 
.A(n_399),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_399),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_399),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_359),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_390),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_395),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_351),
.B(n_194),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_396),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_364),
.B(n_272),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_402),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_355),
.B(n_272),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_359),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_349),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_418),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_350),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_419),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_352),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_420),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_399),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_399),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_363),
.B(n_319),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_421),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_351),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_353),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_360),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_367),
.B(n_201),
.Y(n_467)
);

BUFx10_ASAP7_75t_L g468 ( 
.A(n_356),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_425),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_361),
.Y(n_470)
);

OAI21x1_ASAP7_75t_L g471 ( 
.A1(n_354),
.A2(n_296),
.B(n_225),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_405),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_377),
.B(n_173),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_407),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_424),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_414),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_R g477 ( 
.A(n_409),
.B(n_234),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_426),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_369),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_414),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_415),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_416),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_423),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_429),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_401),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_427),
.B(n_173),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_434),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_424),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_430),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_403),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_L g491 ( 
.A(n_356),
.B(n_186),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_432),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_370),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_435),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_437),
.Y(n_495)
);

AND3x1_ASAP7_75t_L g496 ( 
.A(n_357),
.B(n_254),
.C(n_201),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_440),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_372),
.B(n_254),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_374),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_380),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_358),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_381),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_384),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_398),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_368),
.B(n_319),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_397),
.B(n_179),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_358),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_388),
.B(n_296),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g509 ( 
.A(n_365),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_422),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_439),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_391),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_412),
.B(n_313),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_373),
.Y(n_514)
);

INVx6_ASAP7_75t_L g515 ( 
.A(n_366),
.Y(n_515)
);

OA21x2_ASAP7_75t_L g516 ( 
.A1(n_362),
.A2(n_322),
.B(n_283),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_442),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_444),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_442),
.Y(n_519)
);

AND2x2_ASAP7_75t_SL g520 ( 
.A(n_496),
.B(n_313),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_512),
.B(n_365),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_504),
.B(n_371),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_454),
.Y(n_523)
);

AND2x6_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_504),
.Y(n_524)
);

AND2x6_ASAP7_75t_L g525 ( 
.A(n_512),
.B(n_348),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_442),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_467),
.B(n_412),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_444),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_512),
.B(n_371),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_444),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_454),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_480),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_453),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_479),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_442),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_456),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_453),
.Y(n_537)
);

BUFx10_ASAP7_75t_L g538 ( 
.A(n_447),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_511),
.A2(n_283),
.B1(n_322),
.B2(n_339),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_458),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_458),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_512),
.B(n_376),
.Y(n_542)
);

AND2x6_ASAP7_75t_L g543 ( 
.A(n_504),
.B(n_348),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_512),
.B(n_376),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_480),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_480),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_480),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_465),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_515),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_465),
.Y(n_550)
);

CKINVDCx6p67_ASAP7_75t_R g551 ( 
.A(n_468),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_453),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_485),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_477),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_466),
.Y(n_555)
);

INVx5_ASAP7_75t_L g556 ( 
.A(n_480),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_485),
.B(n_383),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_504),
.B(n_383),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_490),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_490),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_467),
.B(n_385),
.Y(n_561)
);

INVx5_ASAP7_75t_L g562 ( 
.A(n_480),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_510),
.B(n_385),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_510),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_476),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_509),
.B(n_387),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_475),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_449),
.B(n_386),
.Y(n_568)
);

INVx6_ASAP7_75t_L g569 ( 
.A(n_504),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_476),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_442),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_504),
.B(n_488),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_506),
.B(n_473),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_475),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_468),
.B(n_386),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_511),
.A2(n_339),
.B1(n_320),
.B2(n_317),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_476),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_476),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_442),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_468),
.B(n_389),
.Y(n_580)
);

NOR2x1p5_ASAP7_75t_L g581 ( 
.A(n_493),
.B(n_186),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_445),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_466),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_468),
.B(n_389),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_443),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_445),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_443),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_470),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_506),
.B(n_392),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_481),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_515),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_481),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_488),
.B(n_392),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_473),
.B(n_393),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_488),
.B(n_176),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_449),
.B(n_393),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_449),
.B(n_394),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_446),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_443),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_505),
.B(n_394),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_481),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_481),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_443),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_446),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_448),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_496),
.A2(n_408),
.B1(n_436),
.B2(n_433),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_448),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_486),
.B(n_400),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_505),
.B(n_400),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_486),
.B(n_406),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_450),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_516),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_491),
.B(n_406),
.Y(n_613)
);

OR2x2_ASAP7_75t_SL g614 ( 
.A(n_515),
.B(n_326),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_516),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_443),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_443),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_505),
.B(n_410),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_516),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_505),
.B(n_410),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_515),
.B(n_343),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_508),
.B(n_413),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_516),
.A2(n_261),
.B1(n_211),
.B2(n_217),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_501),
.B(n_413),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_460),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_462),
.B(n_192),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_441),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_507),
.B(n_417),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_441),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_516),
.A2(n_261),
.B1(n_286),
.B2(n_277),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_513),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_450),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_493),
.B(n_417),
.Y(n_633)
);

AND2x2_ASAP7_75t_SL g634 ( 
.A(n_513),
.B(n_261),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_452),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_513),
.B(n_375),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_460),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_460),
.Y(n_638)
);

INVx4_ASAP7_75t_SL g639 ( 
.A(n_441),
.Y(n_639)
);

INVxp33_ASAP7_75t_L g640 ( 
.A(n_498),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_451),
.B(n_428),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_441),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_499),
.B(n_428),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_515),
.A2(n_438),
.B1(n_436),
.B2(n_433),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_514),
.Y(n_645)
);

INVxp33_ASAP7_75t_L g646 ( 
.A(n_498),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_452),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_499),
.B(n_431),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_SL g649 ( 
.A(n_513),
.B(n_190),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_462),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_SL g651 ( 
.A1(n_464),
.A2(n_379),
.B1(n_378),
.B2(n_382),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_483),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_441),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_461),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_461),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_483),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_461),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_483),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_508),
.B(n_431),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_508),
.B(n_438),
.Y(n_660)
);

BUFx6f_ASAP7_75t_SL g661 ( 
.A(n_451),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_484),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_484),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_484),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_492),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_492),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_573),
.B(n_451),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_589),
.B(n_451),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_542),
.A2(n_464),
.B1(n_462),
.B2(n_243),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_553),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_594),
.B(n_455),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_633),
.B(n_648),
.C(n_643),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_650),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_608),
.B(n_462),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_534),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_559),
.B(n_500),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_572),
.A2(n_471),
.B(n_500),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_650),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_522),
.A2(n_471),
.B(n_502),
.Y(n_679)
);

O2A1O1Ixp5_ASAP7_75t_L g680 ( 
.A1(n_619),
.A2(n_287),
.B(n_199),
.C(n_214),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_567),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_558),
.B(n_457),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_559),
.B(n_503),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_564),
.B(n_213),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_607),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_524),
.B(n_471),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_520),
.A2(n_342),
.B1(n_189),
.B2(n_259),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_524),
.B(n_218),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_520),
.A2(n_189),
.B1(n_250),
.B2(n_338),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_568),
.B(n_459),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_619),
.A2(n_189),
.B1(n_238),
.B2(n_260),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_619),
.A2(n_230),
.B(n_228),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_521),
.B(n_529),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_568),
.B(n_411),
.C(n_472),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_634),
.B(n_523),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_596),
.A2(n_597),
.B1(n_544),
.B2(n_600),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_596),
.B(n_463),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_634),
.B(n_235),
.Y(n_698)
);

BUFx4_ASAP7_75t_L g699 ( 
.A(n_534),
.Y(n_699)
);

INVx8_ASAP7_75t_L g700 ( 
.A(n_661),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_523),
.B(n_257),
.Y(n_701)
);

AOI221xp5_ASAP7_75t_L g702 ( 
.A1(n_576),
.A2(n_312),
.B1(n_203),
.B2(n_301),
.C(n_302),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_612),
.A2(n_189),
.B1(n_271),
.B2(n_324),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_615),
.A2(n_189),
.B1(n_304),
.B2(n_270),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_610),
.B(n_469),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_531),
.B(n_492),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_531),
.B(n_495),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_565),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_560),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_607),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_615),
.A2(n_189),
.B1(n_301),
.B2(n_312),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_635),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_565),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_569),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_536),
.B(n_495),
.Y(n_715)
);

BUFx2_ASAP7_75t_SL g716 ( 
.A(n_549),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_635),
.Y(n_717)
);

INVx4_ASAP7_75t_L g718 ( 
.A(n_567),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_647),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_538),
.B(n_478),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_647),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_631),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_570),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_538),
.B(n_487),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_540),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_597),
.B(n_494),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_541),
.B(n_472),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_609),
.A2(n_335),
.B1(n_345),
.B2(n_264),
.Y(n_728)
);

NOR3xp33_ASAP7_75t_L g729 ( 
.A(n_557),
.B(n_497),
.C(n_489),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_527),
.B(n_179),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_538),
.B(n_180),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_527),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_613),
.B(n_180),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_640),
.B(n_183),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_646),
.B(n_183),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_548),
.B(n_474),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_618),
.B(n_482),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_548),
.B(n_482),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_550),
.B(n_489),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_561),
.B(n_185),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_620),
.B(n_636),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_561),
.B(n_185),
.Y(n_742)
);

NOR2x1p5_ASAP7_75t_L g743 ( 
.A(n_551),
.B(n_190),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_570),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_645),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_574),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_555),
.B(n_236),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_636),
.B(n_188),
.Y(n_748)
);

INVx8_ASAP7_75t_L g749 ( 
.A(n_661),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_577),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_583),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_588),
.B(n_239),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_622),
.B(n_289),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_577),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_622),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_554),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_641),
.B(n_188),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_578),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_659),
.B(n_191),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_659),
.B(n_191),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_660),
.B(n_195),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_660),
.B(n_195),
.Y(n_762)
);

AND2x6_ASAP7_75t_SL g763 ( 
.A(n_628),
.B(n_203),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_593),
.B(n_198),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_563),
.B(n_198),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_588),
.B(n_242),
.Y(n_766)
);

NOR2xp67_ASAP7_75t_L g767 ( 
.A(n_554),
.B(n_644),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_645),
.Y(n_768)
);

NAND3xp33_ASAP7_75t_L g769 ( 
.A(n_606),
.B(n_291),
.C(n_323),
.Y(n_769)
);

OR2x6_ASAP7_75t_L g770 ( 
.A(n_621),
.B(n_175),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_661),
.A2(n_581),
.B1(n_626),
.B2(n_649),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_578),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_623),
.B(n_246),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_630),
.B(n_249),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_525),
.B(n_189),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_518),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_574),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_595),
.B(n_590),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_595),
.B(n_251),
.Y(n_779)
);

NOR2x1p5_ASAP7_75t_L g780 ( 
.A(n_551),
.B(n_302),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_595),
.B(n_590),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_649),
.B(n_200),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_592),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_525),
.A2(n_347),
.B1(n_315),
.B2(n_321),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_614),
.B(n_202),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_601),
.B(n_602),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_601),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_614),
.B(n_202),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_624),
.B(n_626),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_581),
.B(n_333),
.Y(n_790)
);

BUFx5_ASAP7_75t_L g791 ( 
.A(n_543),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_626),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_528),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_602),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_582),
.Y(n_795)
);

NOR2x1p5_ASAP7_75t_L g796 ( 
.A(n_566),
.B(n_315),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_549),
.B(n_204),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_575),
.B(n_306),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_528),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_580),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_569),
.B(n_253),
.Y(n_801)
);

AND2x2_ASAP7_75t_SL g802 ( 
.A(n_539),
.B(n_175),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_SL g803 ( 
.A(n_591),
.B(n_175),
.Y(n_803)
);

OR2x6_ASAP7_75t_L g804 ( 
.A(n_621),
.B(n_182),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_584),
.B(n_306),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_621),
.B(n_307),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_569),
.B(n_262),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_591),
.B(n_307),
.Y(n_808)
);

O2A1O1Ixp5_ASAP7_75t_L g809 ( 
.A1(n_582),
.A2(n_279),
.B(n_297),
.C(n_268),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_591),
.B(n_310),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_621),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_525),
.A2(n_293),
.B1(n_292),
.B2(n_294),
.Y(n_812)
);

AND2x6_ASAP7_75t_L g813 ( 
.A(n_655),
.B(n_182),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_586),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_530),
.Y(n_815)
);

NAND3xp33_ASAP7_75t_L g816 ( 
.A(n_733),
.B(n_651),
.C(n_611),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_783),
.Y(n_817)
);

NOR3xp33_ASAP7_75t_L g818 ( 
.A(n_672),
.B(n_329),
.C(n_318),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_667),
.B(n_652),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_787),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_670),
.B(n_598),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_692),
.A2(n_547),
.B(n_546),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_794),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_684),
.Y(n_824)
);

O2A1O1Ixp33_ASAP7_75t_SL g825 ( 
.A1(n_686),
.A2(n_666),
.B(n_652),
.C(n_656),
.Y(n_825)
);

OAI321xp33_ASAP7_75t_L g826 ( 
.A1(n_782),
.A2(n_687),
.A3(n_798),
.B1(n_765),
.B2(n_805),
.C(n_784),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_681),
.B(n_662),
.Y(n_827)
);

AO32x1_ASAP7_75t_L g828 ( 
.A1(n_685),
.A2(n_611),
.A3(n_604),
.B1(n_632),
.B2(n_605),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_681),
.B(n_665),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_741),
.B(n_656),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_741),
.B(n_658),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_668),
.B(n_658),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_681),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_737),
.B(n_674),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_679),
.A2(n_525),
.B(n_552),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_731),
.B(n_604),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_737),
.B(n_605),
.Y(n_837)
);

NOR2x1_ASAP7_75t_L g838 ( 
.A(n_716),
.B(n_665),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_681),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_709),
.B(n_632),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_687),
.A2(n_525),
.B1(n_543),
.B2(n_663),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_795),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_815),
.A2(n_781),
.B(n_778),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_777),
.B(n_639),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_693),
.A2(n_663),
.B(n_666),
.C(n_664),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_753),
.B(n_664),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_814),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_732),
.B(n_665),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_684),
.B(n_321),
.Y(n_849)
);

O2A1O1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_695),
.A2(n_530),
.B(n_537),
.C(n_533),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_746),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_696),
.B(n_310),
.Y(n_852)
);

OAI221xp5_ASAP7_75t_L g853 ( 
.A1(n_689),
.A2(n_344),
.B1(n_336),
.B2(n_325),
.C(n_327),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_710),
.B(n_525),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_689),
.A2(n_655),
.B1(n_625),
.B2(n_637),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_798),
.A2(n_537),
.B(n_533),
.C(n_552),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_759),
.A2(n_625),
.B(n_637),
.C(n_638),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_712),
.B(n_517),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_755),
.B(n_311),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_776),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_717),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_719),
.B(n_517),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_800),
.B(n_671),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_721),
.B(n_725),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_759),
.B(n_311),
.Y(n_865)
);

OA21x2_ASAP7_75t_L g866 ( 
.A1(n_680),
.A2(n_288),
.B(n_337),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_677),
.A2(n_532),
.B(n_545),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_746),
.Y(n_868)
);

AO21x1_ASAP7_75t_L g869 ( 
.A1(n_698),
.A2(n_642),
.B(n_543),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_756),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_789),
.B(n_764),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_761),
.B(n_318),
.C(n_346),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_722),
.B(n_639),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_751),
.B(n_625),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_801),
.A2(n_532),
.B(n_545),
.Y(n_875)
);

NOR2x1_ASAP7_75t_L g876 ( 
.A(n_682),
.B(n_767),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_789),
.A2(n_543),
.B1(n_637),
.B2(n_638),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_786),
.B(n_638),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_761),
.A2(n_617),
.B(n_571),
.C(n_587),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_762),
.B(n_325),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_764),
.B(n_517),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_762),
.B(n_327),
.Y(n_882)
);

AOI33xp33_ASAP7_75t_L g883 ( 
.A1(n_702),
.A2(n_347),
.A3(n_330),
.B1(n_328),
.B2(n_308),
.B3(n_182),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_703),
.B(n_543),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_711),
.A2(n_543),
.B1(n_654),
.B2(n_657),
.Y(n_885)
);

NOR2x1_ASAP7_75t_L g886 ( 
.A(n_718),
.B(n_642),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_703),
.B(n_654),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_675),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_807),
.A2(n_562),
.B(n_556),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_704),
.B(n_654),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_705),
.B(n_329),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_706),
.Y(n_892)
);

OR2x2_ASAP7_75t_L g893 ( 
.A(n_768),
.B(n_328),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_746),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_704),
.B(n_654),
.Y(n_895)
);

OAI21xp33_ASAP7_75t_L g896 ( 
.A1(n_765),
.A2(n_330),
.B(n_346),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_707),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_669),
.B(n_332),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_745),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_691),
.A2(n_579),
.B(n_571),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_715),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_746),
.B(n_334),
.Y(n_902)
);

AND2x6_ASAP7_75t_L g903 ( 
.A(n_771),
.B(n_657),
.Y(n_903)
);

BUFx12f_ASAP7_75t_L g904 ( 
.A(n_763),
.Y(n_904)
);

AO21x1_ASAP7_75t_L g905 ( 
.A1(n_782),
.A2(n_642),
.B(n_657),
.Y(n_905)
);

OAI21xp33_ASAP7_75t_L g906 ( 
.A1(n_748),
.A2(n_341),
.B(n_571),
.Y(n_906)
);

OAI21xp33_ASAP7_75t_L g907 ( 
.A1(n_748),
.A2(n_735),
.B(n_734),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_773),
.A2(n_603),
.B(n_526),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_676),
.B(n_587),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_774),
.A2(n_603),
.B(n_526),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_792),
.A2(n_603),
.B(n_526),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_720),
.B(n_535),
.Y(n_912)
);

INVxp67_ASAP7_75t_SL g913 ( 
.A(n_714),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_691),
.A2(n_711),
.B(n_688),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_676),
.B(n_220),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_683),
.B(n_617),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_683),
.B(n_617),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_803),
.B(n_657),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_785),
.A2(n_579),
.B(n_616),
.C(n_599),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_673),
.A2(n_519),
.B1(n_627),
.B2(n_629),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_724),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_727),
.A2(n_585),
.B(n_653),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_678),
.A2(n_627),
.B1(n_629),
.B2(n_653),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_736),
.A2(n_738),
.B(n_739),
.Y(n_924)
);

NAND2xp33_ASAP7_75t_SL g925 ( 
.A(n_811),
.B(n_627),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_811),
.Y(n_926)
);

AO21x1_ASAP7_75t_L g927 ( 
.A1(n_785),
.A2(n_220),
.B(n_273),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_809),
.A2(n_653),
.B(n_585),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_708),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_793),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_779),
.A2(n_629),
.B(n_627),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_802),
.B(n_309),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_718),
.A2(n_627),
.B1(n_309),
.B2(n_308),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_747),
.A2(n_639),
.B(n_124),
.Y(n_934)
);

NAND2x1p5_ASAP7_75t_L g935 ( 
.A(n_714),
.B(n_114),
.Y(n_935)
);

AND2x2_ASAP7_75t_SL g936 ( 
.A(n_802),
.B(n_309),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_713),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_799),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_770),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_723),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_788),
.B(n_308),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_752),
.B(n_220),
.Y(n_942)
);

CKINVDCx10_ASAP7_75t_R g943 ( 
.A(n_699),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_730),
.A2(n_273),
.B(n_12),
.C(n_14),
.Y(n_944)
);

NOR3xp33_ASAP7_75t_L g945 ( 
.A(n_690),
.B(n_273),
.C(n_16),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_766),
.A2(n_168),
.B(n_156),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_744),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_788),
.B(n_136),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_750),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_754),
.Y(n_950)
);

OAI321xp33_ASAP7_75t_L g951 ( 
.A1(n_784),
.A2(n_10),
.A3(n_18),
.B1(n_19),
.B2(n_29),
.C(n_30),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_694),
.Y(n_952)
);

AOI211xp5_ASAP7_75t_L g953 ( 
.A1(n_769),
.A2(n_29),
.B(n_34),
.C(n_35),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_701),
.B(n_125),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_L g955 ( 
.A(n_758),
.B(n_108),
.Y(n_955)
);

AND2x2_ASAP7_75t_SL g956 ( 
.A(n_729),
.B(n_34),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_772),
.B(n_96),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_757),
.A2(n_35),
.B(n_37),
.C(n_39),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_790),
.B(n_84),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_697),
.B(n_43),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_775),
.Y(n_961)
);

AO22x1_ASAP7_75t_L g962 ( 
.A1(n_806),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_797),
.A2(n_810),
.B(n_808),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_728),
.B(n_44),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_760),
.Y(n_965)
);

CKINVDCx8_ASAP7_75t_R g966 ( 
.A(n_700),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_791),
.Y(n_967)
);

AO21x1_ASAP7_75t_L g968 ( 
.A1(n_740),
.A2(n_742),
.B(n_812),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_726),
.A2(n_45),
.B(n_47),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_770),
.A2(n_48),
.B(n_49),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_770),
.A2(n_49),
.B(n_50),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_700),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_804),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_791),
.B(n_51),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_791),
.B(n_55),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_791),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_813),
.B(n_804),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_L g978 ( 
.A(n_700),
.B(n_55),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_749),
.B(n_58),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_804),
.A2(n_58),
.B1(n_749),
.B2(n_796),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_743),
.A2(n_780),
.B(n_813),
.C(n_749),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_SL g982 ( 
.A1(n_822),
.A2(n_914),
.B(n_834),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_861),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_839),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_910),
.A2(n_813),
.B(n_835),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_824),
.B(n_891),
.Y(n_986)
);

AO21x2_ASAP7_75t_L g987 ( 
.A1(n_905),
.A2(n_825),
.B(n_869),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_L g988 ( 
.A1(n_849),
.A2(n_865),
.B(n_880),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_836),
.B(n_907),
.Y(n_989)
);

AOI221x1_ASAP7_75t_L g990 ( 
.A1(n_818),
.A2(n_816),
.B1(n_879),
.B2(n_945),
.C(n_919),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_826),
.A2(n_871),
.B(n_936),
.C(n_960),
.Y(n_991)
);

AO21x1_ASAP7_75t_L g992 ( 
.A1(n_948),
.A2(n_932),
.B(n_974),
.Y(n_992)
);

AO31x2_ASAP7_75t_L g993 ( 
.A1(n_845),
.A2(n_857),
.A3(n_927),
.B(n_856),
.Y(n_993)
);

INVx5_ASAP7_75t_L g994 ( 
.A(n_839),
.Y(n_994)
);

AO31x2_ASAP7_75t_L g995 ( 
.A1(n_819),
.A2(n_832),
.A3(n_975),
.B(n_974),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_924),
.A2(n_890),
.B(n_887),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_882),
.B(n_915),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_949),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_870),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_887),
.A2(n_895),
.B(n_890),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_892),
.B(n_897),
.Y(n_1001)
);

INVxp67_ASAP7_75t_SL g1002 ( 
.A(n_839),
.Y(n_1002)
);

OAI22x1_ASAP7_75t_L g1003 ( 
.A1(n_921),
.A2(n_973),
.B1(n_863),
.B2(n_965),
.Y(n_1003)
);

NOR2xp67_ASAP7_75t_L g1004 ( 
.A(n_872),
.B(n_952),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_820),
.Y(n_1005)
);

AO21x2_ASAP7_75t_L g1006 ( 
.A1(n_881),
.A2(n_831),
.B(n_830),
.Y(n_1006)
);

AOI31xp33_ASAP7_75t_L g1007 ( 
.A1(n_953),
.A2(n_980),
.A3(n_964),
.B(n_977),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_851),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_968),
.A2(n_846),
.B1(n_959),
.B2(n_876),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_851),
.B(n_868),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_899),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_972),
.B(n_844),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_884),
.A2(n_900),
.B(n_850),
.Y(n_1013)
);

OAI222xp33_ASAP7_75t_L g1014 ( 
.A1(n_853),
.A2(n_979),
.B1(n_971),
.B2(n_970),
.C1(n_969),
.C2(n_941),
.Y(n_1014)
);

AO31x2_ASAP7_75t_L g1015 ( 
.A1(n_975),
.A2(n_855),
.A3(n_830),
.B(n_831),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_888),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_931),
.A2(n_875),
.B(n_889),
.Y(n_1017)
);

AO21x1_ASAP7_75t_L g1018 ( 
.A1(n_959),
.A2(n_954),
.B(n_852),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_840),
.B(n_821),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_851),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_926),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_963),
.A2(n_896),
.B(n_901),
.C(n_864),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_837),
.A2(n_864),
.B1(n_841),
.B2(n_884),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_949),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_860),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_878),
.A2(n_961),
.B(n_885),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_823),
.B(n_909),
.Y(n_1027)
);

AOI21x1_ASAP7_75t_SL g1028 ( 
.A1(n_977),
.A2(n_854),
.B(n_954),
.Y(n_1028)
);

NOR3xp33_ASAP7_75t_L g1029 ( 
.A(n_859),
.B(n_978),
.C(n_898),
.Y(n_1029)
);

NAND2x1p5_ASAP7_75t_L g1030 ( 
.A(n_868),
.B(n_833),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_912),
.B(n_916),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_878),
.A2(n_917),
.B(n_894),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_956),
.B(n_893),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_874),
.A2(n_877),
.B(n_957),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_981),
.B(n_939),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_883),
.B(n_942),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_842),
.B(n_847),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_943),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_930),
.B(n_938),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_967),
.A2(n_886),
.B(n_911),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_944),
.A2(n_958),
.B(n_906),
.C(n_951),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_928),
.A2(n_920),
.B(n_829),
.Y(n_1042)
);

INVx6_ASAP7_75t_L g1043 ( 
.A(n_844),
.Y(n_1043)
);

OAI21xp33_ASAP7_75t_SL g1044 ( 
.A1(n_848),
.A2(n_918),
.B(n_858),
.Y(n_1044)
);

AO31x2_ASAP7_75t_L g1045 ( 
.A1(n_957),
.A2(n_934),
.A3(n_828),
.B(n_862),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_827),
.A2(n_829),
.B(n_923),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_L g1047 ( 
.A(n_962),
.B(n_933),
.C(n_902),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_947),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_966),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_929),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_937),
.A2(n_940),
.B(n_950),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_833),
.B(n_903),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_903),
.B(n_913),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_903),
.A2(n_925),
.B1(n_873),
.B2(n_838),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_873),
.Y(n_1055)
);

NAND3xp33_ASAP7_75t_L g1056 ( 
.A(n_946),
.B(n_866),
.C(n_922),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_866),
.A2(n_828),
.B(n_955),
.Y(n_1057)
);

BUFx8_ASAP7_75t_L g1058 ( 
.A(n_904),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_903),
.B(n_935),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_903),
.A2(n_955),
.B(n_935),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_SL g1061 ( 
.A1(n_828),
.A2(n_891),
.B(n_672),
.Y(n_1061)
);

O2A1O1Ixp5_ASAP7_75t_L g1062 ( 
.A1(n_891),
.A2(n_733),
.B(n_865),
.C(n_692),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_826),
.B(n_553),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_888),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_899),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_826),
.B(n_553),
.Y(n_1066)
);

AND2x6_ASAP7_75t_L g1067 ( 
.A(n_976),
.B(n_967),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_926),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_834),
.B(n_573),
.Y(n_1069)
);

NAND3xp33_ASAP7_75t_L g1070 ( 
.A(n_891),
.B(n_865),
.C(n_672),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_834),
.B(n_573),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_834),
.B(n_573),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_817),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_826),
.A2(n_907),
.B(n_865),
.C(n_672),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_870),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_861),
.Y(n_1076)
);

AOI21xp33_ASAP7_75t_L g1077 ( 
.A1(n_826),
.A2(n_907),
.B(n_865),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_861),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_834),
.A2(n_687),
.B1(n_936),
.B2(n_689),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_817),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_834),
.B(n_573),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_834),
.B(n_573),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_822),
.A2(n_692),
.B(n_843),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_914),
.A2(n_826),
.B(n_679),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_914),
.A2(n_826),
.B(n_679),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_834),
.A2(n_687),
.B1(n_936),
.B2(n_689),
.Y(n_1086)
);

AOI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_826),
.A2(n_907),
.B(n_865),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_834),
.B(n_573),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_834),
.B(n_573),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_899),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_849),
.B(n_553),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_834),
.B(n_573),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_822),
.A2(n_692),
.B(n_843),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_834),
.A2(n_687),
.B1(n_936),
.B2(n_689),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_822),
.A2(n_692),
.B(n_843),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_834),
.B(n_573),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_914),
.A2(n_826),
.B(n_679),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_914),
.A2(n_826),
.B(n_679),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_834),
.B(n_573),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_834),
.B(n_573),
.Y(n_1100)
);

AO31x2_ASAP7_75t_L g1101 ( 
.A1(n_905),
.A2(n_869),
.A3(n_879),
.B(n_919),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_817),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_839),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_867),
.A2(n_910),
.B(n_908),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_914),
.A2(n_826),
.B(n_679),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_826),
.A2(n_907),
.B(n_865),
.C(n_672),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_867),
.A2(n_910),
.B(n_908),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_867),
.A2(n_910),
.B(n_908),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_888),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_849),
.B(n_553),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_834),
.B(n_573),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_834),
.B(n_573),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_826),
.B(n_553),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_983),
.Y(n_1114)
);

OR2x6_ASAP7_75t_L g1115 ( 
.A(n_1035),
.B(n_1109),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1088),
.A2(n_1112),
.B1(n_1082),
.B2(n_1111),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1069),
.B(n_1071),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_SL g1118 ( 
.A1(n_1079),
.A2(n_1094),
.B(n_1086),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_1043),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_SL g1120 ( 
.A1(n_1074),
.A2(n_1106),
.B(n_991),
.C(n_1087),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1069),
.B(n_1071),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1011),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1005),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1070),
.A2(n_986),
.B1(n_1029),
.B2(n_988),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_1043),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1076),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_999),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1072),
.A2(n_1082),
.B1(n_1111),
.B2(n_1081),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_SL g1129 ( 
.A(n_1079),
.B(n_1086),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1091),
.B(n_1110),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1019),
.B(n_1033),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1078),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_997),
.B(n_1036),
.Y(n_1133)
);

AND2x2_ASAP7_75t_SL g1134 ( 
.A(n_1059),
.B(n_989),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1043),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1037),
.Y(n_1136)
);

OR2x6_ASAP7_75t_L g1137 ( 
.A(n_1035),
.B(n_1059),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1012),
.B(n_1055),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1073),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1072),
.B(n_1081),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1089),
.B(n_1092),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1037),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_994),
.Y(n_1143)
);

OR2x2_ASAP7_75t_L g1144 ( 
.A(n_1089),
.B(n_1092),
.Y(n_1144)
);

BUFx2_ASAP7_75t_SL g1145 ( 
.A(n_1065),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1077),
.A2(n_1087),
.B(n_1063),
.C(n_1066),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1080),
.Y(n_1147)
);

OR2x6_ASAP7_75t_L g1148 ( 
.A(n_1035),
.B(n_1016),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1039),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_1075),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1102),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_SL g1152 ( 
.A1(n_1094),
.A2(n_1096),
.B1(n_1099),
.B2(n_1100),
.Y(n_1152)
);

NOR2x1p5_ASAP7_75t_L g1153 ( 
.A(n_1047),
.B(n_1038),
.Y(n_1153)
);

NOR2xp67_ASAP7_75t_L g1154 ( 
.A(n_1090),
.B(n_1003),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1021),
.B(n_1068),
.Y(n_1155)
);

INVx2_ASAP7_75t_SL g1156 ( 
.A(n_1064),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_984),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1050),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1004),
.B(n_1001),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1049),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1012),
.B(n_998),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1096),
.A2(n_1099),
.B1(n_1100),
.B2(n_1001),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_984),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1025),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1077),
.A2(n_1027),
.B1(n_1105),
.B2(n_1098),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_1058),
.Y(n_1166)
);

INVx5_ASAP7_75t_L g1167 ( 
.A(n_984),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1007),
.B(n_1113),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_994),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1048),
.B(n_1024),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1014),
.B(n_1009),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1058),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1027),
.A2(n_1085),
.B1(n_1105),
.B2(n_1098),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_1018),
.A2(n_1057),
.A3(n_992),
.B(n_1083),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1060),
.B(n_1010),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1051),
.B(n_1022),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1008),
.B(n_1103),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1020),
.Y(n_1178)
);

AND2x6_ASAP7_75t_L g1179 ( 
.A(n_1054),
.B(n_1052),
.Y(n_1179)
);

NAND2xp33_ASAP7_75t_L g1180 ( 
.A(n_1041),
.B(n_994),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1051),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_994),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1020),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1103),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1030),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1062),
.A2(n_1085),
.B(n_1084),
.C(n_1097),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1030),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1000),
.B(n_1031),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_1084),
.A2(n_1097),
.B(n_985),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_1002),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1044),
.B(n_1053),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1093),
.A2(n_1095),
.B(n_982),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_995),
.B(n_1052),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_SL g1194 ( 
.A1(n_1060),
.A2(n_1053),
.B(n_1034),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1023),
.B(n_1006),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1023),
.B(n_1006),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_990),
.B(n_1046),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_995),
.B(n_996),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_993),
.Y(n_1199)
);

AND2x2_ASAP7_75t_SL g1200 ( 
.A(n_1061),
.B(n_1028),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1034),
.A2(n_1026),
.B(n_1032),
.Y(n_1201)
);

CKINVDCx14_ASAP7_75t_R g1202 ( 
.A(n_1067),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1013),
.A2(n_1040),
.B(n_1042),
.C(n_1056),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1015),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1015),
.B(n_1013),
.Y(n_1205)
);

NAND2xp33_ASAP7_75t_L g1206 ( 
.A(n_1015),
.B(n_1101),
.Y(n_1206)
);

OA21x2_ASAP7_75t_L g1207 ( 
.A1(n_1108),
.A2(n_1107),
.B(n_1104),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1101),
.B(n_987),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1045),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1045),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1017),
.B(n_1091),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1068),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1069),
.B(n_1071),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1012),
.B(n_1055),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1091),
.B(n_1110),
.Y(n_1215)
);

CKINVDCx6p67_ASAP7_75t_R g1216 ( 
.A(n_1011),
.Y(n_1216)
);

INVx5_ASAP7_75t_L g1217 ( 
.A(n_984),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1074),
.A2(n_1106),
.B(n_1077),
.C(n_1087),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_999),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1069),
.B(n_1071),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1012),
.B(n_1055),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_983),
.Y(n_1222)
);

AOI221xp5_ASAP7_75t_L g1223 ( 
.A1(n_1077),
.A2(n_1087),
.B1(n_826),
.B2(n_986),
.C(n_672),
.Y(n_1223)
);

INVx3_ASAP7_75t_SL g1224 ( 
.A(n_999),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1043),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_984),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_983),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1069),
.B(n_1071),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1012),
.B(n_1055),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1062),
.A2(n_826),
.B(n_1070),
.C(n_1077),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_983),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_983),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_986),
.B(n_553),
.Y(n_1233)
);

OR2x6_ASAP7_75t_L g1234 ( 
.A(n_1035),
.B(n_1109),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_986),
.B(n_553),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1070),
.A2(n_891),
.B1(n_865),
.B2(n_369),
.Y(n_1236)
);

BUFx12f_ASAP7_75t_L g1237 ( 
.A(n_1038),
.Y(n_1237)
);

O2A1O1Ixp5_ASAP7_75t_SL g1238 ( 
.A1(n_1077),
.A2(n_1087),
.B(n_932),
.C(n_1066),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_SL g1239 ( 
.A1(n_1077),
.A2(n_891),
.B(n_826),
.C(n_733),
.Y(n_1239)
);

CKINVDCx8_ASAP7_75t_R g1240 ( 
.A(n_999),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1091),
.B(n_1110),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1021),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1069),
.B(n_1071),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_1021),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_986),
.B(n_553),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1043),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1043),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1091),
.B(n_1110),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1068),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1242),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1245),
.B(n_1236),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1123),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1223),
.A2(n_1168),
.B1(n_1129),
.B2(n_1171),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1122),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1223),
.A2(n_1129),
.B1(n_1152),
.B2(n_1124),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1126),
.Y(n_1256)
);

AO21x1_ASAP7_75t_L g1257 ( 
.A1(n_1218),
.A2(n_1146),
.B(n_1180),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1182),
.Y(n_1258)
);

NAND2x1p5_ASAP7_75t_L g1259 ( 
.A(n_1143),
.B(n_1169),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1116),
.B(n_1128),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1155),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_SL g1262 ( 
.A1(n_1146),
.A2(n_1194),
.B(n_1218),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1137),
.B(n_1185),
.Y(n_1263)
);

OAI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1144),
.A2(n_1213),
.B1(n_1141),
.B2(n_1117),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1132),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1152),
.A2(n_1116),
.B1(n_1128),
.B2(n_1162),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1182),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1117),
.A2(n_1140),
.B1(n_1228),
.B2(n_1243),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1162),
.A2(n_1133),
.B1(n_1165),
.B2(n_1131),
.Y(n_1269)
);

INVx6_ASAP7_75t_L g1270 ( 
.A(n_1167),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1165),
.A2(n_1159),
.B1(n_1176),
.B2(n_1141),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1216),
.Y(n_1272)
);

AO21x1_ASAP7_75t_L g1273 ( 
.A1(n_1173),
.A2(n_1191),
.B(n_1186),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1227),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1182),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1121),
.A2(n_1220),
.B1(n_1228),
.B2(n_1140),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1121),
.A2(n_1220),
.B1(n_1213),
.B2(n_1243),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1127),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1150),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1173),
.A2(n_1154),
.B1(n_1142),
.B2(n_1136),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_SL g1281 ( 
.A1(n_1166),
.A2(n_1248),
.B1(n_1215),
.B2(n_1241),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1233),
.B(n_1235),
.Y(n_1282)
);

AO21x1_ASAP7_75t_SL g1283 ( 
.A1(n_1208),
.A2(n_1199),
.B(n_1204),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1244),
.Y(n_1284)
);

OAI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1115),
.A2(n_1234),
.B1(n_1148),
.B2(n_1156),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1153),
.A2(n_1181),
.B1(n_1179),
.B2(n_1188),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1222),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_1219),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1231),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1240),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1237),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1232),
.Y(n_1292)
);

BUFx2_ASAP7_75t_SL g1293 ( 
.A(n_1167),
.Y(n_1293)
);

BUFx4_ASAP7_75t_R g1294 ( 
.A(n_1160),
.Y(n_1294)
);

INVx8_ASAP7_75t_L g1295 ( 
.A(n_1167),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1179),
.A2(n_1188),
.B1(n_1234),
.B2(n_1115),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1167),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1149),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1244),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_1224),
.Y(n_1300)
);

INVx6_ASAP7_75t_SL g1301 ( 
.A(n_1148),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1115),
.A2(n_1234),
.B1(n_1148),
.B2(n_1137),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1130),
.B(n_1212),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1178),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1212),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1158),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1193),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1164),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1134),
.A2(n_1179),
.B1(n_1211),
.B2(n_1137),
.Y(n_1309)
);

NAND2x1p5_ASAP7_75t_L g1310 ( 
.A(n_1143),
.B(n_1169),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1139),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1147),
.Y(n_1312)
);

BUFx2_ASAP7_75t_R g1313 ( 
.A(n_1172),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1177),
.Y(n_1314)
);

INVxp33_ASAP7_75t_L g1315 ( 
.A(n_1249),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1151),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1185),
.B(n_1187),
.Y(n_1317)
);

AO21x2_ASAP7_75t_L g1318 ( 
.A1(n_1192),
.A2(n_1203),
.B(n_1201),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1170),
.Y(n_1319)
);

INVx6_ASAP7_75t_L g1320 ( 
.A(n_1217),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1184),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1230),
.B(n_1120),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1249),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1190),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1163),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1217),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1161),
.Y(n_1327)
);

BUFx2_ASAP7_75t_R g1328 ( 
.A(n_1145),
.Y(n_1328)
);

INVx6_ASAP7_75t_L g1329 ( 
.A(n_1217),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1183),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1187),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1161),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1217),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1179),
.A2(n_1205),
.B1(n_1189),
.B2(n_1200),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1177),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1195),
.A2(n_1196),
.B(n_1198),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1202),
.A2(n_1179),
.B1(n_1239),
.B2(n_1197),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1197),
.A2(n_1175),
.B1(n_1118),
.B2(n_1221),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1175),
.A2(n_1119),
.B1(n_1125),
.B2(n_1135),
.Y(n_1339)
);

AOI222xp33_ASAP7_75t_L g1340 ( 
.A1(n_1138),
.A2(n_1229),
.B1(n_1221),
.B2(n_1214),
.C1(n_1206),
.C2(n_1196),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1138),
.B(n_1229),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1209),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1214),
.A2(n_1175),
.B1(n_1125),
.B2(n_1135),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1119),
.B(n_1247),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1157),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1225),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1207),
.A2(n_1186),
.B(n_1208),
.Y(n_1347)
);

INVx5_ASAP7_75t_L g1348 ( 
.A(n_1157),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1246),
.A2(n_1226),
.B1(n_1210),
.B2(n_1238),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1226),
.B(n_1174),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1174),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1174),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1114),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1116),
.B(n_1128),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1137),
.B(n_1185),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1124),
.B(n_1070),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1155),
.Y(n_1357)
);

OAI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1236),
.A2(n_826),
.B1(n_921),
.B2(n_672),
.Y(n_1358)
);

BUFx12f_ASAP7_75t_L g1359 ( 
.A(n_1219),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1114),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1223),
.A2(n_936),
.B1(n_1087),
.B2(n_1077),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1242),
.Y(n_1362)
);

CKINVDCx6p67_ASAP7_75t_R g1363 ( 
.A(n_1224),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1236),
.A2(n_891),
.B1(n_921),
.B2(n_1088),
.Y(n_1364)
);

OR2x6_ASAP7_75t_L g1365 ( 
.A(n_1148),
.B(n_1137),
.Y(n_1365)
);

OAI21xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1255),
.A2(n_1361),
.B(n_1253),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1342),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1324),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1307),
.B(n_1260),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1284),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1350),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1307),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1354),
.B(n_1334),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1299),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1365),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_1365),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1334),
.B(n_1266),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1365),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1350),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1336),
.B(n_1266),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1347),
.Y(n_1381)
);

AOI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1356),
.A2(n_1349),
.B(n_1273),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1351),
.A2(n_1352),
.B(n_1262),
.Y(n_1383)
);

NAND2x1p5_ASAP7_75t_L g1384 ( 
.A(n_1350),
.B(n_1263),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1297),
.A2(n_1326),
.B(n_1333),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1336),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1295),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1271),
.B(n_1255),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1336),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1352),
.A2(n_1257),
.B(n_1271),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1298),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1253),
.B(n_1269),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1251),
.A2(n_1358),
.B1(n_1364),
.B2(n_1361),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1318),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1269),
.A2(n_1322),
.B(n_1280),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1251),
.A2(n_1276),
.B1(n_1277),
.B2(n_1280),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1292),
.B(n_1276),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1305),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1303),
.B(n_1296),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1263),
.B(n_1355),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1268),
.B(n_1264),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1357),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1286),
.A2(n_1296),
.B(n_1309),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1323),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1277),
.B(n_1286),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1288),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1263),
.B(n_1355),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1261),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1287),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1341),
.B(n_1261),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1340),
.B(n_1289),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1321),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1355),
.Y(n_1413)
);

AOI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1308),
.A2(n_1331),
.B(n_1252),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1282),
.B(n_1281),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1256),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1282),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1265),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1315),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1283),
.B(n_1337),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1338),
.B(n_1319),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1422)
);

INVx5_ASAP7_75t_SL g1423 ( 
.A(n_1363),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1339),
.A2(n_1302),
.B(n_1285),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1301),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1274),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1301),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1353),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1360),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1301),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1315),
.B(n_1250),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1343),
.A2(n_1306),
.B(n_1316),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1311),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1297),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1312),
.B(n_1317),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1317),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1362),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1332),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1330),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1327),
.B(n_1346),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1317),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1293),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1344),
.B(n_1314),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1259),
.Y(n_1444)
);

AND2x4_ASAP7_75t_SL g1445 ( 
.A(n_1400),
.B(n_1363),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1367),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1419),
.B(n_1402),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1373),
.B(n_1335),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1393),
.A2(n_1330),
.B1(n_1290),
.B2(n_1325),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1379),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_1375),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1371),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1374),
.B(n_1278),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1368),
.B(n_1304),
.Y(n_1454)
);

AOI221xp5_ASAP7_75t_L g1455 ( 
.A1(n_1396),
.A2(n_1254),
.B1(n_1272),
.B2(n_1304),
.C(n_1325),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1369),
.B(n_1258),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1417),
.B(n_1288),
.Y(n_1457)
);

NOR2x1_ASAP7_75t_L g1458 ( 
.A(n_1385),
.B(n_1300),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1370),
.B(n_1290),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1431),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1370),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1369),
.B(n_1267),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1375),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1380),
.B(n_1275),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_SL g1465 ( 
.A1(n_1366),
.A2(n_1300),
.B1(n_1329),
.B2(n_1270),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1409),
.Y(n_1466)
);

OAI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1366),
.A2(n_1272),
.B1(n_1310),
.B2(n_1259),
.C(n_1275),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1371),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1412),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1409),
.Y(n_1470)
);

AND2x4_ASAP7_75t_SL g1471 ( 
.A(n_1400),
.B(n_1407),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1409),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1431),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1432),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1371),
.B(n_1376),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1397),
.B(n_1348),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1380),
.B(n_1310),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1432),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1396),
.B(n_1359),
.Y(n_1479)
);

INVxp67_ASAP7_75t_SL g1480 ( 
.A(n_1404),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1376),
.B(n_1378),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1399),
.B(n_1294),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1392),
.A2(n_1359),
.B1(n_1291),
.B2(n_1345),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1432),
.Y(n_1484)
);

OR2x6_ASAP7_75t_L g1485 ( 
.A(n_1376),
.B(n_1270),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1372),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1398),
.B(n_1345),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1378),
.B(n_1294),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1384),
.B(n_1328),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1384),
.B(n_1320),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1415),
.A2(n_1313),
.B1(n_1320),
.B2(n_1329),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1381),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1377),
.B(n_1320),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1392),
.A2(n_1388),
.B1(n_1377),
.B2(n_1424),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1414),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1399),
.B(n_1291),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1414),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1386),
.B(n_1389),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1398),
.B(n_1411),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1411),
.B(n_1401),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1473),
.B(n_1405),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1479),
.A2(n_1388),
.B1(n_1424),
.B2(n_1403),
.Y(n_1502)
);

NAND3xp33_ASAP7_75t_L g1503 ( 
.A(n_1455),
.B(n_1494),
.C(n_1500),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1452),
.B(n_1403),
.Y(n_1504)
);

NAND4xp25_ASAP7_75t_L g1505 ( 
.A(n_1499),
.B(n_1405),
.C(n_1437),
.D(n_1410),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1458),
.B(n_1400),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1452),
.B(n_1468),
.Y(n_1507)
);

AOI21xp33_ASAP7_75t_L g1508 ( 
.A1(n_1496),
.A2(n_1424),
.B(n_1420),
.Y(n_1508)
);

NAND4xp25_ASAP7_75t_L g1509 ( 
.A(n_1449),
.B(n_1437),
.C(n_1421),
.D(n_1440),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1465),
.B(n_1438),
.C(n_1421),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1458),
.B(n_1400),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1460),
.B(n_1408),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1447),
.B(n_1408),
.Y(n_1513)
);

OA211x2_ASAP7_75t_L g1514 ( 
.A1(n_1483),
.A2(n_1422),
.B(n_1423),
.C(n_1385),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1469),
.B(n_1432),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1475),
.B(n_1403),
.Y(n_1516)
);

OAI221xp5_ASAP7_75t_L g1517 ( 
.A1(n_1496),
.A2(n_1378),
.B1(n_1430),
.B2(n_1439),
.C(n_1425),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1480),
.B(n_1418),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1482),
.A2(n_1424),
.B1(n_1420),
.B2(n_1413),
.Y(n_1519)
);

OAI221xp5_ASAP7_75t_SL g1520 ( 
.A1(n_1467),
.A2(n_1482),
.B1(n_1459),
.B2(n_1477),
.C(n_1453),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1461),
.B(n_1418),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1488),
.A2(n_1395),
.B(n_1390),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1475),
.B(n_1383),
.Y(n_1523)
);

OAI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1491),
.A2(n_1430),
.B1(n_1439),
.B2(n_1425),
.C(n_1427),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1446),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1448),
.B(n_1428),
.Y(n_1526)
);

OAI221xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1477),
.A2(n_1440),
.B1(n_1439),
.B2(n_1427),
.C(n_1425),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_R g1528 ( 
.A(n_1489),
.B(n_1406),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1475),
.B(n_1383),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1488),
.A2(n_1423),
.B1(n_1395),
.B2(n_1425),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1448),
.B(n_1383),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1456),
.B(n_1428),
.Y(n_1532)
);

OAI21xp33_ASAP7_75t_L g1533 ( 
.A1(n_1457),
.A2(n_1382),
.B(n_1474),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1456),
.B(n_1428),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1488),
.A2(n_1423),
.B1(n_1395),
.B2(n_1427),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1488),
.A2(n_1423),
.B1(n_1395),
.B2(n_1427),
.Y(n_1536)
);

OAI221xp5_ASAP7_75t_SL g1537 ( 
.A1(n_1487),
.A2(n_1454),
.B1(n_1464),
.B2(n_1484),
.C(n_1478),
.Y(n_1537)
);

OAI21xp33_ASAP7_75t_L g1538 ( 
.A1(n_1493),
.A2(n_1382),
.B(n_1435),
.Y(n_1538)
);

AOI21xp33_ASAP7_75t_L g1539 ( 
.A1(n_1464),
.A2(n_1442),
.B(n_1436),
.Y(n_1539)
);

NOR3xp33_ASAP7_75t_L g1540 ( 
.A(n_1495),
.B(n_1444),
.C(n_1442),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1462),
.B(n_1436),
.Y(n_1541)
);

NOR3xp33_ASAP7_75t_L g1542 ( 
.A(n_1495),
.B(n_1444),
.C(n_1434),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1493),
.A2(n_1413),
.B1(n_1407),
.B2(n_1436),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1462),
.B(n_1416),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1489),
.A2(n_1407),
.B(n_1387),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1481),
.B(n_1450),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_SL g1547 ( 
.A(n_1445),
.B(n_1407),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1481),
.A2(n_1413),
.B1(n_1441),
.B2(n_1443),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1445),
.B(n_1423),
.Y(n_1549)
);

NAND4xp25_ASAP7_75t_L g1550 ( 
.A(n_1497),
.B(n_1426),
.C(n_1429),
.D(n_1433),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1486),
.B(n_1391),
.Y(n_1551)
);

INVxp67_ASAP7_75t_SL g1552 ( 
.A(n_1515),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1501),
.B(n_1466),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1525),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1525),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1533),
.B(n_1466),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1503),
.A2(n_1463),
.B1(n_1490),
.B2(n_1451),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1533),
.B(n_1498),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1523),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1528),
.B(n_1445),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1529),
.Y(n_1561)
);

NOR2xp67_ASAP7_75t_L g1562 ( 
.A(n_1550),
.B(n_1498),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1516),
.B(n_1529),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1531),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1551),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1507),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1504),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1526),
.B(n_1450),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1518),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1532),
.Y(n_1570)
);

NOR2xp67_ASAP7_75t_L g1571 ( 
.A(n_1506),
.B(n_1492),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1507),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1521),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1522),
.B(n_1492),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1540),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1534),
.B(n_1470),
.Y(n_1576)
);

BUFx2_ASAP7_75t_R g1577 ( 
.A(n_1511),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1522),
.B(n_1394),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1546),
.B(n_1541),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1544),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1512),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1538),
.B(n_1472),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1538),
.B(n_1394),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1513),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1575),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1562),
.B(n_1510),
.Y(n_1586)
);

AND2x4_ASAP7_75t_L g1587 ( 
.A(n_1571),
.B(n_1542),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1554),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1554),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1571),
.B(n_1547),
.Y(n_1590)
);

NAND2x1_ASAP7_75t_L g1591 ( 
.A(n_1566),
.B(n_1485),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1562),
.B(n_1549),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1584),
.B(n_1502),
.Y(n_1593)
);

A2O1A1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1575),
.A2(n_1510),
.B(n_1520),
.C(n_1508),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1584),
.B(n_1537),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1566),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1555),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1565),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1579),
.B(n_1471),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1565),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1561),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1566),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1569),
.B(n_1505),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1579),
.B(n_1563),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1569),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1573),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1581),
.B(n_1530),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1573),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1557),
.B(n_1519),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1574),
.B(n_1471),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1576),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1563),
.B(n_1543),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1576),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1553),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1581),
.B(n_1539),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1558),
.B(n_1535),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1577),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1580),
.B(n_1476),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1558),
.B(n_1536),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1568),
.B(n_1548),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1568),
.B(n_1527),
.Y(n_1621)
);

BUFx2_ASAP7_75t_SL g1622 ( 
.A(n_1560),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1601),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1597),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1610),
.B(n_1566),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1603),
.B(n_1580),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1596),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1601),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1597),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1585),
.B(n_1552),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1610),
.B(n_1574),
.Y(n_1631)
);

INVxp33_ASAP7_75t_SL g1632 ( 
.A(n_1617),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1588),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1589),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1603),
.B(n_1570),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1610),
.B(n_1563),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1598),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1600),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1604),
.Y(n_1639)
);

CKINVDCx16_ASAP7_75t_R g1640 ( 
.A(n_1622),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1591),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1606),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1585),
.B(n_1570),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1586),
.A2(n_1514),
.B1(n_1524),
.B2(n_1509),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1590),
.B(n_1567),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1605),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1608),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1590),
.B(n_1567),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1614),
.B(n_1556),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1613),
.B(n_1595),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1590),
.B(n_1596),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1596),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1593),
.B(n_1556),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1615),
.B(n_1552),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1618),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1602),
.Y(n_1657)
);

CKINVDCx16_ASAP7_75t_R g1658 ( 
.A(n_1592),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1607),
.B(n_1582),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1620),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1621),
.B(n_1582),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1602),
.Y(n_1662)
);

AOI322xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1586),
.A2(n_1574),
.A3(n_1577),
.B1(n_1583),
.B2(n_1572),
.C1(n_1578),
.C2(n_1564),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1592),
.B(n_1559),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1651),
.B(n_1616),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1636),
.B(n_1592),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1658),
.B(n_1587),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1660),
.B(n_1619),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1632),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1629),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1626),
.B(n_1594),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1629),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1632),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1623),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1640),
.B(n_1587),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1651),
.B(n_1553),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1636),
.B(n_1587),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1623),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1644),
.B(n_1594),
.Y(n_1679)
);

AND3x1_ASAP7_75t_L g1680 ( 
.A(n_1663),
.B(n_1545),
.C(n_1612),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1633),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1661),
.B(n_1609),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1631),
.B(n_1559),
.Y(n_1683)
);

AND2x2_ASAP7_75t_SL g1684 ( 
.A(n_1663),
.B(n_1578),
.Y(n_1684)
);

INVx4_ASAP7_75t_L g1685 ( 
.A(n_1641),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1661),
.B(n_1564),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1628),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1633),
.Y(n_1688)
);

BUFx3_ASAP7_75t_L g1689 ( 
.A(n_1627),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1652),
.B(n_1599),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1634),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1630),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1628),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1634),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1631),
.B(n_1664),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1654),
.A2(n_1609),
.B1(n_1514),
.B2(n_1517),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1680),
.A2(n_1684),
.B1(n_1679),
.B2(n_1671),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1669),
.B(n_1635),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1691),
.Y(n_1699)
);

OAI31xp33_ASAP7_75t_L g1700 ( 
.A1(n_1696),
.A2(n_1671),
.A3(n_1682),
.B(n_1680),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1675),
.B(n_1625),
.Y(n_1701)
);

A2O1A1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1684),
.A2(n_1641),
.B(n_1655),
.C(n_1659),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1675),
.B(n_1631),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_L g1704 ( 
.A(n_1669),
.B(n_1641),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1691),
.Y(n_1705)
);

NAND2xp33_ASAP7_75t_SL g1706 ( 
.A(n_1675),
.B(n_1630),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1667),
.B(n_1664),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1684),
.A2(n_1643),
.B(n_1649),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1694),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1689),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1667),
.B(n_1645),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1689),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1689),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1673),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1673),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1696),
.A2(n_1656),
.B1(n_1650),
.B2(n_1655),
.Y(n_1716)
);

OAI21xp33_ASAP7_75t_L g1717 ( 
.A1(n_1668),
.A2(n_1656),
.B(n_1648),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1692),
.A2(n_1650),
.B1(n_1624),
.B2(n_1646),
.C(n_1642),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1665),
.B(n_1639),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1692),
.B(n_1668),
.Y(n_1720)
);

NOR4xp25_ASAP7_75t_L g1721 ( 
.A(n_1670),
.B(n_1657),
.C(n_1662),
.D(n_1653),
.Y(n_1721)
);

AOI221x1_ASAP7_75t_L g1722 ( 
.A1(n_1670),
.A2(n_1657),
.B1(n_1637),
.B2(n_1638),
.C(n_1642),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1699),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1699),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1703),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1705),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1705),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1715),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1714),
.B(n_1665),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1700),
.A2(n_1667),
.B1(n_1666),
.B2(n_1695),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1715),
.B(n_1695),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1704),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1698),
.B(n_1676),
.Y(n_1733)
);

NAND2xp33_ASAP7_75t_L g1734 ( 
.A(n_1697),
.B(n_1695),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1709),
.Y(n_1735)
);

BUFx4f_ASAP7_75t_SL g1736 ( 
.A(n_1710),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1711),
.B(n_1666),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1719),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1711),
.B(n_1666),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1719),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1706),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1720),
.B(n_1703),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1712),
.B(n_1666),
.Y(n_1743)
);

NOR2x1_ASAP7_75t_L g1744 ( 
.A(n_1728),
.B(n_1712),
.Y(n_1744)
);

O2A1O1Ixp5_ASAP7_75t_SL g1745 ( 
.A1(n_1741),
.A2(n_1672),
.B(n_1694),
.C(n_1681),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1729),
.B(n_1701),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1730),
.A2(n_1702),
.B1(n_1716),
.B2(n_1732),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1730),
.B(n_1713),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1729),
.B(n_1713),
.Y(n_1749)
);

NAND2x1p5_ASAP7_75t_L g1750 ( 
.A(n_1738),
.B(n_1710),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1736),
.B(n_1701),
.Y(n_1751)
);

NOR3xp33_ASAP7_75t_L g1752 ( 
.A(n_1734),
.B(n_1742),
.C(n_1743),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1737),
.A2(n_1708),
.B(n_1706),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1725),
.B(n_1721),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1740),
.B(n_1707),
.Y(n_1755)
);

AOI222xp33_ASAP7_75t_L g1756 ( 
.A1(n_1736),
.A2(n_1718),
.B1(n_1717),
.B2(n_1707),
.C1(n_1686),
.C2(n_1672),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1755),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1744),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1746),
.B(n_1731),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1753),
.B(n_1739),
.Y(n_1760)
);

AOI211x1_ASAP7_75t_L g1761 ( 
.A1(n_1747),
.A2(n_1735),
.B(n_1727),
.C(n_1726),
.Y(n_1761)
);

A2O1A1Ixp33_ASAP7_75t_L g1762 ( 
.A1(n_1754),
.A2(n_1752),
.B(n_1748),
.C(n_1751),
.Y(n_1762)
);

NAND4xp25_ASAP7_75t_L g1763 ( 
.A(n_1756),
.B(n_1733),
.C(n_1722),
.D(n_1723),
.Y(n_1763)
);

NAND3xp33_ASAP7_75t_L g1764 ( 
.A(n_1745),
.B(n_1722),
.C(n_1724),
.Y(n_1764)
);

NOR3x1_ASAP7_75t_L g1765 ( 
.A(n_1749),
.B(n_1653),
.C(n_1627),
.Y(n_1765)
);

NAND4xp25_ASAP7_75t_L g1766 ( 
.A(n_1750),
.B(n_1685),
.C(n_1677),
.D(n_1686),
.Y(n_1766)
);

NAND3xp33_ASAP7_75t_SL g1767 ( 
.A(n_1762),
.B(n_1764),
.C(n_1760),
.Y(n_1767)
);

NAND3xp33_ASAP7_75t_L g1768 ( 
.A(n_1761),
.B(n_1763),
.C(n_1758),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1757),
.Y(n_1769)
);

NAND3xp33_ASAP7_75t_L g1770 ( 
.A(n_1766),
.B(n_1685),
.C(n_1681),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_L g1771 ( 
.A(n_1759),
.B(n_1685),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1765),
.B(n_1690),
.Y(n_1772)
);

AND3x2_ASAP7_75t_L g1773 ( 
.A(n_1769),
.B(n_1677),
.C(n_1688),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1768),
.B(n_1688),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1771),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1772),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1770),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1767),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1771),
.Y(n_1779)
);

NOR2x1_ASAP7_75t_L g1780 ( 
.A(n_1779),
.B(n_1685),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1774),
.A2(n_1678),
.B(n_1674),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1773),
.B(n_1677),
.Y(n_1782)
);

INVx5_ASAP7_75t_L g1783 ( 
.A(n_1775),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1777),
.Y(n_1784)
);

AND3x4_ASAP7_75t_L g1785 ( 
.A(n_1778),
.B(n_1678),
.C(n_1674),
.Y(n_1785)
);

XNOR2xp5_ASAP7_75t_L g1786 ( 
.A(n_1784),
.B(n_1776),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1782),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1783),
.B(n_1774),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1788),
.Y(n_1789)
);

NOR3xp33_ASAP7_75t_SL g1790 ( 
.A(n_1789),
.B(n_1787),
.C(n_1786),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1790),
.B(n_1783),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1790),
.B(n_1788),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1792),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1791),
.A2(n_1785),
.B1(n_1780),
.B2(n_1781),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1794),
.Y(n_1795)
);

AOI222xp33_ASAP7_75t_L g1796 ( 
.A1(n_1793),
.A2(n_1693),
.B1(n_1678),
.B2(n_1674),
.C1(n_1687),
.C2(n_1683),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1795),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1797),
.A2(n_1796),
.B1(n_1693),
.B2(n_1687),
.Y(n_1798)
);

OAI221xp5_ASAP7_75t_R g1799 ( 
.A1(n_1798),
.A2(n_1693),
.B1(n_1687),
.B2(n_1683),
.C(n_1676),
.Y(n_1799)
);

AOI211xp5_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1683),
.B(n_1647),
.C(n_1638),
.Y(n_1800)
);


endmodule