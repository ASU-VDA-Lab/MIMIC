module fake_jpeg_24976_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_46),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_18),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_29),
.B1(n_17),
.B2(n_35),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_50),
.A2(n_22),
.B1(n_21),
.B2(n_25),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_29),
.B1(n_17),
.B2(n_18),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_55),
.B1(n_63),
.B2(n_69),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_29),
.B1(n_18),
.B2(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_56),
.B(n_59),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_36),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_29),
.B1(n_16),
.B2(n_32),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_73),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_16),
.B1(n_23),
.B2(n_34),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_23),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_34),
.B1(n_26),
.B2(n_33),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_21),
.B1(n_22),
.B2(n_33),
.Y(n_90)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_81),
.Y(n_115)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

CKINVDCx6p67_ASAP7_75t_R g141 ( 
.A(n_76),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_48),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_102),
.Y(n_133)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_39),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_106),
.C(n_107),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_84),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_66),
.Y(n_84)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_89),
.A2(n_37),
.B1(n_26),
.B2(n_31),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_25),
.B1(n_67),
.B2(n_70),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_33),
.B1(n_22),
.B2(n_25),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_54),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_98),
.Y(n_131)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_0),
.B(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_107),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_56),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_101),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_61),
.B(n_21),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_66),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_105),
.B(n_109),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_40),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_40),
.Y(n_107)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_0),
.C(n_1),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_110),
.Y(n_125)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_40),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_44),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_42),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g137 ( 
.A(n_113),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_64),
.B1(n_67),
.B2(n_72),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_86),
.B1(n_106),
.B2(n_82),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_44),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_39),
.C(n_64),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_135),
.C(n_105),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_139),
.B1(n_140),
.B2(n_89),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_83),
.A2(n_26),
.B1(n_30),
.B2(n_27),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_82),
.B(n_39),
.Y(n_132)
);

NOR2x1p5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_112),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_100),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_42),
.C(n_44),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_80),
.A2(n_26),
.B1(n_30),
.B2(n_27),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_145),
.B(n_147),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_146),
.A2(n_148),
.B1(n_160),
.B2(n_175),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_124),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_98),
.B1(n_87),
.B2(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_149),
.B(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_115),
.B(n_87),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_100),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_151),
.B(n_166),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_163),
.B1(n_169),
.B2(n_141),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_76),
.Y(n_153)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_162),
.Y(n_210)
);

AO22x1_ASAP7_75t_L g201 ( 
.A1(n_156),
.A2(n_143),
.B1(n_114),
.B2(n_141),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_159),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_161),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_78),
.Y(n_159)
);

OAI22x1_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_96),
.B1(n_77),
.B2(n_42),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_77),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_88),
.B1(n_99),
.B2(n_111),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_168),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_167),
.C(n_174),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_133),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_95),
.C(n_44),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_123),
.A2(n_110),
.B1(n_104),
.B2(n_103),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_85),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_171),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_85),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_102),
.B(n_2),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_172),
.A2(n_173),
.B(n_138),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_44),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_79),
.C(n_93),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_79),
.B1(n_84),
.B2(n_37),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_31),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_133),
.B(n_136),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_117),
.A2(n_84),
.B1(n_31),
.B2(n_30),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_136),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_185),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_179),
.A2(n_203),
.B1(n_177),
.B2(n_173),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_193),
.B(n_4),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_117),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_120),
.C(n_125),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_167),
.C(n_174),
.Y(n_215)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_197),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_126),
.B1(n_141),
.B2(n_120),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_189),
.A2(n_199),
.B1(n_6),
.B2(n_7),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_126),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_5),
.Y(n_230)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_194),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_126),
.B(n_119),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_195),
.A2(n_209),
.B(n_15),
.Y(n_227)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_119),
.A3(n_138),
.B1(n_114),
.B2(n_129),
.Y(n_196)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_149),
.A2(n_141),
.B1(n_129),
.B2(n_143),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

AO22x1_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_143),
.B1(n_141),
.B2(n_92),
.Y(n_202)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_155),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_207),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_208),
.A2(n_168),
.B1(n_163),
.B2(n_164),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_144),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_213),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_210),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_214),
.B(n_216),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_219),
.C(n_223),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_217),
.Y(n_261)
);

AOI32xp33_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_144),
.A3(n_148),
.B1(n_165),
.B2(n_166),
.Y(n_218)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_158),
.C(n_146),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_173),
.B1(n_176),
.B2(n_162),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_222),
.B1(n_225),
.B2(n_233),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_1),
.C(n_3),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_230),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_236),
.Y(n_240)
);

OA21x2_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_5),
.B(n_6),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_201),
.B1(n_202),
.B2(n_209),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_5),
.C(n_6),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_183),
.C(n_187),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_194),
.A2(n_197),
.B1(n_179),
.B2(n_198),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_6),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_185),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_237),
.B1(n_207),
.B2(n_180),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_181),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_193),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_242),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_245),
.A2(n_251),
.B1(n_231),
.B2(n_211),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_205),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_247),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_224),
.A2(n_204),
.B1(n_201),
.B2(n_191),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_186),
.Y(n_254)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_228),
.Y(n_255)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_186),
.C(n_204),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_219),
.C(n_230),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_212),
.B(n_202),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_258),
.B(n_227),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_224),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_262),
.B(n_239),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_211),
.B1(n_220),
.B2(n_217),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_263),
.A2(n_277),
.B1(n_271),
.B2(n_262),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_266),
.C(n_268),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_221),
.C(n_234),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_249),
.C(n_256),
.Y(n_268)
);

XOR2x2_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_226),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_269),
.B(n_241),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_221),
.C(n_229),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_278),
.C(n_266),
.Y(n_290)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_195),
.B1(n_238),
.B2(n_184),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_240),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_199),
.B1(n_225),
.B2(n_236),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_203),
.C(n_12),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_283),
.A2(n_291),
.B1(n_292),
.B2(n_263),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_289),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_253),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_285),
.B(n_288),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_277),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_287),
.Y(n_300)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_267),
.B(n_275),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_243),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_264),
.C(n_279),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_252),
.B1(n_242),
.B2(n_239),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_295),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_269),
.A2(n_258),
.B(n_259),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_294),
.A2(n_240),
.B(n_284),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_265),
.B1(n_274),
.B2(n_255),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_308),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_302),
.C(n_304),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_303),
.B1(n_307),
.B2(n_250),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_272),
.C(n_276),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_245),
.B1(n_255),
.B2(n_254),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_290),
.C(n_289),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_292),
.A2(n_283),
.B1(n_293),
.B2(n_246),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_288),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_304),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_313),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_298),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_296),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_203),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_317),
.B(n_302),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_243),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_311),
.A2(n_309),
.B(n_300),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_318),
.A2(n_323),
.B(n_322),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_310),
.A2(n_305),
.B(n_309),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_250),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_314),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_313),
.A2(n_250),
.B(n_13),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_325),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_326),
.A2(n_320),
.B1(n_13),
.B2(n_14),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_11),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_328),
.C(n_327),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_13),
.C(n_14),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_14),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_14),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_15),
.Y(n_334)
);


endmodule