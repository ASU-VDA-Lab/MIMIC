module fake_jpeg_19559_n_95 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_49),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_51),
.Y(n_61)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_2),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_2),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_58),
.Y(n_70)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_42),
.B1(n_43),
.B2(n_41),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_64),
.B1(n_3),
.B2(n_4),
.Y(n_72)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_35),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_40),
.B1(n_45),
.B2(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_69),
.Y(n_75)
);

AND2x6_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_5),
.Y(n_78)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_7),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_45),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_3),
.Y(n_76)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_4),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_78),
.B1(n_68),
.B2(n_10),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_81),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_84),
.C(n_78),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_80),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_79),
.B(n_70),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_86),
.A2(n_75),
.B(n_85),
.Y(n_88)
);

OAI322xp33_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_87),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_89),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_8),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_23),
.B(n_24),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_27),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_31),
.C(n_32),
.Y(n_95)
);


endmodule