module fake_netlist_6_3362_n_843 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_843);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_843;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_772;
wire n_656;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_527;
wire n_608;
wire n_474;
wire n_683;
wire n_620;
wire n_420;
wire n_261;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_600;
wire n_464;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_120),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_5),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g172 ( 
.A(n_53),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_128),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_91),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_76),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_35),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_115),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_90),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_157),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_51),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_142),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_60),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_2),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_129),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_102),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_148),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_159),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_18),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_38),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_17),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_6),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_145),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_71),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_62),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_15),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_112),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_45),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_46),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_138),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_75),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_32),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_158),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_28),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_93),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_12),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_12),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_21),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_11),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_8),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_8),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_89),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_164),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_82),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_73),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_37),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_65),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_10),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_83),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_149),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_58),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_117),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_13),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_131),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_146),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_33),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_20),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_21),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_123),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_170),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_181),
.B(n_0),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_181),
.B(n_0),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_172),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_179),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_1),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_179),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_172),
.B(n_1),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_198),
.B(n_2),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_203),
.Y(n_254)
);

AND2x6_ASAP7_75t_L g255 ( 
.A(n_203),
.B(n_29),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_196),
.B(n_206),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_197),
.B(n_3),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_203),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_191),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_198),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_193),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_197),
.B(n_232),
.Y(n_267)
);

AND2x6_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_30),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_3),
.Y(n_269)
);

CKINVDCx6p67_ASAP7_75t_R g270 ( 
.A(n_172),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_185),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_185),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_230),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_31),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_168),
.B(n_171),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_174),
.B(n_4),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_211),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_228),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_176),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g280 ( 
.A(n_202),
.B(n_4),
.Y(n_280)
);

AND2x6_ASAP7_75t_L g281 ( 
.A(n_204),
.B(n_34),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g283 ( 
.A(n_213),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_210),
.B(n_5),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_217),
.B(n_6),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

AOI22x1_ASAP7_75t_SL g287 ( 
.A1(n_237),
.A2(n_215),
.B1(n_234),
.B2(n_224),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_L g288 ( 
.A1(n_249),
.A2(n_194),
.B1(n_235),
.B2(n_199),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_237),
.B(n_220),
.Y(n_289)
);

OR2x6_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_7),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_169),
.Y(n_292)
);

AND2x4_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_173),
.Y(n_293)
);

CKINVDCx8_ASAP7_75t_R g294 ( 
.A(n_262),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_271),
.A2(n_233),
.B1(n_231),
.B2(n_227),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_240),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_272),
.A2(n_226),
.B1(n_225),
.B2(n_223),
.Y(n_298)
);

AO22x2_ASAP7_75t_L g299 ( 
.A1(n_274),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_247),
.A2(n_222),
.B1(n_221),
.B2(n_219),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_175),
.Y(n_301)
);

AO22x2_ASAP7_75t_L g302 ( 
.A1(n_274),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_238),
.Y(n_305)
);

BUFx6f_ASAP7_75t_SL g306 ( 
.A(n_276),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_240),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_189),
.B1(n_208),
.B2(n_207),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_177),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_259),
.A2(n_218),
.B1(n_205),
.B2(n_201),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_266),
.B(n_178),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_180),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_283),
.A2(n_195),
.B1(n_192),
.B2(n_190),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_248),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_253),
.B(n_14),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_248),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_267),
.A2(n_188),
.B1(n_187),
.B2(n_184),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_248),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_L g324 ( 
.A1(n_270),
.A2(n_183),
.B1(n_182),
.B2(n_16),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_247),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_L g326 ( 
.A1(n_260),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_L g327 ( 
.A1(n_260),
.A2(n_259),
.B1(n_239),
.B2(n_242),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_273),
.B(n_36),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_263),
.B(n_39),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_276),
.B(n_19),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_243),
.A2(n_280),
.B1(n_269),
.B2(n_285),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_243),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_273),
.B(n_40),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_280),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_241),
.B(n_22),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_258),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_292),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_291),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_312),
.Y(n_340)
);

NOR2xp67_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_245),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_41),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_316),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_275),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_321),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_318),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_286),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_319),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_287),
.B(n_42),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_303),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_43),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_304),
.Y(n_354)
);

INVxp33_ASAP7_75t_L g355 ( 
.A(n_320),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_307),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_317),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_323),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_295),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_337),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_284),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_337),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_294),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_311),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_269),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_310),
.B(n_244),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_311),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_311),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_305),
.B(n_256),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_311),
.Y(n_370)
);

XOR2x2_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_24),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_305),
.B(n_256),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_309),
.B(n_250),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_310),
.B(n_251),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_334),
.Y(n_381)
);

XOR2x2_ASAP7_75t_L g382 ( 
.A(n_330),
.B(n_25),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_334),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_293),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_300),
.Y(n_385)
);

XNOR2x2_ASAP7_75t_L g386 ( 
.A(n_299),
.B(n_26),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_313),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_293),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

OR2x6_ASAP7_75t_L g390 ( 
.A(n_290),
.B(n_250),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_288),
.B(n_245),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_298),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_296),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_322),
.B(n_44),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_306),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_306),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_331),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_301),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_290),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_288),
.B(n_26),
.Y(n_400)
);

INVx4_ASAP7_75t_SL g401 ( 
.A(n_290),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_299),
.B(n_245),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_299),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_302),
.Y(n_404)
);

INVx4_ASAP7_75t_SL g405 ( 
.A(n_302),
.Y(n_405)
);

BUFx8_ASAP7_75t_L g406 ( 
.A(n_302),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_325),
.B(n_332),
.Y(n_407)
);

XNOR2x2_ASAP7_75t_L g408 ( 
.A(n_326),
.B(n_27),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_338),
.B(n_324),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_281),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_368),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_281),
.Y(n_412)
);

AND2x2_ASAP7_75t_SL g413 ( 
.A(n_361),
.B(n_365),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_373),
.B(n_281),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_374),
.B(n_281),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_375),
.B(n_281),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_377),
.B(n_255),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_387),
.B(n_336),
.Y(n_418)
);

AND2x2_ASAP7_75t_SL g419 ( 
.A(n_361),
.B(n_255),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_359),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_360),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_384),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_389),
.B(n_252),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_378),
.A2(n_255),
.B(n_268),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_362),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_379),
.B(n_255),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_351),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_370),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_398),
.B(n_255),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_352),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_268),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_354),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_356),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_390),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_381),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_339),
.B(n_268),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_364),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_357),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_345),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_344),
.B(n_268),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_383),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_405),
.B(n_365),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_338),
.B(n_399),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_344),
.B(n_268),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_363),
.Y(n_446)
);

OR2x6_ASAP7_75t_L g447 ( 
.A(n_390),
.B(n_326),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_340),
.B(n_245),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_363),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_405),
.B(n_380),
.Y(n_450)
);

AND2x2_ASAP7_75t_SL g451 ( 
.A(n_407),
.B(n_252),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_358),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_366),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_343),
.B(n_246),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_346),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_348),
.B(n_246),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_366),
.B(n_324),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_376),
.B(n_246),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_349),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_390),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_376),
.B(n_246),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_367),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_368),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_391),
.B(n_254),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_402),
.B(n_403),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_404),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_399),
.B(n_254),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_399),
.B(n_393),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_401),
.B(n_252),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_347),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_392),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_401),
.Y(n_472)
);

NAND2x1p5_ASAP7_75t_L g473 ( 
.A(n_341),
.B(n_254),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_401),
.B(n_252),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_391),
.B(n_265),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_386),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_342),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_395),
.B(n_254),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_396),
.B(n_47),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_406),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_397),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_432),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_446),
.B(n_355),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_413),
.B(n_355),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_455),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_443),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_413),
.B(n_400),
.Y(n_489)
);

AND2x6_ASAP7_75t_L g490 ( 
.A(n_432),
.B(n_406),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_426),
.B(n_385),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_449),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_413),
.B(n_419),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_419),
.B(n_394),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_470),
.B(n_385),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_420),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_420),
.Y(n_497)
);

OR2x6_ASAP7_75t_L g498 ( 
.A(n_447),
.B(n_408),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_455),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_436),
.B(n_353),
.Y(n_500)
);

OR2x6_ASAP7_75t_L g501 ( 
.A(n_447),
.B(n_477),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_421),
.Y(n_502)
);

INVx6_ASAP7_75t_L g503 ( 
.A(n_422),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_419),
.B(n_265),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_421),
.Y(n_505)
);

INVx8_ASAP7_75t_L g506 ( 
.A(n_432),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_425),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_465),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_476),
.B(n_350),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_466),
.B(n_265),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_466),
.B(n_265),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_425),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_463),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_443),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_463),
.Y(n_515)
);

NAND2x1p5_ASAP7_75t_L g516 ( 
.A(n_432),
.B(n_278),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_447),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_449),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_465),
.Y(n_519)
);

AND2x2_ASAP7_75t_SL g520 ( 
.A(n_451),
.B(n_278),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_423),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_462),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_436),
.B(n_27),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_423),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_462),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_428),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_428),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_429),
.Y(n_528)
);

AO21x2_ASAP7_75t_L g529 ( 
.A1(n_424),
.A2(n_48),
.B(n_49),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_478),
.B(n_50),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_451),
.B(n_278),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_478),
.B(n_52),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_410),
.B(n_278),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_426),
.B(n_54),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_481),
.B(n_55),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_479),
.B(n_56),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_431),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_422),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_431),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_442),
.Y(n_540)
);

AO21x2_ASAP7_75t_L g541 ( 
.A1(n_417),
.A2(n_57),
.B(n_59),
.Y(n_541)
);

INVxp67_ASAP7_75t_SL g542 ( 
.A(n_538),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_501),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_503),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_488),
.B(n_451),
.Y(n_545)
);

INVx3_ASAP7_75t_SL g546 ( 
.A(n_506),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_484),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_486),
.A2(n_457),
.B1(n_409),
.B2(n_468),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_515),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_515),
.Y(n_550)
);

INVx3_ASAP7_75t_SL g551 ( 
.A(n_506),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_497),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_484),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_512),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_538),
.Y(n_555)
);

INVx8_ASAP7_75t_L g556 ( 
.A(n_506),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_484),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_485),
.Y(n_558)
);

CKINVDCx14_ASAP7_75t_R g559 ( 
.A(n_518),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_483),
.B(n_471),
.Y(n_560)
);

INVx6_ASAP7_75t_SL g561 ( 
.A(n_501),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_492),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_484),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_512),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_497),
.Y(n_565)
);

BUFx12f_ASAP7_75t_L g566 ( 
.A(n_536),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_518),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_538),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_530),
.Y(n_569)
);

BUFx12f_ASAP7_75t_L g570 ( 
.A(n_491),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_496),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_488),
.B(n_422),
.Y(n_572)
);

BUFx4_ASAP7_75t_SL g573 ( 
.A(n_498),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_538),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_503),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_508),
.B(n_477),
.Y(n_576)
);

INVx3_ASAP7_75t_SL g577 ( 
.A(n_491),
.Y(n_577)
);

BUFx6f_ASAP7_75t_SL g578 ( 
.A(n_490),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_532),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_503),
.Y(n_580)
);

NAND2x1p5_ASAP7_75t_L g581 ( 
.A(n_535),
.B(n_528),
.Y(n_581)
);

BUFx8_ASAP7_75t_SL g582 ( 
.A(n_498),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_495),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_528),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_513),
.Y(n_585)
);

NAND2x1p5_ASAP7_75t_L g586 ( 
.A(n_535),
.B(n_438),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_501),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_514),
.Y(n_588)
);

BUFx2_ASAP7_75t_R g589 ( 
.A(n_494),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_560),
.A2(n_489),
.B1(n_471),
.B2(n_483),
.Y(n_590)
);

CKINVDCx12_ASAP7_75t_R g591 ( 
.A(n_576),
.Y(n_591)
);

BUFx10_ASAP7_75t_L g592 ( 
.A(n_578),
.Y(n_592)
);

INVx6_ASAP7_75t_L g593 ( 
.A(n_547),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_548),
.A2(n_498),
.B1(n_494),
.B2(n_493),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_585),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_576),
.B(n_508),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_545),
.B(n_519),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_545),
.A2(n_493),
.B1(n_517),
.B2(n_487),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_585),
.Y(n_599)
);

INVx6_ASAP7_75t_L g600 ( 
.A(n_547),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_554),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_574),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_549),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_554),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_549),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_582),
.A2(n_499),
.B1(n_520),
.B2(n_447),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_558),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_564),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_550),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_582),
.A2(n_520),
.B1(n_526),
.B2(n_539),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_569),
.A2(n_500),
.B1(n_444),
.B2(n_534),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_564),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_550),
.B(n_519),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_559),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_578),
.Y(n_615)
);

CKINVDCx11_ASAP7_75t_R g616 ( 
.A(n_570),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_583),
.B(n_579),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_588),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_588),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_546),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_552),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_570),
.A2(n_540),
.B1(n_534),
.B2(n_442),
.Y(n_622)
);

BUFx8_ASAP7_75t_L g623 ( 
.A(n_578),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_562),
.A2(n_509),
.B(n_418),
.Y(n_624)
);

BUFx6f_ASAP7_75t_SL g625 ( 
.A(n_567),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_574),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_567),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_SL g628 ( 
.A1(n_566),
.A2(n_523),
.B1(n_490),
.B2(n_482),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_552),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_SL g630 ( 
.A1(n_566),
.A2(n_490),
.B1(n_481),
.B2(n_410),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_543),
.A2(n_527),
.B1(n_537),
.B2(n_521),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_565),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_546),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_610),
.A2(n_587),
.B1(n_543),
.B2(n_577),
.Y(n_634)
);

BUFx12f_ASAP7_75t_L g635 ( 
.A(n_616),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_594),
.A2(n_587),
.B1(n_577),
.B2(n_422),
.Y(n_636)
);

AOI222xp33_ASAP7_75t_L g637 ( 
.A1(n_594),
.A2(n_577),
.B1(n_502),
.B2(n_505),
.C1(n_507),
.C2(n_481),
.Y(n_637)
);

OAI22xp33_ASAP7_75t_L g638 ( 
.A1(n_596),
.A2(n_561),
.B1(n_524),
.B2(n_571),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_610),
.A2(n_422),
.B1(n_561),
.B2(n_572),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_606),
.A2(n_561),
.B1(n_571),
.B2(n_572),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_606),
.A2(n_572),
.B1(n_434),
.B2(n_439),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_625),
.A2(n_412),
.B1(n_435),
.B2(n_460),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_625),
.A2(n_412),
.B1(n_459),
.B2(n_433),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_611),
.A2(n_586),
.B1(n_522),
.B2(n_525),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_622),
.A2(n_589),
.B1(n_586),
.B2(n_581),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_SL g646 ( 
.A1(n_590),
.A2(n_573),
.B1(n_490),
.B2(n_529),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_617),
.A2(n_459),
.B1(n_452),
.B2(n_433),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_591),
.B(n_467),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_595),
.Y(n_649)
);

BUFx4f_ASAP7_75t_SL g650 ( 
.A(n_623),
.Y(n_650)
);

BUFx4f_ASAP7_75t_SL g651 ( 
.A(n_623),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_607),
.A2(n_598),
.B1(n_627),
.B2(n_630),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_598),
.A2(n_452),
.B1(n_475),
.B2(n_434),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_618),
.A2(n_475),
.B1(n_439),
.B2(n_415),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_618),
.A2(n_416),
.B1(n_415),
.B2(n_529),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_628),
.A2(n_416),
.B1(n_430),
.B2(n_458),
.Y(n_656)
);

BUFx12f_ASAP7_75t_L g657 ( 
.A(n_616),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_SL g658 ( 
.A1(n_623),
.A2(n_614),
.B1(n_490),
.B2(n_619),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_619),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_631),
.A2(n_586),
.B1(n_581),
.B2(n_551),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_592),
.Y(n_661)
);

CKINVDCx11_ASAP7_75t_R g662 ( 
.A(n_592),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_597),
.B(n_565),
.Y(n_663)
);

OR2x6_ASAP7_75t_L g664 ( 
.A(n_620),
.B(n_556),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_624),
.A2(n_414),
.B1(n_480),
.B2(n_450),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_613),
.B(n_553),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_631),
.A2(n_461),
.B1(n_414),
.B2(n_440),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_SL g668 ( 
.A1(n_615),
.A2(n_581),
.B1(n_541),
.B2(n_531),
.Y(n_668)
);

OAI22xp33_ASAP7_75t_L g669 ( 
.A1(n_599),
.A2(n_531),
.B1(n_504),
.B2(n_551),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_601),
.B(n_450),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_604),
.A2(n_441),
.B(n_445),
.Y(n_671)
);

OAI21xp33_ASAP7_75t_L g672 ( 
.A1(n_608),
.A2(n_427),
.B(n_437),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_620),
.A2(n_472),
.B1(n_553),
.B2(n_469),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_615),
.A2(n_440),
.B1(n_557),
.B2(n_563),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_633),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_633),
.A2(n_546),
.B1(n_551),
.B2(n_504),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_603),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_593),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_612),
.B(n_557),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_SL g680 ( 
.A1(n_602),
.A2(n_541),
.B1(n_556),
.B2(n_574),
.Y(n_680)
);

BUFx12f_ASAP7_75t_L g681 ( 
.A(n_602),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_632),
.Y(n_682)
);

OAI22xp33_ASAP7_75t_L g683 ( 
.A1(n_603),
.A2(n_574),
.B1(n_510),
.B2(n_511),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_605),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_652),
.A2(n_553),
.B1(n_593),
.B2(n_600),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_682),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_637),
.A2(n_440),
.B1(n_563),
.B2(n_533),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_659),
.B(n_605),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_L g689 ( 
.A1(n_665),
.A2(n_602),
.B1(n_626),
.B2(n_575),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_641),
.A2(n_600),
.B1(n_593),
.B2(n_542),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_663),
.B(n_609),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_640),
.A2(n_533),
.B1(n_547),
.B2(n_469),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_640),
.A2(n_533),
.B1(n_547),
.B2(n_474),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_666),
.B(n_609),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_634),
.A2(n_533),
.B1(n_547),
.B2(n_474),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_679),
.B(n_621),
.Y(n_696)
);

AOI222xp33_ASAP7_75t_L g697 ( 
.A1(n_645),
.A2(n_464),
.B1(n_629),
.B2(n_621),
.C1(n_510),
.C2(n_511),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_649),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_641),
.A2(n_600),
.B1(n_555),
.B2(n_473),
.Y(n_699)
);

AOI221xp5_ASAP7_75t_L g700 ( 
.A1(n_644),
.A2(n_638),
.B1(n_642),
.B2(n_648),
.C(n_669),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_639),
.A2(n_533),
.B1(n_580),
.B2(n_438),
.Y(n_701)
);

OAI221xp5_ASAP7_75t_SL g702 ( 
.A1(n_646),
.A2(n_629),
.B1(n_544),
.B2(n_584),
.C(n_568),
.Y(n_702)
);

OAI222xp33_ASAP7_75t_L g703 ( 
.A1(n_636),
.A2(n_584),
.B1(n_544),
.B2(n_473),
.C1(n_516),
.C2(n_575),
.Y(n_703)
);

OAI221xp5_ASAP7_75t_L g704 ( 
.A1(n_643),
.A2(n_473),
.B1(n_516),
.B2(n_584),
.C(n_575),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_644),
.A2(n_580),
.B1(n_438),
.B2(n_556),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_656),
.A2(n_657),
.B1(n_635),
.B2(n_654),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_661),
.A2(n_580),
.B1(n_438),
.B2(n_556),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_677),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_684),
.B(n_568),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_SL g710 ( 
.A1(n_650),
.A2(n_626),
.B1(n_602),
.B2(n_574),
.Y(n_710)
);

AOI222xp33_ASAP7_75t_L g711 ( 
.A1(n_650),
.A2(n_651),
.B1(n_653),
.B2(n_647),
.C1(n_638),
.C2(n_670),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_683),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_651),
.A2(n_580),
.B1(n_438),
.B2(n_429),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_678),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_673),
.A2(n_411),
.B1(n_626),
.B2(n_568),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_658),
.A2(n_580),
.B1(n_429),
.B2(n_626),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_669),
.A2(n_429),
.B1(n_454),
.B2(n_448),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_662),
.A2(n_429),
.B1(n_456),
.B2(n_261),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_660),
.A2(n_261),
.B1(n_63),
.B2(n_64),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_667),
.A2(n_261),
.B1(n_66),
.B2(n_67),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_664),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_SL g722 ( 
.A1(n_676),
.A2(n_261),
.B1(n_68),
.B2(n_69),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_675),
.B(n_61),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_721),
.Y(n_724)
);

AOI21xp33_ASAP7_75t_L g725 ( 
.A1(n_711),
.A2(n_668),
.B(n_672),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_714),
.B(n_680),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_688),
.B(n_683),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_719),
.A2(n_664),
.B1(n_671),
.B2(n_681),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_700),
.B(n_674),
.C(n_655),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_691),
.B(n_664),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_686),
.B(n_714),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_686),
.B(n_70),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_694),
.B(n_72),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_721),
.B(n_167),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_696),
.B(n_698),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_689),
.B(n_702),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_698),
.B(n_74),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_708),
.B(n_77),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_708),
.B(n_78),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_709),
.B(n_79),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_719),
.B(n_80),
.C(n_81),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_706),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_697),
.B(n_87),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_704),
.B(n_88),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_709),
.B(n_92),
.Y(n_745)
);

OAI21xp5_ASAP7_75t_SL g746 ( 
.A1(n_722),
.A2(n_94),
.B(n_95),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_712),
.B(n_96),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_712),
.B(n_97),
.Y(n_748)
);

NOR3xp33_ASAP7_75t_L g749 ( 
.A(n_723),
.B(n_98),
.C(n_100),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_718),
.B(n_101),
.C(n_103),
.Y(n_750)
);

OA21x2_ASAP7_75t_L g751 ( 
.A1(n_717),
.A2(n_104),
.B(n_105),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_724),
.B(n_717),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_731),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_728),
.B(n_705),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_735),
.Y(n_755)
);

AO21x2_ASAP7_75t_L g756 ( 
.A1(n_743),
.A2(n_703),
.B(n_690),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_L g757 ( 
.A(n_743),
.B(n_685),
.C(n_699),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_724),
.B(n_695),
.Y(n_758)
);

NAND4xp75_ASAP7_75t_L g759 ( 
.A(n_751),
.B(n_710),
.C(n_716),
.D(n_707),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_724),
.B(n_693),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_729),
.A2(n_720),
.B1(n_692),
.B2(n_687),
.Y(n_761)
);

AND2x2_ASAP7_75t_SL g762 ( 
.A(n_751),
.B(n_701),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_SL g763 ( 
.A(n_736),
.B(n_715),
.Y(n_763)
);

AOI21xp33_ASAP7_75t_L g764 ( 
.A1(n_744),
.A2(n_713),
.B(n_107),
.Y(n_764)
);

NOR3xp33_ASAP7_75t_L g765 ( 
.A(n_741),
.B(n_106),
.C(n_108),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_730),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_727),
.B(n_109),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_753),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_766),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_755),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_766),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_752),
.B(n_726),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_752),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_758),
.Y(n_774)
);

INVx4_ASAP7_75t_L g775 ( 
.A(n_756),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_760),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_767),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_760),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_762),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_774),
.B(n_756),
.Y(n_780)
);

XNOR2xp5_ASAP7_75t_L g781 ( 
.A(n_777),
.B(n_759),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_769),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_768),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_773),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_769),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_783),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_784),
.Y(n_787)
);

OA22x2_ASAP7_75t_L g788 ( 
.A1(n_781),
.A2(n_775),
.B1(n_779),
.B2(n_776),
.Y(n_788)
);

AO22x2_ASAP7_75t_L g789 ( 
.A1(n_780),
.A2(n_775),
.B1(n_779),
.B2(n_778),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_782),
.A2(n_754),
.B1(n_775),
.B2(n_762),
.Y(n_790)
);

OA22x2_ASAP7_75t_L g791 ( 
.A1(n_782),
.A2(n_772),
.B1(n_773),
.B2(n_754),
.Y(n_791)
);

XOR2xp5_ASAP7_75t_L g792 ( 
.A(n_784),
.B(n_742),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_787),
.Y(n_793)
);

OAI322xp33_ASAP7_75t_L g794 ( 
.A1(n_788),
.A2(n_790),
.A3(n_791),
.B1(n_786),
.B2(n_763),
.C1(n_792),
.C2(n_770),
.Y(n_794)
);

XOR2xp5_ASAP7_75t_L g795 ( 
.A(n_789),
.B(n_750),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_789),
.Y(n_796)
);

OAI322xp33_ASAP7_75t_L g797 ( 
.A1(n_788),
.A2(n_770),
.A3(n_768),
.B1(n_736),
.B2(n_785),
.C1(n_744),
.C2(n_728),
.Y(n_797)
);

OAI322xp33_ASAP7_75t_L g798 ( 
.A1(n_788),
.A2(n_772),
.A3(n_771),
.B1(n_747),
.B2(n_748),
.C1(n_733),
.C2(n_745),
.Y(n_798)
);

AOI221xp5_ASAP7_75t_L g799 ( 
.A1(n_794),
.A2(n_757),
.B1(n_725),
.B2(n_764),
.C(n_765),
.Y(n_799)
);

OA22x2_ASAP7_75t_L g800 ( 
.A1(n_795),
.A2(n_746),
.B1(n_734),
.B2(n_737),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_796),
.A2(n_749),
.B1(n_751),
.B2(n_761),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_800),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_801),
.A2(n_793),
.B1(n_797),
.B2(n_761),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_799),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_802),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_803),
.B(n_798),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_804),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_803),
.B(n_740),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_802),
.Y(n_809)
);

OA22x2_ASAP7_75t_L g810 ( 
.A1(n_804),
.A2(n_732),
.B1(n_739),
.B2(n_738),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_805),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_809),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_807),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_806),
.A2(n_808),
.B1(n_810),
.B2(n_113),
.Y(n_814)
);

NOR2x1_ASAP7_75t_L g815 ( 
.A(n_807),
.B(n_110),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_805),
.B(n_111),
.Y(n_816)
);

AOI211xp5_ASAP7_75t_SL g817 ( 
.A1(n_811),
.A2(n_114),
.B(n_116),
.C(n_118),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_815),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_814),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_819)
);

NAND2x1_ASAP7_75t_L g820 ( 
.A(n_812),
.B(n_124),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_813),
.A2(n_126),
.B1(n_127),
.B2(n_130),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_818),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_820),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_821),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_819),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_817),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_820),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_818),
.B(n_816),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_822),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_823),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_828),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_826),
.A2(n_825),
.B1(n_824),
.B2(n_827),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_828),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_833)
);

OAI22x1_ASAP7_75t_L g834 ( 
.A1(n_823),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_830),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_831),
.Y(n_836)
);

OAI22xp33_ASAP7_75t_L g837 ( 
.A1(n_836),
.A2(n_832),
.B1(n_829),
.B2(n_833),
.Y(n_837)
);

NAND4xp25_ASAP7_75t_L g838 ( 
.A(n_835),
.B(n_834),
.C(n_140),
.D(n_141),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_838),
.Y(n_839)
);

OAI22xp33_ASAP7_75t_L g840 ( 
.A1(n_839),
.A2(n_837),
.B1(n_143),
.B2(n_147),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_840),
.Y(n_841)
);

AOI221xp5_ASAP7_75t_L g842 ( 
.A1(n_841),
.A2(n_139),
.B1(n_150),
.B2(n_151),
.C(n_152),
.Y(n_842)
);

AOI211xp5_ASAP7_75t_L g843 ( 
.A1(n_842),
.A2(n_153),
.B(n_154),
.C(n_155),
.Y(n_843)
);


endmodule