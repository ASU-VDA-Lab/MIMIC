module fake_jpeg_13157_n_587 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_587);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_587;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_2),
.B(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_57),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g176 ( 
.A(n_65),
.Y(n_176)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_9),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_67),
.B(n_68),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_32),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_78),
.Y(n_159)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_81),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_82),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_83),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_84),
.Y(n_189)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_85),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_87),
.Y(n_193)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_89),
.Y(n_198)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_92),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_95),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_98),
.Y(n_191)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_22),
.B(n_15),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_100),
.B(n_105),
.Y(n_154)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_22),
.B(n_15),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_123),
.Y(n_142)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_103),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_24),
.B(n_15),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_20),
.Y(n_106)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_20),
.Y(n_110)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_24),
.B(n_14),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_111),
.B(n_118),
.Y(n_170)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_26),
.Y(n_112)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_27),
.B(n_14),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_115),
.B(n_116),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_27),
.B(n_14),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_31),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_39),
.Y(n_120)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_23),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_62),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_125),
.A2(n_148),
.B1(n_152),
.B2(n_160),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_85),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_128),
.B(n_150),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_60),
.A2(n_35),
.B1(n_34),
.B2(n_42),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_135),
.A2(n_31),
.B(n_89),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_61),
.A2(n_35),
.B1(n_28),
.B2(n_23),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_101),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_151),
.B(n_123),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_77),
.A2(n_47),
.B1(n_23),
.B2(n_28),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_110),
.A2(n_47),
.B1(n_23),
.B2(n_28),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_63),
.A2(n_28),
.B1(n_52),
.B2(n_47),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_162),
.A2(n_87),
.B1(n_92),
.B2(n_96),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_37),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_166),
.B(n_178),
.Y(n_256)
);

OA22x2_ASAP7_75t_SL g171 ( 
.A1(n_65),
.A2(n_42),
.B1(n_41),
.B2(n_43),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_171),
.B(n_184),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_93),
.A2(n_52),
.B1(n_47),
.B2(n_98),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_172),
.A2(n_184),
.B1(n_188),
.B2(n_199),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_83),
.B(n_32),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_106),
.B(n_48),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_41),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_70),
.A2(n_52),
.B1(n_58),
.B2(n_53),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_71),
.A2(n_37),
.B1(n_43),
.B2(n_52),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_75),
.B(n_25),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_192),
.B(n_196),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_76),
.B(n_25),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_80),
.A2(n_49),
.B1(n_48),
.B2(n_39),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_81),
.B(n_58),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_203),
.B(n_1),
.Y(n_273)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_204),
.Y(n_290)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_206),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_175),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_207),
.B(n_242),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_49),
.B1(n_51),
.B2(n_56),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_208),
.A2(n_224),
.B1(n_247),
.B2(n_249),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_131),
.B(n_144),
.C(n_155),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_209),
.B(n_217),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_210),
.Y(n_291)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_213),
.B(n_238),
.Y(n_298)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_214),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_215),
.B(n_230),
.Y(n_302)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_216),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_51),
.C(n_119),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_219),
.Y(n_293)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_220),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_221),
.A2(n_236),
.B1(n_271),
.B2(n_160),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_222),
.Y(n_309)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_223),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_129),
.A2(n_46),
.B1(n_56),
.B2(n_53),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_170),
.B(n_46),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_225),
.B(n_239),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_142),
.B(n_0),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_L g284 ( 
.A1(n_226),
.A2(n_245),
.B(n_273),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_227),
.A2(n_5),
.B(n_6),
.Y(n_316)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_130),
.Y(n_228)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_228),
.Y(n_282)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_231),
.Y(n_283)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_232),
.Y(n_310)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_233),
.Y(n_314)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_134),
.Y(n_234)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_234),
.Y(n_317)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_235),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_180),
.A2(n_104),
.B1(n_121),
.B2(n_114),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_127),
.A2(n_113),
.B1(n_109),
.B2(n_107),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_237),
.A2(n_267),
.B1(n_167),
.B2(n_149),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_175),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_89),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_141),
.Y(n_240)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_240),
.Y(n_329)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_241),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

INVx4_ASAP7_75t_SL g243 ( 
.A(n_164),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_243),
.B(n_246),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_140),
.Y(n_244)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_244),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_156),
.B(n_0),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_159),
.B(n_1),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_129),
.A2(n_84),
.B1(n_83),
.B2(n_82),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_165),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_250),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_157),
.A2(n_84),
.B1(n_31),
.B2(n_10),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_134),
.Y(n_251)
);

BUFx6f_ASAP7_75t_SL g332 ( 
.A(n_251),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_252),
.Y(n_301)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_190),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_253),
.B(n_257),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_145),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_254),
.Y(n_318)
);

AOI32xp33_ASAP7_75t_L g255 ( 
.A1(n_154),
.A2(n_31),
.A3(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_255),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_138),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_161),
.B(n_12),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_258),
.B(n_264),
.Y(n_289)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_146),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_259),
.Y(n_322)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_146),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_260),
.B(n_261),
.Y(n_319)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_187),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_262),
.B(n_263),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_199),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_148),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_163),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_265),
.A2(n_269),
.B1(n_274),
.B2(n_147),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_152),
.A2(n_31),
.B1(n_11),
.B2(n_4),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_133),
.B(n_1),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_4),
.Y(n_311)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_198),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_168),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_270),
.B(n_272),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_167),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_140),
.B(n_11),
.Y(n_272)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_181),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_275),
.A2(n_278),
.B1(n_279),
.B2(n_292),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_229),
.A2(n_149),
.B1(n_136),
.B2(n_133),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_212),
.A2(n_136),
.B1(n_197),
.B2(n_139),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_280),
.A2(n_215),
.B1(n_230),
.B2(n_245),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_263),
.A2(n_158),
.B1(n_193),
.B2(n_186),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_300),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_L g303 ( 
.A1(n_256),
.A2(n_172),
.B(n_3),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_L g353 ( 
.A1(n_303),
.A2(n_308),
.B(n_5),
.Y(n_353)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_266),
.B(n_177),
.CI(n_168),
.CON(n_304),
.SN(n_304)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_304),
.B(n_313),
.Y(n_355)
);

AND2x2_ASAP7_75t_SL g306 ( 
.A(n_246),
.B(n_191),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_307),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_242),
.A2(n_139),
.B(n_193),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_311),
.B(n_268),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g313 ( 
.A(n_209),
.B(n_194),
.CI(n_197),
.CON(n_313),
.SN(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_226),
.B(n_153),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_323),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_231),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_226),
.B(n_153),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_246),
.B(n_137),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_325),
.B(n_7),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_210),
.A2(n_186),
.B1(n_137),
.B2(n_158),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_327),
.A2(n_221),
.B1(n_232),
.B2(n_205),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_227),
.A2(n_185),
.B1(n_6),
.B2(n_7),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_328),
.A2(n_243),
.B(n_7),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_218),
.B(n_185),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_330),
.B(n_285),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_333),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_334),
.B(n_346),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_335),
.A2(n_341),
.B1(n_358),
.B2(n_367),
.Y(n_405)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_337),
.A2(n_342),
.B1(n_356),
.B2(n_357),
.Y(n_377)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_338),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_287),
.B(n_215),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_340),
.B(n_370),
.C(n_326),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_278),
.A2(n_217),
.B1(n_240),
.B2(n_241),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_302),
.A2(n_245),
.B1(n_248),
.B2(n_250),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_314),
.Y(n_343)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_309),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_344),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_288),
.B(n_265),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_345),
.B(n_349),
.Y(n_396)
);

AO22x1_ASAP7_75t_SL g346 ( 
.A1(n_302),
.A2(n_220),
.B1(n_233),
.B2(n_235),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_274),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_347),
.B(n_294),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_348),
.A2(n_354),
.B1(n_310),
.B2(n_324),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_305),
.B(n_252),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_286),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_361),
.Y(n_378)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_297),
.Y(n_352)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_353),
.A2(n_310),
.B1(n_331),
.B2(n_324),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_280),
.A2(n_244),
.B1(n_214),
.B2(n_260),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_289),
.A2(n_228),
.B1(n_204),
.B2(n_206),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_291),
.A2(n_216),
.B1(n_234),
.B2(n_251),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_279),
.A2(n_270),
.B1(n_259),
.B2(n_269),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_309),
.Y(n_394)
);

A2O1A1Ixp33_ASAP7_75t_SL g360 ( 
.A1(n_295),
.A2(n_6),
.B(n_7),
.C(n_222),
.Y(n_360)
);

O2A1O1Ixp33_ASAP7_75t_L g387 ( 
.A1(n_360),
.A2(n_332),
.B(n_322),
.C(n_301),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_296),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_362),
.B(n_365),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_311),
.B(n_287),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_306),
.A2(n_320),
.B1(n_325),
.B2(n_284),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_366),
.A2(n_374),
.B1(n_318),
.B2(n_322),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_328),
.A2(n_275),
.B1(n_321),
.B2(n_316),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_313),
.B(n_323),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_372),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_313),
.A2(n_304),
.B1(n_292),
.B2(n_327),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_369),
.A2(n_355),
.B1(n_367),
.B2(n_339),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_306),
.B(n_320),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_371),
.B(n_334),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_315),
.B(n_304),
.Y(n_372)
);

INVx13_ASAP7_75t_L g373 ( 
.A(n_276),
.Y(n_373)
);

BUFx5_ASAP7_75t_L g407 ( 
.A(n_373),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_320),
.A2(n_307),
.B1(n_308),
.B2(n_293),
.Y(n_374)
);

AO22x1_ASAP7_75t_SL g375 ( 
.A1(n_293),
.A2(n_312),
.B1(n_277),
.B2(n_329),
.Y(n_375)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_375),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_331),
.A2(n_276),
.B1(n_318),
.B2(n_298),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_376),
.A2(n_283),
.B(n_294),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_368),
.A2(n_277),
.B1(n_319),
.B2(n_317),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_381),
.A2(n_395),
.B1(n_398),
.B2(n_335),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_382),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_383),
.A2(n_390),
.B(n_394),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_312),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_340),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_386),
.Y(n_446)
);

OR2x6_ASAP7_75t_SL g427 ( 
.A(n_387),
.B(n_400),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_376),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_397),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_361),
.B(n_329),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_389),
.B(n_409),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_339),
.A2(n_283),
.B(n_299),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_392),
.A2(n_359),
.B(n_348),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_374),
.A2(n_290),
.B1(n_317),
.B2(n_282),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_375),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_372),
.A2(n_290),
.B1(n_282),
.B2(n_281),
.Y(n_398)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_375),
.Y(n_403)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_403),
.Y(n_434)
);

AOI21xp33_ASAP7_75t_SL g404 ( 
.A1(n_347),
.A2(n_299),
.B(n_326),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_SL g423 ( 
.A(n_404),
.B(n_412),
.C(n_347),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_336),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_411),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_385),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_351),
.B(n_281),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_343),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_413),
.A2(n_355),
.B1(n_366),
.B2(n_348),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_415),
.B(n_379),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_418),
.A2(n_438),
.B1(n_441),
.B2(n_377),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_420),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_386),
.A2(n_369),
.B1(n_363),
.B2(n_339),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_421),
.A2(n_424),
.B1(n_433),
.B2(n_444),
.Y(n_448)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_407),
.Y(n_422)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_423),
.A2(n_418),
.B1(n_432),
.B2(n_442),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_401),
.A2(n_363),
.B1(n_341),
.B2(n_358),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_350),
.Y(n_425)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_425),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_350),
.Y(n_426)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_426),
.Y(n_466)
);

AOI21x1_ASAP7_75t_L g468 ( 
.A1(n_429),
.A2(n_400),
.B(n_380),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_436),
.Y(n_453)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_410),
.Y(n_431)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_431),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_378),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_432),
.B(n_437),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_403),
.A2(n_364),
.B1(n_362),
.B2(n_360),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_352),
.Y(n_435)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_435),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_408),
.B(n_370),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_378),
.B(n_338),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_405),
.A2(n_342),
.B1(n_356),
.B2(n_357),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_346),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_439),
.B(n_384),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_405),
.A2(n_346),
.B1(n_360),
.B2(n_344),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_389),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_442),
.B(n_443),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_406),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_388),
.A2(n_360),
.B1(n_333),
.B2(n_373),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_445),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_377),
.A2(n_333),
.B1(n_360),
.B2(n_381),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_447),
.A2(n_390),
.B1(n_383),
.B2(n_394),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_449),
.A2(n_459),
.B1(n_469),
.B2(n_427),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_450),
.A2(n_455),
.B1(n_458),
.B2(n_472),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_452),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_446),
.A2(n_395),
.B1(n_384),
.B2(n_387),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_440),
.A2(n_387),
.B1(n_412),
.B2(n_396),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_421),
.A2(n_413),
.B1(n_394),
.B2(n_392),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_461),
.B(n_428),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_437),
.B(n_396),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_462),
.B(n_467),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_463),
.B(n_465),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_436),
.B(n_379),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_419),
.B(n_399),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_468),
.A2(n_475),
.B(n_416),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_434),
.A2(n_393),
.B1(n_399),
.B2(n_411),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_419),
.B(n_407),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_470),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_441),
.A2(n_393),
.B1(n_414),
.B2(n_391),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_430),
.B(n_391),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_415),
.C(n_423),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_416),
.A2(n_414),
.B(n_410),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_434),
.A2(n_402),
.B1(n_410),
.B2(n_438),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_476),
.A2(n_420),
.B1(n_447),
.B2(n_424),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_450),
.A2(n_451),
.B1(n_455),
.B2(n_464),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_477),
.A2(n_489),
.B1(n_466),
.B2(n_474),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_491),
.Y(n_509)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_457),
.Y(n_483)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_483),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_473),
.B(n_422),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_484),
.B(n_502),
.Y(n_506)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_454),
.Y(n_486)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_486),
.Y(n_504)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_454),
.Y(n_487)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_487),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_488),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_490),
.B(n_472),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_469),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_453),
.B(n_426),
.C(n_425),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_496),
.C(n_465),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_464),
.B(n_443),
.Y(n_493)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_493),
.Y(n_514)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_460),
.Y(n_494)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_494),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_495),
.B(n_468),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_435),
.C(n_429),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_448),
.A2(n_451),
.B1(n_449),
.B2(n_459),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_497),
.B(n_499),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_471),
.Y(n_498)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_498),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_458),
.A2(n_427),
.B(n_428),
.Y(n_499)
);

FAx1_ASAP7_75t_L g500 ( 
.A(n_461),
.B(n_427),
.CI(n_448),
.CON(n_500),
.SN(n_500)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_500),
.B(n_501),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_466),
.B(n_417),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_452),
.B(n_445),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_505),
.B(n_508),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_507),
.B(n_517),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_496),
.Y(n_508)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_494),
.Y(n_511)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_511),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_513),
.A2(n_516),
.B1(n_521),
.B2(n_486),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_489),
.A2(n_474),
.B1(n_439),
.B2(n_427),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_490),
.B(n_463),
.C(n_475),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_518),
.B(n_519),
.C(n_523),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_482),
.B(n_476),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_492),
.B(n_417),
.C(n_433),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_503),
.B(n_480),
.Y(n_525)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_525),
.Y(n_553)
);

A2O1A1Ixp33_ASAP7_75t_SL g527 ( 
.A1(n_522),
.A2(n_499),
.B(n_500),
.C(n_488),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_527),
.B(n_520),
.C(n_479),
.Y(n_549)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_506),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_529),
.Y(n_541)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_515),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_521),
.A2(n_478),
.B1(n_477),
.B2(n_491),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_530),
.B(n_534),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_510),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_493),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_507),
.B(n_485),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_504),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_535),
.B(n_536),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_518),
.B(n_495),
.C(n_497),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_512),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_L g550 ( 
.A(n_537),
.B(n_540),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_538),
.A2(n_478),
.B1(n_520),
.B2(n_522),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_514),
.B(n_480),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_539),
.A2(n_483),
.B(n_501),
.Y(n_547)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_510),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_542),
.B(n_546),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_531),
.B(n_519),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_544),
.B(n_545),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_531),
.B(n_508),
.Y(n_545)
);

AOI21x1_ASAP7_75t_L g564 ( 
.A1(n_547),
.A2(n_549),
.B(n_539),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_538),
.A2(n_517),
.B1(n_523),
.B2(n_500),
.Y(n_551)
);

OAI21xp33_ASAP7_75t_L g558 ( 
.A1(n_551),
.A2(n_509),
.B(n_500),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_532),
.B(n_513),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_552),
.B(n_554),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_526),
.A2(n_509),
.B(n_481),
.Y(n_554)
);

AOI21x1_ASAP7_75t_SL g573 ( 
.A1(n_558),
.A2(n_559),
.B(n_546),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_553),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_548),
.B(n_532),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_560),
.B(n_561),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_551),
.B(n_536),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_552),
.B(n_530),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_562),
.B(n_542),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_527),
.C(n_533),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_563),
.B(n_565),
.Y(n_566)
);

OAI21xp33_ASAP7_75t_L g571 ( 
.A1(n_564),
.A2(n_487),
.B(n_527),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_541),
.B(n_525),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_557),
.B(n_549),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_567),
.B(n_572),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_559),
.A2(n_545),
.B(n_550),
.Y(n_568)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_568),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_570),
.B(n_573),
.Y(n_574)
);

A2O1A1O1Ixp25_ASAP7_75t_L g578 ( 
.A1(n_571),
.A2(n_558),
.B(n_505),
.C(n_516),
.D(n_524),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_555),
.B(n_544),
.C(n_527),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_569),
.B(n_555),
.C(n_556),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_576),
.B(n_566),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_578),
.A2(n_566),
.B(n_511),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_579),
.A2(n_580),
.B(n_581),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_575),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_580),
.B(n_574),
.C(n_577),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g584 ( 
.A1(n_582),
.A2(n_574),
.B(n_456),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_584),
.B(n_583),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_585),
.A2(n_460),
.B(n_471),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_586),
.A2(n_431),
.B(n_444),
.Y(n_587)
);


endmodule