module fake_jpeg_3941_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_49),
.Y(n_60)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_30),
.B1(n_26),
.B2(n_23),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_30),
.B1(n_26),
.B2(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_56),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_62),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_64),
.B(n_66),
.Y(n_94)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_67),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_73),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_40),
.B1(n_34),
.B2(n_35),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_17),
.B1(n_32),
.B2(n_28),
.Y(n_95)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_71),
.B(n_75),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_24),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_74),
.B(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_26),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_25),
.C(n_17),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_24),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_18),
.Y(n_84)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_60),
.CI(n_59),
.CON(n_109),
.SN(n_109)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_25),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_37),
.B1(n_36),
.B2(n_38),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_62),
.B1(n_32),
.B2(n_22),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_114),
.B1(n_16),
.B2(n_21),
.Y(n_119)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_37),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_SL g141 ( 
.A(n_98),
.B(n_101),
.C(n_105),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_73),
.C(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_109),
.B(n_22),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_17),
.B1(n_16),
.B2(n_28),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_134),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_61),
.C(n_57),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_139),
.C(n_58),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_76),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_113),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_21),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_123),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_119),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_82),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_121),
.B(n_138),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_78),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_70),
.Y(n_122)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_90),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_111),
.B1(n_110),
.B2(n_103),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_18),
.B1(n_29),
.B2(n_72),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_130),
.A2(n_132),
.B1(n_114),
.B2(n_97),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_27),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_135),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_89),
.A2(n_82),
.B1(n_27),
.B2(n_20),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_99),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_25),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_80),
.C(n_58),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_25),
.C(n_15),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_100),
.B(n_110),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_145),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_153),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_96),
.B(n_113),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_156),
.B(n_157),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_130),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_104),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_120),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_103),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_155),
.Y(n_181)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_100),
.B(n_92),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_124),
.A2(n_27),
.B(n_20),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_108),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_161),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_80),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_3),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_132),
.C(n_118),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_20),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_13),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_169),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_172),
.C(n_174),
.Y(n_204)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_188),
.Y(n_198)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_134),
.C(n_138),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_138),
.C(n_125),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_0),
.B(n_1),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_112),
.B1(n_111),
.B2(n_15),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_177),
.A2(n_143),
.B1(n_148),
.B2(n_163),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_149),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_2),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_146),
.Y(n_196)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_4),
.Y(n_189)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_161),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_203),
.Y(n_213)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

OA21x2_ASAP7_75t_SL g201 ( 
.A1(n_170),
.A2(n_160),
.B(n_147),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_166),
.A3(n_5),
.B1(n_6),
.B2(n_9),
.C1(n_4),
.C2(n_11),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_164),
.B(n_144),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_167),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_205),
.Y(n_212)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_184),
.B1(n_171),
.B2(n_188),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_216),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_181),
.B1(n_168),
.B2(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_211),
.B(n_215),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_198),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_172),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_175),
.B1(n_183),
.B2(n_174),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_217),
.Y(n_230)
);

A2O1A1O1Ixp25_ASAP7_75t_L g218 ( 
.A1(n_203),
.A2(n_156),
.B(n_157),
.C(n_176),
.D(n_154),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_218),
.B(n_5),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_205),
.B(n_196),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_220),
.A2(n_193),
.B1(n_200),
.B2(n_192),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_204),
.C(n_194),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_231),
.C(n_213),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_202),
.B(n_195),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_225),
.B(n_226),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_209),
.A2(n_191),
.B1(n_204),
.B2(n_194),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_228),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_4),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_R g233 ( 
.A(n_224),
.B(n_218),
.C(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_207),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_238),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_222),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_223),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_239),
.C(n_221),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_212),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_208),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_216),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_233),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_214),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_243),
.B(n_244),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_230),
.Y(n_244)
);

AOI31xp67_ASAP7_75t_SL g252 ( 
.A1(n_246),
.A2(n_248),
.A3(n_247),
.B(n_9),
.Y(n_252)
);

INVxp33_ASAP7_75t_SL g251 ( 
.A(n_247),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_237),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_249),
.A2(n_241),
.B1(n_240),
.B2(n_225),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_252),
.C(n_6),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_253),
.A2(n_254),
.B(n_10),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_251),
.A2(n_6),
.B(n_10),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_11),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_11),
.Y(n_257)
);


endmodule