module fake_jpeg_28487_n_163 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

INVx8_ASAP7_75t_SL g66 ( 
.A(n_16),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_77),
.Y(n_90)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_0),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_64),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_0),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_57),
.B(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_67),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_54),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_58),
.B1(n_51),
.B2(n_65),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_88),
.B1(n_91),
.B2(n_54),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_93),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_64),
.B1(n_51),
.B2(n_65),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_47),
.B1(n_49),
.B2(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_66),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_100),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

AO22x1_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_69),
.B1(n_54),
.B2(n_60),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_109),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_108),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_3),
.B(n_6),
.Y(n_125)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_63),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_1),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_61),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_59),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_56),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_2),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_128),
.Y(n_134)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_122),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_25),
.B(n_27),
.Y(n_140)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_6),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_7),
.B1(n_14),
.B2(n_17),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_142),
.B1(n_34),
.B2(n_36),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_132),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_139),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_40),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_142),
.C(n_141),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_24),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_140),
.A2(n_118),
.B(n_35),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_28),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_117),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_37),
.Y(n_153)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_149),
.C(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_150),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_114),
.B(n_123),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_152),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_153),
.A2(n_38),
.B1(n_116),
.B2(n_115),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_154),
.C(n_151),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_157),
.A2(n_156),
.B1(n_136),
.B2(n_135),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_144),
.B(n_145),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_134),
.CI(n_147),
.CON(n_160),
.SN(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_160),
.Y(n_162)
);

NOR2xp67_ASAP7_75t_R g163 ( 
.A(n_162),
.B(n_149),
.Y(n_163)
);


endmodule