module fake_jpeg_21810_n_69 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_69);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_69;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_55;
wire n_27;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_24;
wire n_28;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_25;
wire n_67;
wire n_43;
wire n_29;
wire n_50;
wire n_37;
wire n_32;
wire n_66;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_6),
.B(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_49)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_3),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

NOR3xp33_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_50),
.C(n_53),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_35),
.B2(n_36),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_53),
.C(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_58),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_34),
.B1(n_24),
.B2(n_39),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_25),
.C(n_18),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_18),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_62),
.C(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_63),
.B(n_6),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_32),
.B(n_27),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_33),
.C(n_23),
.Y(n_66)
);

OAI321xp33_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_66),
.A3(n_48),
.B1(n_49),
.B2(n_28),
.C(n_23),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_38),
.B1(n_44),
.B2(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_45),
.Y(n_69)
);


endmodule