module fake_aes_6464_n_25 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_25);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
NOR2x1p5_ASAP7_75t_L g9 ( .A(n_8), .B(n_4), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_6), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_3), .Y(n_11) );
BUFx2_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_14), .B(n_0), .Y(n_15) );
CKINVDCx16_ASAP7_75t_R g16 ( .A(n_15), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_16), .B(n_12), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_17), .B(n_12), .Y(n_19) );
AOI21xp33_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_18), .B(n_10), .Y(n_20) );
O2A1O1Ixp33_ASAP7_75t_L g21 ( .A1(n_18), .A2(n_11), .B(n_13), .C(n_9), .Y(n_21) );
CKINVDCx16_ASAP7_75t_R g22 ( .A(n_20), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
OAI22xp5_ASAP7_75t_SL g24 ( .A1(n_22), .A2(n_11), .B1(n_10), .B2(n_14), .Y(n_24) );
AOI222xp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_23), .B1(n_1), .B2(n_2), .C1(n_3), .C2(n_0), .Y(n_25) );
endmodule