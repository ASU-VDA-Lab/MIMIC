module fake_netlist_5_1985_n_1817 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1817);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1817;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1752;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_9),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_94),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_48),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_15),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_130),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_48),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_67),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_35),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_12),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_65),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_68),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_32),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_0),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_42),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_159),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_7),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_39),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_95),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_29),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_150),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_24),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_104),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_14),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_33),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_11),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_1),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_134),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_127),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_93),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_42),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_133),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_55),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_45),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_63),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_4),
.Y(n_207)
);

INVxp33_ASAP7_75t_SL g208 ( 
.A(n_96),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_24),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_12),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_29),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_142),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_88),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_23),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_129),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_2),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_70),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_19),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_126),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_92),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_118),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_9),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_163),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_10),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_112),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_145),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_98),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_56),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_83),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_2),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_61),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_122),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_40),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_101),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_38),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_138),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_105),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_151),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_135),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_74),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_4),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_27),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_34),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_110),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_44),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_27),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_30),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_141),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_58),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_44),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_56),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_140),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_35),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_152),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_111),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_40),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_49),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_161),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_6),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_156),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_148),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_37),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_28),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_51),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_37),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_117),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_11),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_66),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_124),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_69),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_23),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_75),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_116),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_85),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_41),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_5),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_34),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_16),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_107),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_72),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_36),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_115),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_160),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_50),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_59),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_49),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_125),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_19),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_144),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_102),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_32),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_139),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_28),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_43),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_6),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_7),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_18),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_71),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_79),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_22),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_155),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_26),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_97),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_132),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_106),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_123),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_80),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_22),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_136),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_73),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_131),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_120),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_50),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_162),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_14),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_91),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_17),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_109),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_20),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_119),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_8),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_45),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_62),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_21),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_31),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_17),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_165),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_208),
.B(n_0),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_167),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_292),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_239),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_289),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_172),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_292),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_177),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_292),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_292),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_180),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_181),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_216),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_187),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_192),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_194),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_200),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_216),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_216),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_216),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_201),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_203),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_258),
.B(n_1),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_216),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_213),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_215),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_219),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_246),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_221),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_223),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_225),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_226),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_227),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_229),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_231),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_179),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_179),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_246),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_258),
.B(n_3),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_232),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_246),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_234),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_236),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_248),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_246),
.Y(n_377)
);

INVxp33_ASAP7_75t_SL g378 ( 
.A(n_309),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_238),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_252),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_246),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_188),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_260),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_261),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_266),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_269),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_188),
.Y(n_387)
);

INVxp33_ASAP7_75t_SL g388 ( 
.A(n_309),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_233),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_233),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_217),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_270),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_173),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_272),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_235),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_235),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_274),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_280),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_242),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_282),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_242),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_314),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_285),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_238),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_314),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_299),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_391),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_345),
.B(n_300),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g409 ( 
.A(n_328),
.B(n_184),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_345),
.B(n_302),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_328),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_350),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_350),
.B(n_231),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_351),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_391),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_351),
.B(n_304),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_331),
.B(n_238),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_335),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_356),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_393),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_360),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_338),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_360),
.Y(n_432)
);

AND2x2_ASAP7_75t_SL g433 ( 
.A(n_355),
.B(n_184),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_340),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_370),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_340),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_341),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_370),
.B(n_169),
.Y(n_439)
);

AND3x1_ASAP7_75t_L g440 ( 
.A(n_369),
.B(n_290),
.C(n_170),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_371),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_373),
.B(n_169),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_373),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_343),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_377),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_377),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_381),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_381),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_343),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_387),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_368),
.B(n_175),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_387),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_389),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_389),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_378),
.B(n_168),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_390),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_390),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_395),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_395),
.B(n_396),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_L g462 ( 
.A(n_396),
.B(n_290),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_399),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_399),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_401),
.B(n_174),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_401),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_402),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_402),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_405),
.B(n_174),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_405),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_330),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_332),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_337),
.B(n_305),
.Y(n_473)
);

BUFx8_ASAP7_75t_L g474 ( 
.A(n_379),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_342),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_344),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_346),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_347),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_348),
.Y(n_479)
);

OAI22xp33_ASAP7_75t_L g480 ( 
.A1(n_441),
.A2(n_404),
.B1(n_388),
.B2(n_247),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_427),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_411),
.Y(n_482)
);

NAND2xp33_ASAP7_75t_L g483 ( 
.A(n_420),
.B(n_349),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_416),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_R g485 ( 
.A(n_457),
.B(n_353),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_422),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_441),
.B(n_354),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_416),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_418),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_465),
.B(n_357),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_416),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_406),
.B(n_359),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_418),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_R g494 ( 
.A(n_457),
.B(n_362),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_406),
.B(n_363),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_433),
.B(n_365),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_418),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_471),
.B(n_375),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_L g500 ( 
.A(n_420),
.B(n_383),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_422),
.Y(n_501)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_427),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_471),
.B(n_190),
.Y(n_503)
);

OAI22xp33_ASAP7_75t_L g504 ( 
.A1(n_453),
.A2(n_241),
.B1(n_193),
.B2(n_326),
.Y(n_504)
);

NAND3xp33_ASAP7_75t_L g505 ( 
.A(n_433),
.B(n_183),
.C(n_176),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_433),
.B(n_384),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_433),
.B(n_385),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_409),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_473),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_474),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_411),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_477),
.B(n_386),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_418),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_409),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

AO22x2_ASAP7_75t_L g516 ( 
.A1(n_477),
.A2(n_224),
.B1(n_327),
.B2(n_170),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_453),
.A2(n_414),
.B1(n_442),
.B2(n_439),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_414),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_407),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_407),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_429),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_440),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_411),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_471),
.B(n_392),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_416),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_416),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_429),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_408),
.B(n_410),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_429),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_416),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_412),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_412),
.Y(n_534)
);

AND2x6_ASAP7_75t_L g535 ( 
.A(n_471),
.B(n_190),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_471),
.B(n_394),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_471),
.B(n_398),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_474),
.B(n_339),
.Y(n_538)
);

AND2x2_ASAP7_75t_SL g539 ( 
.A(n_440),
.B(n_199),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_429),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_436),
.Y(n_541)
);

AND2x2_ASAP7_75t_SL g542 ( 
.A(n_471),
.B(n_199),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_436),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_477),
.B(n_358),
.Y(n_544)
);

NOR2x1p5_ASAP7_75t_L g545 ( 
.A(n_478),
.B(n_166),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_408),
.B(n_410),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_471),
.B(n_361),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_422),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_412),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_412),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_479),
.B(n_364),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_465),
.B(n_176),
.Y(n_552)
);

INVx5_ASAP7_75t_L g553 ( 
.A(n_409),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_416),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_479),
.B(n_473),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_479),
.B(n_366),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_414),
.A2(n_230),
.B1(n_327),
.B2(n_224),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_475),
.B(n_372),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_465),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_416),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_417),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_436),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_469),
.B(n_439),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_436),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_414),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_407),
.Y(n_566)
);

BUFx10_ASAP7_75t_L g567 ( 
.A(n_471),
.Y(n_567)
);

NOR2x1p5_ASAP7_75t_L g568 ( 
.A(n_478),
.B(n_475),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_416),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_409),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_422),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_469),
.B(n_439),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_414),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_419),
.B(n_475),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_436),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_417),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_407),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_475),
.B(n_403),
.Y(n_578)
);

AND2x2_ASAP7_75t_SL g579 ( 
.A(n_476),
.B(n_254),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_417),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_417),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_419),
.B(n_220),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_449),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_422),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_474),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_469),
.B(n_183),
.Y(n_586)
);

NAND3xp33_ASAP7_75t_L g587 ( 
.A(n_442),
.B(n_237),
.C(n_212),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_476),
.B(n_374),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_422),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_449),
.Y(n_590)
);

AND2x4_ASAP7_75t_SL g591 ( 
.A(n_476),
.B(n_376),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_449),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_476),
.B(n_380),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_449),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_442),
.B(n_212),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_478),
.B(n_397),
.Y(n_596)
);

AND2x6_ASAP7_75t_L g597 ( 
.A(n_478),
.B(n_254),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_472),
.B(n_400),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_445),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_462),
.A2(n_214),
.B1(n_320),
.B2(n_323),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_445),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_414),
.A2(n_478),
.B1(n_409),
.B2(n_262),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_409),
.A2(n_209),
.B1(n_249),
.B2(n_230),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_422),
.Y(n_604)
);

CKINVDCx6p67_ASAP7_75t_R g605 ( 
.A(n_474),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_445),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_422),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_451),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_472),
.B(n_306),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_461),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_422),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_415),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_413),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_413),
.Y(n_614)
);

AND2x6_ASAP7_75t_L g615 ( 
.A(n_423),
.B(n_279),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_425),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_415),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_474),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_415),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_421),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_421),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_461),
.B(n_237),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_451),
.Y(n_623)
);

AO21x2_ASAP7_75t_L g624 ( 
.A1(n_462),
.A2(n_255),
.B(n_206),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_423),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_466),
.B(n_240),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_425),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_421),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_452),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_426),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_518),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_623),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_518),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_510),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_518),
.Y(n_635)
);

AND2x6_ASAP7_75t_L g636 ( 
.A(n_574),
.B(n_530),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_555),
.B(n_423),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_509),
.B(n_293),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_573),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_542),
.B(n_423),
.Y(n_640)
);

NOR3xp33_ASAP7_75t_L g641 ( 
.A(n_480),
.B(n_182),
.C(n_178),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_487),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_610),
.B(n_185),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_546),
.B(n_423),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_487),
.B(n_186),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_496),
.B(n_189),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_481),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_506),
.B(n_197),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_579),
.B(n_423),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_L g650 ( 
.A(n_568),
.B(n_217),
.Y(n_650)
);

A2O1A1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_505),
.A2(n_171),
.B(n_295),
.C(n_278),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_579),
.B(n_563),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_507),
.A2(n_505),
.B1(n_517),
.B2(n_579),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_559),
.A2(n_171),
.B(n_295),
.C(n_278),
.Y(n_654)
);

A2O1A1Ixp33_ASAP7_75t_L g655 ( 
.A1(n_563),
.A2(n_279),
.B(n_324),
.C(n_315),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_572),
.B(n_582),
.Y(n_656)
);

NOR2xp67_ASAP7_75t_L g657 ( 
.A(n_544),
.B(n_452),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_573),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_512),
.B(n_492),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_573),
.Y(n_660)
);

A2O1A1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_572),
.A2(n_301),
.B(n_303),
.C(n_298),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_490),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_519),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_608),
.B(n_423),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_608),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_520),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_L g667 ( 
.A1(n_600),
.A2(n_301),
.B1(n_303),
.B2(n_298),
.Y(n_667)
);

BUFx5_ASAP7_75t_L g668 ( 
.A(n_567),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_629),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_629),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_495),
.B(n_542),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_520),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_490),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_520),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_542),
.B(n_423),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_SL g676 ( 
.A(n_605),
.B(n_474),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_519),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_599),
.B(n_423),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_613),
.Y(n_679)
);

NAND2x1_ASAP7_75t_L g680 ( 
.A(n_565),
.B(n_424),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_565),
.B(n_430),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_L g682 ( 
.A(n_568),
.B(n_217),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_521),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_599),
.B(n_430),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_567),
.B(n_430),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_613),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_601),
.B(n_430),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_601),
.B(n_430),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_606),
.B(n_430),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_545),
.A2(n_336),
.B1(n_334),
.B2(n_317),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_521),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_545),
.A2(n_310),
.B1(n_319),
.B2(n_321),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_606),
.B(n_430),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_614),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_614),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_502),
.B(n_466),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_567),
.B(n_430),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_493),
.B(n_430),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_602),
.A2(n_244),
.B1(n_240),
.B2(n_291),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_552),
.B(n_431),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_552),
.B(n_431),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_521),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_551),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_566),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_616),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_516),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_591),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_591),
.B(n_466),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_586),
.B(n_431),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_616),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_586),
.B(n_431),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_595),
.B(n_431),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_595),
.B(n_431),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_567),
.B(n_431),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_489),
.B(n_431),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_627),
.B(n_431),
.Y(n_716)
);

BUFx6f_ASAP7_75t_SL g717 ( 
.A(n_539),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_523),
.B(n_198),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_627),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_622),
.A2(n_166),
.B(n_191),
.C(n_195),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_504),
.B(n_204),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_626),
.B(n_244),
.Y(n_722)
);

AND2x2_ASAP7_75t_SL g723 ( 
.A(n_539),
.B(n_483),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_630),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_591),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_630),
.B(n_434),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_489),
.B(n_434),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_497),
.B(n_513),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_497),
.B(n_434),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_578),
.B(n_207),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_513),
.B(n_434),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_515),
.B(n_434),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_612),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_515),
.B(n_434),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_571),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_612),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_499),
.A2(n_268),
.B1(n_313),
.B2(n_315),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_485),
.Y(n_738)
);

BUFx8_ASAP7_75t_L g739 ( 
.A(n_585),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_617),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_522),
.B(n_434),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_525),
.A2(n_268),
.B1(n_313),
.B2(n_291),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_522),
.B(n_434),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_566),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_617),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_609),
.B(n_536),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_619),
.Y(n_747)
);

NOR2xp67_ASAP7_75t_L g748 ( 
.A(n_556),
.B(n_455),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_537),
.B(n_210),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_600),
.B(n_211),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_619),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_527),
.B(n_529),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_539),
.B(n_218),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_571),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_500),
.A2(n_312),
.B1(n_311),
.B2(n_308),
.Y(n_755)
);

NAND3xp33_ASAP7_75t_L g756 ( 
.A(n_494),
.B(n_593),
.C(n_558),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_566),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_527),
.B(n_434),
.Y(n_758)
);

AND2x4_ASAP7_75t_SL g759 ( 
.A(n_605),
.B(n_273),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_529),
.B(n_437),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_531),
.B(n_437),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_531),
.B(n_540),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_SL g763 ( 
.A1(n_598),
.A2(n_243),
.B1(n_222),
.B2(n_228),
.Y(n_763)
);

INVxp33_ASAP7_75t_L g764 ( 
.A(n_588),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_516),
.A2(n_191),
.B1(n_264),
.B2(n_195),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_SL g766 ( 
.A1(n_538),
.A2(n_273),
.B1(n_283),
.B2(n_287),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_516),
.A2(n_249),
.B1(n_202),
.B2(n_209),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_620),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_540),
.B(n_437),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_541),
.B(n_437),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_541),
.B(n_437),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_543),
.B(n_437),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_543),
.B(n_245),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_577),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_547),
.A2(n_597),
.B1(n_596),
.B2(n_622),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_562),
.B(n_437),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_516),
.A2(n_250),
.B1(n_202),
.B2(n_262),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_562),
.B(n_437),
.Y(n_778)
);

CKINVDCx11_ASAP7_75t_R g779 ( 
.A(n_585),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_577),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_626),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_564),
.B(n_575),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_564),
.B(n_437),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_580),
.Y(n_784)
);

AND2x6_ASAP7_75t_SL g785 ( 
.A(n_622),
.B(n_196),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_575),
.B(n_438),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_622),
.B(n_618),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_620),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_589),
.B(n_438),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_SL g790 ( 
.A(n_557),
.B(n_251),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_622),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_587),
.B(n_253),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_484),
.B(n_438),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_597),
.A2(n_307),
.B1(n_287),
.B2(n_283),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_621),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_484),
.B(n_438),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_484),
.B(n_438),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_621),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_580),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_484),
.B(n_438),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_488),
.B(n_438),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_659),
.B(n_597),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_668),
.B(n_488),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_644),
.A2(n_501),
.B(n_486),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_659),
.A2(n_587),
.B(n_196),
.C(n_250),
.Y(n_805)
);

CKINVDCx10_ASAP7_75t_R g806 ( 
.A(n_717),
.Y(n_806)
);

NOR2x2_ASAP7_75t_L g807 ( 
.A(n_667),
.B(n_628),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_636),
.B(n_597),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_685),
.A2(n_501),
.B(n_486),
.Y(n_809)
);

O2A1O1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_652),
.A2(n_628),
.B(n_581),
.C(n_583),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_671),
.A2(n_603),
.B1(n_324),
.B2(n_607),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_685),
.A2(n_501),
.B(n_486),
.Y(n_812)
);

OAI21xp33_ASAP7_75t_L g813 ( 
.A1(n_638),
.A2(n_257),
.B(n_256),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_697),
.A2(n_501),
.B(n_486),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_697),
.A2(n_548),
.B(n_604),
.Y(n_815)
);

NOR3xp33_ASAP7_75t_L g816 ( 
.A(n_756),
.B(n_259),
.C(n_205),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_754),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_750),
.A2(n_264),
.B(n_297),
.C(n_455),
.Y(n_818)
);

AO21x1_ASAP7_75t_L g819 ( 
.A1(n_653),
.A2(n_583),
.B(n_581),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_636),
.B(n_597),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_714),
.A2(n_548),
.B(n_625),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_668),
.B(n_663),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_658),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_733),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_663),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_714),
.A2(n_548),
.B(n_625),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_636),
.B(n_597),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_679),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_696),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_649),
.A2(n_548),
.B(n_625),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_637),
.A2(n_607),
.B(n_604),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_638),
.B(n_624),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_725),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_789),
.A2(n_607),
.B(n_604),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_636),
.B(n_597),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_706),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_686),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_636),
.B(n_488),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_736),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_675),
.A2(n_571),
.B(n_491),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_700),
.A2(n_709),
.B(n_701),
.Y(n_841)
);

CKINVDCx10_ASAP7_75t_R g842 ( 
.A(n_717),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_711),
.A2(n_571),
.B(n_491),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_712),
.A2(n_571),
.B(n_491),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_713),
.A2(n_491),
.B(n_526),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_656),
.B(n_488),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_651),
.A2(n_706),
.B(n_661),
.C(n_654),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_781),
.B(n_526),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_651),
.A2(n_594),
.B(n_580),
.C(n_524),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_646),
.B(n_526),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_646),
.B(n_526),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_750),
.A2(n_297),
.B(n_455),
.C(n_594),
.Y(n_852)
);

AO21x1_ASAP7_75t_L g853 ( 
.A1(n_753),
.A2(n_511),
.B(n_482),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_648),
.B(n_528),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_707),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_640),
.A2(n_554),
.B(n_528),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_640),
.A2(n_554),
.B(n_528),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_632),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_681),
.A2(n_554),
.B(n_528),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_681),
.A2(n_554),
.B(n_532),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_698),
.A2(n_762),
.B(n_752),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_775),
.A2(n_723),
.B1(n_677),
.B2(n_746),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_648),
.B(n_532),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_677),
.A2(n_663),
.B(n_650),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_723),
.A2(n_560),
.B1(n_532),
.B2(n_569),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_668),
.B(n_532),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_752),
.A2(n_550),
.B(n_498),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_658),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_668),
.B(n_560),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_643),
.B(n_624),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_661),
.A2(n_533),
.B(n_482),
.C(n_592),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_703),
.B(n_584),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_708),
.B(n_624),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_643),
.B(n_263),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_748),
.B(n_560),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_663),
.A2(n_560),
.B(n_569),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_682),
.A2(n_569),
.B(n_611),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_746),
.A2(n_503),
.B1(n_535),
.B2(n_569),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_735),
.A2(n_584),
.B(n_611),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_665),
.B(n_669),
.Y(n_880)
);

OAI21xp33_ASAP7_75t_L g881 ( 
.A1(n_721),
.A2(n_276),
.B(n_267),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_670),
.B(n_694),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_738),
.Y(n_883)
);

AOI21x1_ASAP7_75t_L g884 ( 
.A1(n_762),
.A2(n_511),
.B(n_498),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_754),
.Y(n_885)
);

AOI21xp33_ASAP7_75t_L g886 ( 
.A1(n_645),
.A2(n_275),
.B(n_271),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_728),
.A2(n_561),
.B(n_534),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_791),
.A2(n_584),
.B1(n_611),
.B2(n_592),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_695),
.B(n_584),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_705),
.Y(n_890)
);

BUFx12f_ASAP7_75t_L g891 ( 
.A(n_779),
.Y(n_891)
);

AO21x1_ASAP7_75t_L g892 ( 
.A1(n_753),
.A2(n_742),
.B(n_737),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_654),
.A2(n_550),
.B(n_533),
.C(n_590),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_782),
.A2(n_549),
.B(n_590),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_SL g895 ( 
.A(n_676),
.B(n_265),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_754),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_662),
.B(n_611),
.Y(n_897)
);

BUFx4f_ASAP7_75t_L g898 ( 
.A(n_787),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_668),
.B(n_524),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_754),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_642),
.B(n_534),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_710),
.B(n_719),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_667),
.A2(n_655),
.B(n_699),
.C(n_720),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_764),
.B(n_549),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_668),
.B(n_561),
.Y(n_905)
);

AOI33xp33_ASAP7_75t_L g906 ( 
.A1(n_765),
.A2(n_432),
.A3(n_426),
.B1(n_428),
.B2(n_468),
.B3(n_454),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_735),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_724),
.B(n_576),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_639),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_657),
.B(n_576),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_L g911 ( 
.A(n_660),
.B(n_503),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_793),
.A2(n_514),
.B(n_570),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_673),
.B(n_716),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_645),
.B(n_277),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_740),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_722),
.B(n_503),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_792),
.A2(n_428),
.B(n_432),
.C(n_424),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_722),
.B(n_773),
.Y(n_918)
);

AND2x4_ASAP7_75t_SL g919 ( 
.A(n_634),
.B(n_455),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_792),
.A2(n_455),
.B(n_294),
.C(n_281),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_726),
.B(n_508),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_745),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_796),
.A2(n_570),
.B(n_553),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_749),
.B(n_508),
.Y(n_924)
);

NOR2x1_ASAP7_75t_L g925 ( 
.A(n_730),
.B(n_424),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_678),
.A2(n_503),
.B(n_535),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_773),
.B(n_503),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_721),
.A2(n_286),
.B(n_284),
.C(n_325),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_797),
.A2(n_508),
.B(n_570),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_800),
.A2(n_508),
.B(n_570),
.Y(n_930)
);

AO21x1_ASAP7_75t_L g931 ( 
.A1(n_749),
.A2(n_443),
.B(n_446),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_747),
.B(n_503),
.Y(n_932)
);

BUFx2_ASAP7_75t_SL g933 ( 
.A(n_690),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_680),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_684),
.A2(n_503),
.B(n_535),
.Y(n_935)
);

NAND3xp33_ASAP7_75t_SL g936 ( 
.A(n_641),
.B(n_766),
.C(n_718),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_801),
.A2(n_508),
.B(n_570),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_664),
.A2(n_508),
.B(n_570),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_751),
.B(n_535),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_718),
.B(n_288),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_768),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_763),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_788),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_765),
.A2(n_318),
.B1(n_296),
.B2(n_322),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_647),
.B(n_790),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_687),
.A2(n_689),
.B(n_688),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_693),
.A2(n_514),
.B(n_553),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_767),
.A2(n_777),
.B1(n_794),
.B2(n_795),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_798),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_767),
.A2(n_316),
.B(n_456),
.C(n_454),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_727),
.A2(n_514),
.B(n_553),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_777),
.A2(n_535),
.B1(n_615),
.B2(n_217),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_631),
.B(n_633),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_784),
.B(n_799),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_729),
.A2(n_514),
.B(n_553),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_692),
.A2(n_443),
.B1(n_446),
.B2(n_447),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_785),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_731),
.A2(n_786),
.B(n_741),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_739),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_715),
.A2(n_772),
.B(n_783),
.C(n_734),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_732),
.A2(n_758),
.B(n_760),
.Y(n_961)
);

OAI21xp33_ASAP7_75t_L g962 ( 
.A1(n_755),
.A2(n_435),
.B(n_448),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_635),
.Y(n_963)
);

BUFx2_ASAP7_75t_SL g964 ( 
.A(n_666),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_715),
.A2(n_443),
.B(n_446),
.C(n_447),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_672),
.Y(n_966)
);

AOI21x1_ASAP7_75t_L g967 ( 
.A1(n_734),
.A2(n_435),
.B(n_447),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_674),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_683),
.B(n_535),
.Y(n_969)
);

BUFx4f_ASAP7_75t_L g970 ( 
.A(n_759),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_769),
.A2(n_535),
.B(n_615),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_743),
.A2(n_448),
.B(n_435),
.C(n_468),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_691),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_739),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_702),
.Y(n_975)
);

NOR2x1_ASAP7_75t_L g976 ( 
.A(n_743),
.B(n_448),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_770),
.A2(n_468),
.B(n_463),
.C(n_470),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_704),
.B(n_514),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_744),
.A2(n_615),
.B1(n_409),
.B2(n_438),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_757),
.B(n_438),
.Y(n_980)
);

AO21x1_ASAP7_75t_L g981 ( 
.A1(n_761),
.A2(n_771),
.B(n_783),
.Y(n_981)
);

AOI21x1_ASAP7_75t_L g982 ( 
.A1(n_761),
.A2(n_464),
.B(n_456),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_776),
.A2(n_553),
.B(n_514),
.Y(n_983)
);

CKINVDCx8_ASAP7_75t_R g984 ( 
.A(n_771),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_772),
.A2(n_553),
.B(n_444),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_778),
.A2(n_615),
.B(n_409),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_774),
.Y(n_987)
);

NOR2x1_ASAP7_75t_L g988 ( 
.A(n_778),
.B(n_454),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_780),
.B(n_454),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_649),
.A2(n_615),
.B(n_409),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_644),
.A2(n_444),
.B(n_470),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_659),
.A2(n_615),
.B1(n_409),
.B2(n_444),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_781),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_832),
.B(n_409),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_862),
.A2(n_463),
.B1(n_470),
.B2(n_468),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_918),
.A2(n_459),
.B1(n_470),
.B2(n_467),
.Y(n_996)
);

NOR3xp33_ASAP7_75t_SL g997 ( 
.A(n_883),
.B(n_936),
.C(n_928),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_864),
.A2(n_841),
.B(n_802),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_817),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_858),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_886),
.B(n_456),
.C(n_459),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_825),
.B(n_444),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_825),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_914),
.B(n_8),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_822),
.A2(n_444),
.B(n_467),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_903),
.A2(n_459),
.B(n_467),
.C(n_464),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_SL g1007 ( 
.A(n_942),
.B(n_456),
.C(n_459),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_963),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_828),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_870),
.B(n_444),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_836),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_872),
.B(n_444),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_861),
.A2(n_615),
.B(n_467),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_SL g1014 ( 
.A1(n_816),
.A2(n_464),
.B(n_463),
.C(n_217),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_833),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_822),
.A2(n_444),
.B(n_463),
.Y(n_1016)
);

INVx5_ASAP7_75t_L g1017 ( 
.A(n_817),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_829),
.B(n_464),
.Y(n_1018)
);

AO21x1_ASAP7_75t_L g1019 ( 
.A1(n_850),
.A2(n_217),
.B(n_13),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_993),
.B(n_10),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_940),
.B(n_460),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_873),
.A2(n_444),
.B1(n_458),
.B2(n_450),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_875),
.A2(n_460),
.B(n_458),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_966),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_933),
.A2(n_217),
.B1(n_458),
.B2(n_450),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_824),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_873),
.A2(n_460),
.B1(n_458),
.B2(n_450),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_993),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_839),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_823),
.A2(n_460),
.B1(n_458),
.B2(n_450),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_922),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_941),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_898),
.B(n_217),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_SL g1034 ( 
.A(n_974),
.B(n_460),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_817),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_891),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_907),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_928),
.A2(n_13),
.B(n_15),
.C(n_16),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_R g1039 ( 
.A(n_806),
.B(n_64),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_874),
.B(n_18),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_851),
.A2(n_460),
.B(n_458),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_884),
.A2(n_76),
.B(n_158),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_854),
.A2(n_460),
.B(n_458),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_837),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_898),
.B(n_460),
.Y(n_1045)
);

NAND3xp33_ASAP7_75t_L g1046 ( 
.A(n_881),
.B(n_460),
.C(n_458),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_817),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_863),
.A2(n_846),
.B(n_924),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_872),
.B(n_458),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_SL g1050 ( 
.A1(n_920),
.A2(n_852),
.B(n_950),
.C(n_818),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_813),
.B(n_20),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_836),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_945),
.B(n_450),
.Y(n_1053)
);

CKINVDCx8_ASAP7_75t_R g1054 ( 
.A(n_842),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_904),
.B(n_450),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_919),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_885),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_920),
.A2(n_21),
.B(n_25),
.C(n_26),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_904),
.B(n_450),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_890),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_847),
.A2(n_450),
.B(n_30),
.C(n_31),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_805),
.A2(n_25),
.B(n_33),
.C(n_36),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_949),
.Y(n_1063)
);

CKINVDCx6p67_ASAP7_75t_R g1064 ( 
.A(n_959),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_902),
.B(n_450),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_960),
.A2(n_38),
.B(n_39),
.C(n_41),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_833),
.B(n_43),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_SL g1068 ( 
.A1(n_816),
.A2(n_84),
.B(n_137),
.C(n_128),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_949),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_901),
.B(n_81),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_901),
.B(n_82),
.Y(n_1071)
);

CKINVDCx11_ASAP7_75t_R g1072 ( 
.A(n_957),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_882),
.A2(n_46),
.B(n_47),
.C(n_51),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_SL g1074 ( 
.A(n_944),
.B(n_46),
.C(n_47),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_880),
.B(n_52),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_915),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_913),
.B(n_87),
.Y(n_1077)
);

O2A1O1Ixp5_ASAP7_75t_L g1078 ( 
.A1(n_931),
.A2(n_86),
.B(n_114),
.C(n_113),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_805),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_927),
.A2(n_78),
.B(n_108),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_855),
.B(n_53),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_924),
.A2(n_89),
.B(n_103),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_823),
.B(n_77),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_925),
.A2(n_54),
.B(n_55),
.C(n_57),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_943),
.Y(n_1085)
);

OR2x6_ASAP7_75t_L g1086 ( 
.A(n_855),
.B(n_60),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_984),
.B(n_57),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_913),
.B(n_90),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_897),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_804),
.A2(n_99),
.B(n_100),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_868),
.A2(n_58),
.B1(n_143),
.B2(n_948),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_803),
.A2(n_869),
.B(n_866),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_909),
.Y(n_1093)
);

O2A1O1Ixp5_ASAP7_75t_L g1094 ( 
.A1(n_892),
.A2(n_853),
.B(n_819),
.C(n_888),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_908),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_856),
.A2(n_857),
.B(n_840),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_897),
.A2(n_895),
.B1(n_916),
.B2(n_909),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_803),
.A2(n_869),
.B(n_866),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_906),
.B(n_950),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_885),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_906),
.B(n_848),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_852),
.A2(n_818),
.B(n_810),
.C(n_917),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_807),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_899),
.A2(n_905),
.B(n_830),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_970),
.B(n_868),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_970),
.B(n_910),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_907),
.B(n_885),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_878),
.A2(n_962),
.B(n_871),
.C(n_990),
.Y(n_1108)
);

INVx4_ASAP7_75t_L g1109 ( 
.A(n_885),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_958),
.A2(n_961),
.B(n_808),
.C(n_835),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_820),
.A2(n_827),
.B(n_893),
.C(n_849),
.Y(n_1111)
);

NAND2x1p5_ASAP7_75t_L g1112 ( 
.A(n_900),
.B(n_896),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_889),
.A2(n_865),
.B1(n_838),
.B2(n_964),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_956),
.A2(n_977),
.B(n_811),
.C(n_968),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_973),
.B(n_975),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_987),
.A2(n_981),
.B1(n_952),
.B2(n_976),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_989),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_954),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_900),
.B(n_896),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_988),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_934),
.B(n_992),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_899),
.A2(n_905),
.B(n_812),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_934),
.A2(n_877),
.B1(n_814),
.B2(n_809),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_953),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_921),
.B(n_953),
.Y(n_1125)
);

INVxp67_ASAP7_75t_L g1126 ( 
.A(n_978),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_946),
.A2(n_844),
.B(n_843),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_SL g1128 ( 
.A1(n_926),
.A2(n_935),
.B(n_971),
.C(n_911),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_921),
.A2(n_978),
.B1(n_939),
.B2(n_932),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_952),
.A2(n_815),
.B1(n_821),
.B2(n_826),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_876),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_980),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_845),
.A2(n_831),
.B(n_834),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_967),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_859),
.A2(n_860),
.B(n_991),
.C(n_969),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_979),
.A2(n_986),
.B1(n_867),
.B2(n_985),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_887),
.B(n_894),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_982),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_977),
.B(n_879),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_965),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_951),
.B(n_983),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_972),
.A2(n_947),
.B(n_955),
.C(n_938),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_912),
.A2(n_923),
.B1(n_929),
.B2(n_930),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_937),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_864),
.A2(n_668),
.B(n_685),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_864),
.A2(n_668),
.B(n_685),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_862),
.A2(n_659),
.B1(n_756),
.B2(n_918),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_832),
.B(n_636),
.Y(n_1148)
);

AOI21x1_ASAP7_75t_L g1149 ( 
.A1(n_924),
.A2(n_822),
.B(n_899),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_829),
.B(n_509),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_1054),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_998),
.A2(n_1048),
.B(n_1123),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1127),
.A2(n_1110),
.B(n_1137),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1133),
.A2(n_1096),
.B(n_1145),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1137),
.A2(n_1108),
.B(n_1146),
.Y(n_1155)
);

CKINVDCx16_ASAP7_75t_R g1156 ( 
.A(n_1036),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_1015),
.Y(n_1157)
);

NOR2xp67_ASAP7_75t_L g1158 ( 
.A(n_1106),
.B(n_1105),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1130),
.A2(n_1121),
.B(n_1128),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_1148),
.A2(n_1102),
.B(n_1141),
.Y(n_1160)
);

OAI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_1040),
.A2(n_1004),
.B(n_1051),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1122),
.A2(n_1104),
.B(n_1149),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_L g1163 ( 
.A(n_997),
.B(n_1074),
.C(n_1087),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1150),
.B(n_1028),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1147),
.A2(n_1075),
.B(n_1071),
.C(n_1070),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1044),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1103),
.B(n_1052),
.Y(n_1167)
);

BUFx12f_ASAP7_75t_L g1168 ( 
.A(n_1072),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1064),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1124),
.Y(n_1170)
);

AO21x2_ASAP7_75t_L g1171 ( 
.A1(n_1148),
.A2(n_1139),
.B(n_1013),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_1019),
.A2(n_1111),
.A3(n_1143),
.B(n_1113),
.Y(n_1172)
);

INVx3_ASAP7_75t_SL g1173 ( 
.A(n_1056),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1010),
.A2(n_1135),
.B(n_1021),
.Y(n_1174)
);

O2A1O1Ixp5_ASAP7_75t_L g1175 ( 
.A1(n_1094),
.A2(n_1078),
.B(n_1071),
.C(n_1070),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_995),
.A2(n_1139),
.A3(n_1061),
.B(n_1006),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1066),
.A2(n_1084),
.B(n_1038),
.C(n_1073),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1010),
.A2(n_1142),
.B(n_1114),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1117),
.A2(n_1095),
.B1(n_1116),
.B2(n_1097),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1099),
.A2(n_1049),
.A3(n_1091),
.B(n_1012),
.Y(n_1180)
);

AND2x2_ASAP7_75t_SL g1181 ( 
.A(n_1034),
.B(n_1081),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1060),
.Y(n_1182)
);

O2A1O1Ixp5_ASAP7_75t_L g1183 ( 
.A1(n_1053),
.A2(n_1131),
.B(n_1033),
.C(n_1083),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_1086),
.B(n_1003),
.Y(n_1184)
);

NAND2x1_ASAP7_75t_L g1185 ( 
.A(n_1037),
.B(n_1003),
.Y(n_1185)
);

AOI221x1_ASAP7_75t_L g1186 ( 
.A1(n_1080),
.A2(n_1046),
.B1(n_1090),
.B2(n_1099),
.C(n_1098),
.Y(n_1186)
);

OAI22x1_ASAP7_75t_L g1187 ( 
.A1(n_1020),
.A2(n_1069),
.B1(n_1063),
.B2(n_1076),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_994),
.A2(n_1125),
.B(n_1092),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1089),
.A2(n_1086),
.B1(n_1118),
.B2(n_1029),
.Y(n_1189)
);

BUFx8_ASAP7_75t_L g1190 ( 
.A(n_1067),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1037),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1049),
.A2(n_1012),
.A3(n_1043),
.B(n_1144),
.Y(n_1192)
);

BUFx2_ASAP7_75t_R g1193 ( 
.A(n_1107),
.Y(n_1193)
);

CKINVDCx11_ASAP7_75t_R g1194 ( 
.A(n_1086),
.Y(n_1194)
);

INVxp67_ASAP7_75t_SL g1195 ( 
.A(n_1011),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1005),
.A2(n_1016),
.B(n_1042),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1043),
.A2(n_1041),
.B(n_1134),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1026),
.B(n_1032),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1132),
.A2(n_994),
.B(n_1050),
.Y(n_1199)
);

AND2x6_ASAP7_75t_L g1200 ( 
.A(n_999),
.B(n_1047),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_996),
.A2(n_1027),
.A3(n_1131),
.B(n_1022),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1039),
.Y(n_1202)
);

OR2x2_ASAP7_75t_L g1203 ( 
.A(n_1031),
.B(n_1085),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1065),
.A2(n_1017),
.B(n_1059),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1101),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1017),
.A2(n_1055),
.B(n_1136),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1115),
.Y(n_1207)
);

O2A1O1Ixp5_ASAP7_75t_L g1208 ( 
.A1(n_1080),
.A2(n_1045),
.B(n_1088),
.C(n_1077),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1093),
.B(n_1126),
.Y(n_1209)
);

NOR4xp25_ASAP7_75t_L g1210 ( 
.A(n_1058),
.B(n_1062),
.C(n_1079),
.D(n_1007),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1134),
.A2(n_1023),
.B(n_1088),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1077),
.A2(n_1101),
.A3(n_1030),
.B(n_1082),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1017),
.A2(n_1140),
.B(n_1115),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1120),
.B(n_1008),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1018),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1024),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1025),
.A2(n_1129),
.B(n_1001),
.C(n_1068),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1035),
.A2(n_1057),
.A3(n_1109),
.B(n_1014),
.Y(n_1218)
);

AO21x2_ASAP7_75t_L g1219 ( 
.A1(n_1119),
.A2(n_1138),
.B(n_1002),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1035),
.B(n_1109),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1057),
.A2(n_1138),
.A3(n_1002),
.B(n_1112),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_999),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1112),
.A2(n_1138),
.B(n_1047),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_999),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1047),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1100),
.Y(n_1226)
);

NAND2x1p5_ASAP7_75t_L g1227 ( 
.A(n_1100),
.B(n_1017),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1100),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1095),
.B(n_659),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_SL g1230 ( 
.A1(n_1061),
.A2(n_1066),
.B(n_920),
.C(n_1099),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1004),
.A2(n_659),
.B(n_1040),
.C(n_756),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1102),
.A2(n_931),
.A3(n_853),
.B(n_819),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1095),
.B(n_659),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1015),
.B(n_833),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_999),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1102),
.A2(n_931),
.A3(n_853),
.B(n_819),
.Y(n_1236)
);

AO32x2_ASAP7_75t_L g1237 ( 
.A1(n_1147),
.A2(n_862),
.A3(n_1091),
.B1(n_653),
.B2(n_995),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1103),
.B(n_703),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1095),
.B(n_659),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1004),
.A2(n_703),
.B(n_659),
.C(n_420),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1102),
.A2(n_931),
.A3(n_853),
.B(n_819),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1102),
.A2(n_931),
.A3(n_853),
.B(n_819),
.Y(n_1243)
);

INVx6_ASAP7_75t_L g1244 ( 
.A(n_1000),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1127),
.A2(n_1133),
.B(n_1096),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_1028),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1127),
.A2(n_1133),
.B(n_1096),
.Y(n_1247)
);

AOI221x1_ASAP7_75t_L g1248 ( 
.A1(n_1147),
.A2(n_1066),
.B1(n_1061),
.B2(n_756),
.C(n_998),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1124),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1252)
);

AOI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1049),
.A2(n_998),
.B(n_1048),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1254)
);

BUFx4_ASAP7_75t_SL g1255 ( 
.A(n_1000),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1009),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1095),
.B(n_659),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1094),
.A2(n_1048),
.B(n_1148),
.Y(n_1261)
);

NAND3xp33_ASAP7_75t_SL g1262 ( 
.A(n_1004),
.B(n_659),
.C(n_703),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1103),
.B(n_703),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1000),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1127),
.A2(n_1133),
.B(n_1096),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1127),
.A2(n_1133),
.B(n_1096),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1095),
.B(n_659),
.Y(n_1270)
);

AO21x1_ASAP7_75t_L g1271 ( 
.A1(n_1147),
.A2(n_659),
.B(n_862),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1147),
.A2(n_659),
.B(n_671),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1147),
.A2(n_659),
.B(n_671),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1095),
.B(n_659),
.Y(n_1274)
);

AO31x2_ASAP7_75t_L g1275 ( 
.A1(n_1102),
.A2(n_931),
.A3(n_853),
.B(n_819),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1103),
.B(n_703),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1004),
.A2(n_659),
.B(n_1040),
.C(n_756),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1096),
.A2(n_931),
.B(n_998),
.Y(n_1279)
);

NAND3x1_ASAP7_75t_L g1280 ( 
.A(n_1087),
.B(n_750),
.C(n_600),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1036),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1103),
.B(n_829),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1094),
.A2(n_1048),
.B(n_1148),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1103),
.B(n_829),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1009),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1095),
.B(n_659),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1004),
.A2(n_703),
.B(n_659),
.C(n_420),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1127),
.A2(n_1133),
.B(n_1096),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_SL g1290 ( 
.A1(n_1061),
.A2(n_1066),
.B(n_920),
.C(n_1099),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1103),
.B(n_703),
.Y(n_1291)
);

AOI221x1_ASAP7_75t_L g1292 ( 
.A1(n_1147),
.A2(n_1066),
.B1(n_1061),
.B2(n_756),
.C(n_998),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1102),
.A2(n_931),
.A3(n_853),
.B(n_819),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1037),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1102),
.A2(n_931),
.A3(n_853),
.B(n_819),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1004),
.A2(n_703),
.B(n_659),
.C(n_420),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1004),
.A2(n_659),
.B(n_1040),
.C(n_756),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1036),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1000),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_998),
.A2(n_668),
.B(n_1048),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1095),
.B(n_659),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1124),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1161),
.A2(n_1262),
.B1(n_1271),
.B2(n_1163),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1229),
.A2(n_1259),
.B1(n_1301),
.B2(n_1286),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1170),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1181),
.A2(n_1280),
.B1(n_1273),
.B2(n_1272),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1282),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1233),
.A2(n_1240),
.B1(n_1270),
.B2(n_1274),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1182),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1231),
.A2(n_1278),
.B1(n_1297),
.B2(n_1238),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1265),
.A2(n_1277),
.B1(n_1291),
.B2(n_1189),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1165),
.A2(n_1241),
.B1(n_1296),
.B2(n_1287),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1244),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1234),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1266),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1191),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1285),
.Y(n_1317)
);

BUFx10_ASAP7_75t_L g1318 ( 
.A(n_1234),
.Y(n_1318)
);

CKINVDCx14_ASAP7_75t_R g1319 ( 
.A(n_1151),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_1156),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1194),
.A2(n_1179),
.B1(n_1207),
.B2(n_1159),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1184),
.A2(n_1158),
.B1(n_1284),
.B2(n_1246),
.Y(n_1322)
);

BUFx12f_ASAP7_75t_L g1323 ( 
.A(n_1281),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1215),
.B(n_1214),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1166),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1200),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1184),
.A2(n_1195),
.B1(n_1193),
.B2(n_1164),
.Y(n_1327)
);

CKINVDCx11_ASAP7_75t_R g1328 ( 
.A(n_1168),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1187),
.A2(n_1155),
.B1(n_1205),
.B2(n_1178),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1294),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1249),
.Y(n_1331)
);

OAI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1248),
.A2(n_1292),
.B1(n_1203),
.B2(n_1257),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1302),
.Y(n_1333)
);

BUFx4f_ASAP7_75t_SL g1334 ( 
.A(n_1173),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1205),
.A2(n_1216),
.B1(n_1209),
.B2(n_1188),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1235),
.Y(n_1336)
);

BUFx10_ASAP7_75t_L g1337 ( 
.A(n_1202),
.Y(n_1337)
);

INVx8_ASAP7_75t_L g1338 ( 
.A(n_1200),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1171),
.A2(n_1198),
.B1(n_1160),
.B2(n_1190),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1171),
.A2(n_1199),
.B1(n_1279),
.B2(n_1174),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1299),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1228),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1157),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1224),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1217),
.A2(n_1177),
.B(n_1186),
.Y(n_1345)
);

BUFx10_ASAP7_75t_L g1346 ( 
.A(n_1298),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1255),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1169),
.A2(n_1294),
.B1(n_1210),
.B2(n_1206),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1279),
.A2(n_1261),
.B1(n_1283),
.B2(n_1153),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1213),
.A2(n_1220),
.B1(n_1204),
.B2(n_1185),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1226),
.B(n_1225),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1237),
.A2(n_1223),
.B1(n_1152),
.B2(n_1154),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1261),
.A2(n_1283),
.B1(n_1237),
.B2(n_1289),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1235),
.Y(n_1354)
);

BUFx2_ASAP7_75t_SL g1355 ( 
.A(n_1200),
.Y(n_1355)
);

AOI21xp33_ASAP7_75t_L g1356 ( 
.A1(n_1175),
.A2(n_1208),
.B(n_1183),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1222),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1237),
.A2(n_1230),
.B1(n_1290),
.B2(n_1268),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1227),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1245),
.A2(n_1247),
.B1(n_1267),
.B2(n_1211),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1172),
.B(n_1212),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1239),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1219),
.A2(n_1251),
.B1(n_1288),
.B2(n_1276),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1162),
.A2(n_1197),
.B1(n_1219),
.B2(n_1300),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1221),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1250),
.A2(n_1263),
.B1(n_1254),
.B2(n_1256),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1221),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1172),
.B(n_1212),
.Y(n_1368)
);

INVx4_ASAP7_75t_L g1369 ( 
.A(n_1218),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1218),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1252),
.A2(n_1269),
.B1(n_1264),
.B2(n_1258),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1172),
.B(n_1212),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1218),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1260),
.Y(n_1374)
);

INVx11_ASAP7_75t_L g1375 ( 
.A(n_1232),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1232),
.Y(n_1376)
);

INVx6_ASAP7_75t_L g1377 ( 
.A(n_1176),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1180),
.B(n_1242),
.Y(n_1378)
);

INVx3_ASAP7_75t_SL g1379 ( 
.A(n_1236),
.Y(n_1379)
);

OAI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1253),
.A2(n_1176),
.B1(n_1180),
.B2(n_1236),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1242),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1196),
.A2(n_1176),
.B1(n_1180),
.B2(n_1243),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1243),
.A2(n_1275),
.B1(n_1293),
.B2(n_1295),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1243),
.Y(n_1384)
);

CKINVDCx11_ASAP7_75t_R g1385 ( 
.A(n_1275),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1293),
.A2(n_1295),
.B1(n_1201),
.B2(n_1192),
.Y(n_1386)
);

INVx6_ASAP7_75t_L g1387 ( 
.A(n_1295),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_1201),
.Y(n_1388)
);

INVx2_ASAP7_75t_R g1389 ( 
.A(n_1201),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1167),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1167),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1182),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1167),
.Y(n_1393)
);

INVx3_ASAP7_75t_SL g1394 ( 
.A(n_1244),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1182),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1161),
.A2(n_1262),
.B1(n_1271),
.B2(n_936),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1167),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1182),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1161),
.A2(n_1262),
.B1(n_1271),
.B2(n_936),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1151),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1161),
.A2(n_1262),
.B1(n_1271),
.B2(n_936),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1181),
.A2(n_756),
.B1(n_538),
.B2(n_659),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1182),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1244),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1280),
.A2(n_1161),
.B1(n_659),
.B2(n_738),
.Y(n_1405)
);

INVx3_ASAP7_75t_SL g1406 ( 
.A(n_1244),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1181),
.A2(n_756),
.B1(n_538),
.B2(n_659),
.Y(n_1407)
);

BUFx12f_ASAP7_75t_L g1408 ( 
.A(n_1281),
.Y(n_1408)
);

CKINVDCx11_ASAP7_75t_R g1409 ( 
.A(n_1168),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1181),
.A2(n_756),
.B1(n_538),
.B2(n_659),
.Y(n_1410)
);

BUFx2_ASAP7_75t_SL g1411 ( 
.A(n_1151),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1182),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1182),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1151),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1167),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1151),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1181),
.A2(n_756),
.B1(n_538),
.B2(n_659),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1161),
.A2(n_1262),
.B1(n_1271),
.B2(n_936),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1181),
.A2(n_756),
.B1(n_538),
.B2(n_659),
.Y(n_1419)
);

BUFx4f_ASAP7_75t_SL g1420 ( 
.A(n_1151),
.Y(n_1420)
);

BUFx8_ASAP7_75t_L g1421 ( 
.A(n_1168),
.Y(n_1421)
);

INVx2_ASAP7_75t_SL g1422 ( 
.A(n_1244),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1244),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1181),
.A2(n_756),
.B1(n_538),
.B2(n_659),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1182),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1280),
.A2(n_1161),
.B1(n_659),
.B2(n_738),
.Y(n_1426)
);

CKINVDCx6p67_ASAP7_75t_R g1427 ( 
.A(n_1281),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1305),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1400),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1378),
.B(n_1361),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1384),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1371),
.A2(n_1364),
.B(n_1366),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1367),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1331),
.Y(n_1434)
);

INVx4_ASAP7_75t_SL g1435 ( 
.A(n_1387),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1414),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1312),
.A2(n_1399),
.B(n_1396),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1333),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1379),
.B(n_1376),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1365),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1364),
.A2(n_1366),
.B(n_1360),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1304),
.B(n_1308),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1338),
.Y(n_1443)
);

AO21x2_ASAP7_75t_L g1444 ( 
.A1(n_1356),
.A2(n_1380),
.B(n_1345),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1379),
.B(n_1383),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1394),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1381),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1318),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1390),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1370),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1388),
.B(n_1385),
.Y(n_1451)
);

AO21x2_ASAP7_75t_L g1452 ( 
.A1(n_1380),
.A2(n_1335),
.B(n_1368),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1375),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_SL g1454 ( 
.A(n_1421),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1393),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1318),
.Y(n_1456)
);

BUFx8_ASAP7_75t_L g1457 ( 
.A(n_1323),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1372),
.Y(n_1458)
);

AOI21xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1310),
.A2(n_1405),
.B(n_1426),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_R g1460 ( 
.A(n_1416),
.B(n_1319),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1360),
.A2(n_1349),
.B(n_1340),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1306),
.A2(n_1321),
.B1(n_1417),
.B2(n_1410),
.Y(n_1462)
);

AO21x2_ASAP7_75t_L g1463 ( 
.A1(n_1335),
.A2(n_1332),
.B(n_1350),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1377),
.Y(n_1464)
);

NAND2x1p5_ASAP7_75t_L g1465 ( 
.A(n_1369),
.B(n_1373),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1386),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1386),
.B(n_1389),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1362),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1332),
.A2(n_1304),
.B(n_1325),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1326),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1389),
.B(n_1339),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1382),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1341),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1329),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1329),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1303),
.B(n_1324),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1339),
.B(n_1374),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1321),
.B(n_1353),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1394),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1309),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1391),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1303),
.B(n_1397),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1415),
.B(n_1401),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1317),
.Y(n_1484)
);

AO21x1_ASAP7_75t_SL g1485 ( 
.A1(n_1401),
.A2(n_1418),
.B(n_1340),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1392),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1395),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1418),
.B(n_1307),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1315),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1398),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1403),
.Y(n_1491)
);

AO21x2_ASAP7_75t_L g1492 ( 
.A1(n_1344),
.A2(n_1363),
.B(n_1425),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1412),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1402),
.B(n_1424),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1413),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1406),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1358),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1407),
.A2(n_1419),
.B(n_1311),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1349),
.A2(n_1353),
.B(n_1316),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1352),
.B(n_1330),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1348),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1355),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1406),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1322),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1338),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1351),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1506),
.B(n_1327),
.Y(n_1507)
);

O2A1O1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1459),
.A2(n_1437),
.B(n_1498),
.C(n_1442),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1438),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1459),
.A2(n_1343),
.B(n_1359),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1506),
.B(n_1342),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1439),
.B(n_1431),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1462),
.A2(n_1411),
.B1(n_1320),
.B2(n_1319),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1494),
.A2(n_1314),
.B(n_1357),
.C(n_1354),
.Y(n_1514)
);

OR2x6_ASAP7_75t_L g1515 ( 
.A(n_1477),
.B(n_1323),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1449),
.B(n_1347),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1451),
.B(n_1500),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1501),
.A2(n_1468),
.B1(n_1504),
.B2(n_1483),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1446),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1444),
.A2(n_1336),
.B(n_1422),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1453),
.B(n_1313),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1444),
.A2(n_1313),
.B(n_1423),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1455),
.B(n_1404),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1446),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1468),
.B(n_1423),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1479),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1428),
.Y(n_1527)
);

AOI211xp5_ASAP7_75t_L g1528 ( 
.A1(n_1501),
.A2(n_1482),
.B(n_1488),
.C(n_1476),
.Y(n_1528)
);

AOI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1474),
.A2(n_1427),
.B1(n_1328),
.B2(n_1334),
.C(n_1421),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1489),
.B(n_1337),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1492),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1481),
.B(n_1420),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1430),
.B(n_1420),
.Y(n_1533)
);

OAI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1432),
.A2(n_1400),
.B(n_1346),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1489),
.B(n_1337),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1473),
.B(n_1346),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1479),
.A2(n_1408),
.B1(n_1328),
.B2(n_1409),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1496),
.A2(n_1408),
.B1(n_1503),
.B2(n_1429),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1435),
.B(n_1464),
.Y(n_1539)
);

OAI211xp5_ASAP7_75t_L g1540 ( 
.A1(n_1474),
.A2(n_1475),
.B(n_1478),
.C(n_1497),
.Y(n_1540)
);

AO21x2_ASAP7_75t_L g1541 ( 
.A1(n_1441),
.A2(n_1463),
.B(n_1461),
.Y(n_1541)
);

AOI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1475),
.A2(n_1463),
.B1(n_1466),
.B2(n_1472),
.C(n_1469),
.Y(n_1542)
);

AO32x2_ASAP7_75t_L g1543 ( 
.A1(n_1434),
.A2(n_1473),
.A3(n_1448),
.B1(n_1456),
.B2(n_1430),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1477),
.A2(n_1432),
.B(n_1478),
.C(n_1445),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1445),
.B(n_1477),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1429),
.A2(n_1503),
.B1(n_1496),
.B2(n_1443),
.Y(n_1546)
);

AO32x2_ASAP7_75t_L g1547 ( 
.A1(n_1448),
.A2(n_1456),
.A3(n_1469),
.B1(n_1433),
.B2(n_1466),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1480),
.B(n_1484),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1463),
.A2(n_1436),
.B1(n_1457),
.B2(n_1470),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1492),
.Y(n_1550)
);

AOI221xp5_ASAP7_75t_L g1551 ( 
.A1(n_1469),
.A2(n_1444),
.B1(n_1495),
.B2(n_1490),
.C(n_1487),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_SL g1552 ( 
.A1(n_1505),
.A2(n_1502),
.B1(n_1443),
.B2(n_1470),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1461),
.A2(n_1441),
.B(n_1499),
.Y(n_1553)
);

AOI221xp5_ASAP7_75t_L g1554 ( 
.A1(n_1486),
.A2(n_1490),
.B1(n_1493),
.B2(n_1491),
.C(n_1487),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1553),
.B(n_1541),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1542),
.B(n_1458),
.Y(n_1556)
);

NOR2x1_ASAP7_75t_L g1557 ( 
.A(n_1522),
.B(n_1492),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1542),
.B(n_1458),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1509),
.B(n_1452),
.Y(n_1559)
);

CKINVDCx14_ASAP7_75t_R g1560 ( 
.A(n_1537),
.Y(n_1560)
);

INVxp67_ASAP7_75t_SL g1561 ( 
.A(n_1531),
.Y(n_1561)
);

BUFx2_ASAP7_75t_L g1562 ( 
.A(n_1543),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1527),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1527),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1543),
.B(n_1467),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1543),
.B(n_1499),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1531),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1543),
.B(n_1471),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1547),
.B(n_1544),
.Y(n_1569)
);

INVxp67_ASAP7_75t_SL g1570 ( 
.A(n_1550),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1539),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1547),
.B(n_1471),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1533),
.B(n_1454),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1548),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1547),
.B(n_1447),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1544),
.B(n_1545),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1554),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1515),
.A2(n_1485),
.B1(n_1513),
.B2(n_1534),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1552),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1561),
.B(n_1551),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1566),
.B(n_1551),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1563),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1571),
.Y(n_1583)
);

NAND3xp33_ASAP7_75t_L g1584 ( 
.A(n_1577),
.B(n_1508),
.C(n_1528),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1563),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1562),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1564),
.Y(n_1587)
);

OAI33xp33_ASAP7_75t_L g1588 ( 
.A1(n_1577),
.A2(n_1508),
.A3(n_1511),
.B1(n_1538),
.B2(n_1546),
.B3(n_1507),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1555),
.A2(n_1465),
.B(n_1522),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1566),
.B(n_1517),
.Y(n_1590)
);

BUFx12f_ASAP7_75t_L g1591 ( 
.A(n_1579),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1575),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1578),
.A2(n_1513),
.B1(n_1485),
.B2(n_1518),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1569),
.B(n_1512),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1575),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1561),
.B(n_1520),
.Y(n_1596)
);

OR2x6_ASAP7_75t_L g1597 ( 
.A(n_1569),
.B(n_1515),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1575),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1569),
.B(n_1450),
.Y(n_1599)
);

AND4x1_ASAP7_75t_L g1600 ( 
.A(n_1557),
.B(n_1529),
.C(n_1549),
.D(n_1514),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1579),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1565),
.B(n_1572),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1562),
.B(n_1440),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1567),
.B(n_1520),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1599),
.B(n_1556),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1602),
.B(n_1572),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1602),
.B(n_1572),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1582),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1582),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1583),
.B(n_1567),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1592),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1599),
.B(n_1556),
.Y(n_1612)
);

INVxp67_ASAP7_75t_SL g1613 ( 
.A(n_1596),
.Y(n_1613)
);

NOR2x1_ASAP7_75t_L g1614 ( 
.A(n_1580),
.B(n_1557),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1583),
.Y(n_1615)
);

AO21x1_ASAP7_75t_SL g1616 ( 
.A1(n_1580),
.A2(n_1558),
.B(n_1586),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1591),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1599),
.B(n_1558),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1602),
.B(n_1568),
.Y(n_1619)
);

BUFx2_ASAP7_75t_SL g1620 ( 
.A(n_1583),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1602),
.B(n_1568),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1586),
.B(n_1559),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1583),
.B(n_1570),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1591),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1582),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1592),
.B(n_1568),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1595),
.B(n_1576),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1603),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1595),
.B(n_1576),
.Y(n_1629)
);

AOI21xp33_ASAP7_75t_L g1630 ( 
.A1(n_1584),
.A2(n_1540),
.B(n_1510),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1595),
.B(n_1576),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1599),
.B(n_1574),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1585),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1585),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1585),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1598),
.B(n_1570),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1587),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1605),
.B(n_1596),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1630),
.B(n_1594),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1608),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1608),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1628),
.Y(n_1642)
);

O2A1O1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1630),
.A2(n_1584),
.B(n_1588),
.C(n_1580),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1609),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1609),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1605),
.B(n_1596),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1619),
.B(n_1590),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1616),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1612),
.B(n_1604),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1619),
.B(n_1621),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1625),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1625),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1619),
.B(n_1590),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1621),
.B(n_1590),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1633),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1613),
.B(n_1617),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1612),
.B(n_1604),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1613),
.B(n_1594),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1633),
.Y(n_1659)
);

NOR2x1_ASAP7_75t_L g1660 ( 
.A(n_1624),
.B(n_1584),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1634),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1628),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1611),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1634),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1621),
.B(n_1590),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1611),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1618),
.B(n_1632),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1635),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1606),
.B(n_1597),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1611),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1614),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1635),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1637),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1637),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1632),
.Y(n_1675)
);

NAND2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1614),
.B(n_1600),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1618),
.B(n_1604),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1636),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1606),
.B(n_1597),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1617),
.B(n_1560),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1676),
.B(n_1624),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1663),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1676),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1680),
.B(n_1624),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1676),
.B(n_1616),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1663),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1645),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1650),
.B(n_1616),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1643),
.B(n_1573),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1650),
.B(n_1606),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1648),
.A2(n_1588),
.B1(n_1581),
.B2(n_1601),
.C(n_1593),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1645),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1666),
.Y(n_1693)
);

OAI21xp33_ASAP7_75t_L g1694 ( 
.A1(n_1660),
.A2(n_1639),
.B(n_1671),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1651),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1675),
.B(n_1581),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1656),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1638),
.B(n_1622),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1638),
.B(n_1622),
.Y(n_1699)
);

AND3x1_ASAP7_75t_L g1700 ( 
.A(n_1669),
.B(n_1529),
.C(n_1581),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1666),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1669),
.B(n_1679),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1646),
.B(n_1600),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1651),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1642),
.Y(n_1705)
);

NOR2xp67_ASAP7_75t_L g1706 ( 
.A(n_1662),
.B(n_1601),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1647),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1646),
.B(n_1622),
.Y(n_1708)
);

INVx2_ASAP7_75t_SL g1709 ( 
.A(n_1678),
.Y(n_1709)
);

NAND4xp25_ASAP7_75t_L g1710 ( 
.A(n_1658),
.B(n_1593),
.C(n_1581),
.D(n_1532),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1652),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1649),
.B(n_1594),
.Y(n_1712)
);

O2A1O1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1649),
.A2(n_1677),
.B(n_1657),
.C(n_1579),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1675),
.B(n_1627),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1657),
.B(n_1594),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1679),
.B(n_1607),
.Y(n_1716)
);

INVx2_ASAP7_75t_SL g1717 ( 
.A(n_1683),
.Y(n_1717)
);

OAI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1710),
.A2(n_1597),
.B1(n_1591),
.B2(n_1667),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1694),
.A2(n_1703),
.B1(n_1689),
.B2(n_1691),
.C(n_1697),
.Y(n_1719)
);

INVxp67_ASAP7_75t_L g1720 ( 
.A(n_1683),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1694),
.A2(n_1678),
.B1(n_1677),
.B2(n_1664),
.C(n_1644),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1705),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1684),
.B(n_1457),
.Y(n_1723)
);

AOI21xp33_ASAP7_75t_L g1724 ( 
.A1(n_1685),
.A2(n_1591),
.B(n_1667),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1707),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1709),
.Y(n_1726)
);

AOI21xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1685),
.A2(n_1546),
.B(n_1526),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1688),
.B(n_1647),
.Y(n_1728)
);

NAND4xp75_ASAP7_75t_L g1729 ( 
.A(n_1681),
.B(n_1457),
.C(n_1600),
.D(n_1530),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1706),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1700),
.A2(n_1597),
.B1(n_1653),
.B2(n_1654),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1697),
.B(n_1681),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1688),
.B(n_1653),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1706),
.A2(n_1589),
.B(n_1640),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1710),
.A2(n_1589),
.B(n_1641),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1709),
.Y(n_1736)
);

INVx1_ASAP7_75t_SL g1737 ( 
.A(n_1683),
.Y(n_1737)
);

AOI322xp5_ASAP7_75t_L g1738 ( 
.A1(n_1696),
.A2(n_1607),
.A3(n_1627),
.B1(n_1629),
.B2(n_1631),
.C1(n_1665),
.C2(n_1654),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1702),
.A2(n_1597),
.B1(n_1515),
.B2(n_1631),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1707),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1700),
.A2(n_1597),
.B1(n_1631),
.B2(n_1629),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1707),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1726),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1726),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1736),
.Y(n_1745)
);

AOI211x1_ASAP7_75t_L g1746 ( 
.A1(n_1718),
.A2(n_1696),
.B(n_1702),
.C(n_1714),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1736),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1728),
.B(n_1716),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1728),
.B(n_1716),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1737),
.B(n_1713),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1732),
.B(n_1712),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1723),
.B(n_1457),
.Y(n_1752)
);

OAI332xp33_ASAP7_75t_L g1753 ( 
.A1(n_1722),
.A2(n_1687),
.A3(n_1692),
.B1(n_1711),
.B2(n_1695),
.B3(n_1704),
.C1(n_1699),
.C2(n_1698),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1719),
.A2(n_1707),
.B1(n_1597),
.B2(n_1715),
.Y(n_1754)
);

XNOR2x2_ASAP7_75t_L g1755 ( 
.A(n_1729),
.B(n_1698),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1722),
.B(n_1714),
.Y(n_1756)
);

NAND4xp25_ASAP7_75t_L g1757 ( 
.A(n_1721),
.B(n_1516),
.C(n_1687),
.D(n_1704),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1720),
.B(n_1690),
.Y(n_1758)
);

OAI221xp5_ASAP7_75t_SL g1759 ( 
.A1(n_1741),
.A2(n_1708),
.B1(n_1699),
.B2(n_1597),
.C(n_1690),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1717),
.B(n_1708),
.Y(n_1760)
);

AOI32xp33_ASAP7_75t_L g1761 ( 
.A1(n_1731),
.A2(n_1627),
.A3(n_1629),
.B1(n_1695),
.B2(n_1711),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1717),
.B(n_1665),
.Y(n_1762)
);

INVx1_ASAP7_75t_SL g1763 ( 
.A(n_1755),
.Y(n_1763)
);

NAND3xp33_ASAP7_75t_L g1764 ( 
.A(n_1746),
.B(n_1730),
.C(n_1724),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1748),
.B(n_1733),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1757),
.A2(n_1729),
.B1(n_1733),
.B2(n_1739),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1743),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1750),
.A2(n_1727),
.B1(n_1735),
.B2(n_1734),
.Y(n_1768)
);

NOR2x1_ASAP7_75t_L g1769 ( 
.A(n_1744),
.B(n_1725),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1749),
.B(n_1725),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1762),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1762),
.B(n_1740),
.Y(n_1772)
);

A2O1A1Ixp33_ASAP7_75t_L g1773 ( 
.A1(n_1757),
.A2(n_1738),
.B(n_1740),
.C(n_1742),
.Y(n_1773)
);

INVxp67_ASAP7_75t_SL g1774 ( 
.A(n_1760),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1763),
.B(n_1753),
.Y(n_1775)
);

NOR3xp33_ASAP7_75t_L g1776 ( 
.A(n_1763),
.B(n_1753),
.C(n_1754),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1765),
.B(n_1758),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1764),
.B(n_1747),
.C(n_1745),
.Y(n_1778)
);

CKINVDCx14_ASAP7_75t_R g1779 ( 
.A(n_1771),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1769),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1768),
.B(n_1761),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1770),
.B(n_1772),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_L g1783 ( 
.A(n_1773),
.B(n_1759),
.C(n_1756),
.Y(n_1783)
);

NOR3x1_ASAP7_75t_L g1784 ( 
.A(n_1774),
.B(n_1751),
.C(n_1692),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1767),
.Y(n_1785)
);

NAND4xp25_ASAP7_75t_L g1786 ( 
.A(n_1776),
.B(n_1766),
.C(n_1752),
.D(n_1768),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_SL g1787 ( 
.A(n_1782),
.B(n_1742),
.Y(n_1787)
);

AOI222xp33_ASAP7_75t_L g1788 ( 
.A1(n_1775),
.A2(n_1701),
.B1(n_1693),
.B2(n_1686),
.C1(n_1682),
.C2(n_1674),
.Y(n_1788)
);

AOI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1776),
.A2(n_1701),
.B1(n_1693),
.B2(n_1686),
.C(n_1682),
.Y(n_1789)
);

OAI211xp5_ASAP7_75t_L g1790 ( 
.A1(n_1781),
.A2(n_1460),
.B(n_1693),
.C(n_1686),
.Y(n_1790)
);

OAI211xp5_ASAP7_75t_L g1791 ( 
.A1(n_1786),
.A2(n_1778),
.B(n_1780),
.C(n_1779),
.Y(n_1791)
);

AOI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1790),
.A2(n_1783),
.B1(n_1777),
.B2(n_1785),
.C(n_1784),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1787),
.B(n_1682),
.Y(n_1793)
);

AOI221x1_ASAP7_75t_L g1794 ( 
.A1(n_1788),
.A2(n_1701),
.B1(n_1674),
.B2(n_1673),
.C(n_1672),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1789),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1787),
.B(n_1668),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1792),
.B(n_1607),
.Y(n_1797)
);

NOR3xp33_ASAP7_75t_L g1798 ( 
.A(n_1791),
.B(n_1535),
.C(n_1536),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1793),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1795),
.B(n_1626),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_SL g1801 ( 
.A1(n_1796),
.A2(n_1620),
.B1(n_1519),
.B2(n_1524),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1797),
.B(n_1800),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1799),
.B(n_1794),
.Y(n_1803)
);

NAND4xp75_ASAP7_75t_L g1804 ( 
.A(n_1801),
.B(n_1615),
.C(n_1672),
.D(n_1661),
.Y(n_1804)
);

NAND3xp33_ASAP7_75t_SL g1805 ( 
.A(n_1803),
.B(n_1798),
.C(n_1525),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1805),
.A2(n_1802),
.B1(n_1804),
.B2(n_1670),
.Y(n_1806)
);

INVxp33_ASAP7_75t_SL g1807 ( 
.A(n_1806),
.Y(n_1807)
);

XNOR2xp5_ASAP7_75t_L g1808 ( 
.A(n_1806),
.B(n_1521),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1807),
.A2(n_1670),
.B1(n_1620),
.B2(n_1615),
.Y(n_1809)
);

CKINVDCx20_ASAP7_75t_R g1810 ( 
.A(n_1808),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1809),
.B(n_1615),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1810),
.A2(n_1655),
.B(n_1652),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1811),
.A2(n_1673),
.B1(n_1661),
.B2(n_1659),
.Y(n_1813)
);

OA21x2_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1812),
.B(n_1659),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1814),
.Y(n_1815)
);

AOI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1815),
.A2(n_1655),
.B1(n_1623),
.B2(n_1610),
.C(n_1524),
.Y(n_1816)
);

AOI211xp5_ASAP7_75t_L g1817 ( 
.A1(n_1816),
.A2(n_1519),
.B(n_1524),
.C(n_1523),
.Y(n_1817)
);


endmodule