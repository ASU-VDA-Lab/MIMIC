module fake_jpeg_7954_n_227 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_35),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

NOR2x1_ASAP7_75t_R g57 ( 
.A(n_36),
.B(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_40),
.B(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_20),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_42),
.B1(n_36),
.B2(n_20),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_33),
.B1(n_32),
.B2(n_43),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_20),
.B1(n_26),
.B2(n_23),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_25),
.B1(n_24),
.B2(n_29),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_62),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_26),
.Y(n_59)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_17),
.C(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_24),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_22),
.Y(n_83)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_69),
.B(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_73),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_80),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_26),
.B1(n_23),
.B2(n_17),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_75),
.A2(n_76),
.B1(n_7),
.B2(n_8),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_18),
.B1(n_28),
.B2(n_21),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_22),
.B1(n_34),
.B2(n_25),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_33),
.B1(n_32),
.B2(n_64),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_98),
.B(n_3),
.C(n_4),
.Y(n_106)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_47),
.B(n_21),
.C(n_34),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_85),
.B1(n_86),
.B2(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_83),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_1),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_94),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_1),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_33),
.B1(n_32),
.B2(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_97),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_115),
.B1(n_116),
.B2(n_120),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_102),
.B(n_111),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_16),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_11),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_33),
.B1(n_32),
.B2(n_45),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_119),
.B1(n_95),
.B2(n_91),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_45),
.B(n_4),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_94),
.B(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_10),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_3),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_114),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_73),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_5),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_14),
.B1(n_12),
.B2(n_9),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_9),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_94),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_109),
.B1(n_121),
.B2(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_124),
.B(n_128),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_74),
.B1(n_91),
.B2(n_71),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_132),
.B(n_134),
.Y(n_153)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_73),
.Y(n_130)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_138),
.Y(n_156)
);

OR2x2_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_68),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_10),
.B(n_11),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_97),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_139),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_116),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_71),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_77),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_142),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_110),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_77),
.Y(n_144)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_84),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_103),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_152),
.C(n_155),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_127),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_150),
.B(n_123),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_99),
.C(n_113),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_105),
.C(n_107),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_163),
.C(n_134),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_107),
.C(n_101),
.Y(n_163)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_172),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_143),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_171),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_126),
.C(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

OAI321xp33_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_126),
.A3(n_133),
.B1(n_124),
.B2(n_106),
.C(n_129),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_153),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_138),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_177),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_147),
.C(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_180),
.A2(n_181),
.B(n_182),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_131),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_189),
.C(n_179),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_183),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_164),
.C(n_152),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_148),
.B1(n_125),
.B2(n_158),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_168),
.B1(n_180),
.B2(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_200),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_203),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_175),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_201),
.C(n_204),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_153),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_194),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_202),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_169),
.B1(n_182),
.B2(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_178),
.C(n_155),
.Y(n_204)
);

AOI21x1_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_192),
.B(n_188),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_206),
.A2(n_193),
.B(n_146),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_211),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_185),
.C(n_184),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_212),
.B(n_213),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_202),
.A3(n_195),
.B1(n_185),
.B2(n_190),
.C1(n_193),
.C2(n_201),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_205),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_190),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_154),
.B(n_141),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_157),
.C(n_118),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_220),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_215),
.A2(n_210),
.B(n_197),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_154),
.C(n_114),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_222),
.C(n_114),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_224),
.B(n_225),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_84),
.B(n_137),
.C(n_88),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_93),
.Y(n_227)
);


endmodule