module fake_netlist_6_4039_n_2211 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2211);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2211;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_1159;
wire n_276;
wire n_995;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2052;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_54),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_132),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_98),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_179),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_31),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_4),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_101),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_146),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_42),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_190),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_39),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_111),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_194),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_16),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_33),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_77),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_45),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_25),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_151),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_105),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_85),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_155),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_106),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_96),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_176),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_68),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_72),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_18),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_136),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_181),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_133),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_187),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_149),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_213),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_171),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_50),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_66),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_202),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_49),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_109),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_39),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_157),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_1),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_56),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_26),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_154),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_112),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_75),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_99),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_124),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_69),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_9),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_51),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_85),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_121),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_25),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_158),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_118),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_13),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_72),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_162),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_19),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_11),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_209),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_167),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_90),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_200),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_3),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_160),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_6),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_174),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_218),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_82),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_89),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_100),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_172),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_135),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_1),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_168),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_35),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_198),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_55),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_142),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_108),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_33),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_166),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_113),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_97),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_70),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_8),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_139),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_0),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_18),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_183),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_87),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_67),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_65),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_73),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_66),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_47),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_28),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_114),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_49),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_56),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_10),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_140),
.Y(n_329)
);

BUFx5_ASAP7_75t_L g330 ( 
.A(n_3),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_26),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_88),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_77),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_8),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_4),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_145),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_11),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_75),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_70),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_92),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_93),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_63),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_102),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_148),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_192),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_34),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_134),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_207),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_116),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_10),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_27),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_24),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_120),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_82),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_141),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_215),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_117),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_51),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_150),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_95),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_9),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_47),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_138),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_40),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_186),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_208),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_211),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_60),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_54),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_0),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_177),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_60),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_52),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_83),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_74),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_42),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_76),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_48),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_5),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_23),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_203),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_217),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_74),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_175),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_69),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_193),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_119),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_104),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_5),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_214),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_48),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_83),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_195),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_204),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_165),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_27),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_156),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_159),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_127),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_137),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_22),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_164),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_131),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_196),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_94),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_13),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_52),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_23),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_34),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_110),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_43),
.Y(n_411)
);

BUFx10_ASAP7_75t_L g412 ( 
.A(n_125),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_115),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_169),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_43),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_22),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_126),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_65),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_128),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_7),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_216),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_76),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_67),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_180),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_20),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_31),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_41),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_123),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_143),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_153),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_44),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_30),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_30),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_170),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_224),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_234),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_232),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_241),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_225),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_330),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_330),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_295),
.Y(n_442)
);

INVxp33_ASAP7_75t_L g443 ( 
.A(n_378),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_228),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_330),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_231),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_245),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_330),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_221),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_330),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_330),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_226),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_330),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_330),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_330),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_295),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_279),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_279),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_279),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_279),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_237),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_279),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_237),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_256),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_282),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_282),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_282),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_306),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_246),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_282),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_250),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_233),
.B(n_2),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_282),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_233),
.B(n_2),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_291),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_331),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_255),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_331),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_331),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_259),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_264),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_331),
.Y(n_483)
);

INVxp33_ASAP7_75t_SL g484 ( 
.A(n_227),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_252),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_220),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_220),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_269),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_271),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_272),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_331),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_260),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_369),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_280),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_260),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_380),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_380),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_401),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_281),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_353),
.B(n_6),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_288),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_230),
.B(n_7),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_289),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_222),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_292),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_230),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_237),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_309),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_222),
.Y(n_512)
);

INVxp33_ASAP7_75t_L g513 ( 
.A(n_242),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_235),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_242),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_266),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_266),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_267),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_267),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_270),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_294),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_244),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_270),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_311),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_297),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_229),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_229),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_299),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_240),
.Y(n_529)
);

CKINVDCx14_ASAP7_75t_R g530 ( 
.A(n_223),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_301),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_301),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_240),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_243),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_303),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_363),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_303),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_300),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_402),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_424),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_315),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_304),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_315),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_316),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_316),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_236),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_321),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_314),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_253),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_317),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_254),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_458),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_446),
.A2(n_443),
.B1(n_505),
.B2(n_319),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_458),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_459),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_459),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_512),
.B(n_329),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_489),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_442),
.B(n_425),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_522),
.B(n_318),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_460),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_484),
.B(n_353),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_483),
.B(n_325),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_452),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_452),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_489),
.B(n_336),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_489),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_440),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_460),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_461),
.Y(n_570)
);

BUFx8_ASAP7_75t_L g571 ( 
.A(n_450),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_489),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_489),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_457),
.B(n_343),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_435),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_440),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_441),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_439),
.B(n_340),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_473),
.B(n_344),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_461),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_513),
.B(n_425),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_476),
.B(n_321),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_441),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_463),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_463),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_445),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_466),
.Y(n_587)
);

AND2x2_ASAP7_75t_SL g588 ( 
.A(n_475),
.B(n_271),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_500),
.B(n_466),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_516),
.B(n_322),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_449),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_467),
.B(n_348),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_449),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_467),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_468),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_451),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_451),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_468),
.B(n_345),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_471),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_471),
.B(n_355),
.Y(n_601)
);

AND2x2_ASAP7_75t_SL g602 ( 
.A(n_505),
.B(n_348),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_514),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_474),
.B(n_243),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_474),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_477),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_477),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_479),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_454),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_454),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_479),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_480),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_455),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_480),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_491),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_455),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_491),
.B(n_251),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_456),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_486),
.B(n_251),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_444),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_487),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_456),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_533),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_533),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_507),
.B(n_262),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_534),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_509),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_534),
.Y(n_628)
);

NOR2x1_ASAP7_75t_L g629 ( 
.A(n_485),
.B(n_262),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_509),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_492),
.Y(n_631)
);

INVx6_ASAP7_75t_L g632 ( 
.A(n_485),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_515),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_526),
.B(n_268),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_492),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_527),
.B(n_356),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_495),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_495),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_515),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_496),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_517),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_529),
.B(n_268),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_578),
.B(n_447),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_564),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_568),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_562),
.B(n_448),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_558),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_564),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_602),
.A2(n_588),
.B1(n_559),
.B2(n_579),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_581),
.B(n_470),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_568),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_568),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_583),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_564),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_574),
.B(n_472),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_583),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_602),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_574),
.B(n_478),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_583),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_582),
.B(n_450),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_565),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_602),
.A2(n_453),
.B1(n_337),
.B2(n_352),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_609),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_563),
.B(n_481),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_558),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_619),
.B(n_278),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_609),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_609),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_565),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_565),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_603),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_610),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_610),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_610),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_559),
.B(n_496),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_558),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_613),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_613),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_613),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_576),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_579),
.B(n_482),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_588),
.A2(n_551),
.B1(n_549),
.B2(n_488),
.Y(n_682)
);

BUFx10_ASAP7_75t_L g683 ( 
.A(n_632),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_622),
.Y(n_684)
);

INVx5_ASAP7_75t_L g685 ( 
.A(n_576),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_581),
.B(n_490),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_622),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_563),
.B(n_494),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_622),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_632),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_588),
.A2(n_453),
.B1(n_337),
.B2(n_352),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_595),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_619),
.B(n_497),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_619),
.A2(n_376),
.B1(n_377),
.B2(n_322),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_619),
.B(n_497),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_595),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_576),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_558),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_576),
.Y(n_699)
);

INVx4_ASAP7_75t_L g700 ( 
.A(n_576),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_595),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_576),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_577),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_576),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_577),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_566),
.B(n_499),
.Y(n_706)
);

AND2x6_ASAP7_75t_L g707 ( 
.A(n_577),
.B(n_278),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_632),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_557),
.A2(n_530),
.B1(n_506),
.B2(n_508),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_632),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_625),
.A2(n_377),
.B1(n_385),
.B2(n_376),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_586),
.Y(n_712)
);

INVx8_ASAP7_75t_L g713 ( 
.A(n_557),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_632),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_586),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_557),
.B(n_504),
.Y(n_716)
);

INVxp33_ASAP7_75t_SL g717 ( 
.A(n_603),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_575),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_586),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_577),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_586),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_566),
.B(n_521),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_582),
.B(n_437),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_597),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_597),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_586),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_558),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_597),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_597),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_558),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_558),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_586),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_599),
.B(n_525),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_586),
.Y(n_734)
);

CKINVDCx16_ASAP7_75t_R g735 ( 
.A(n_553),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_572),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_620),
.B(n_528),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_629),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_623),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_625),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_623),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_621),
.Y(n_742)
);

INVx4_ASAP7_75t_SL g743 ( 
.A(n_590),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_572),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_572),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_590),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_572),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_590),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_599),
.B(n_538),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_601),
.B(n_542),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_620),
.B(n_548),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_552),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_552),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_601),
.B(n_550),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_590),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_620),
.B(n_493),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_590),
.Y(n_757)
);

BUFx10_ASAP7_75t_L g758 ( 
.A(n_625),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_572),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_590),
.Y(n_760)
);

NOR3xp33_ASAP7_75t_L g761 ( 
.A(n_553),
.B(n_464),
.C(n_462),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_572),
.Y(n_762)
);

BUFx10_ASAP7_75t_L g763 ( 
.A(n_625),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_590),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_589),
.B(n_546),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_620),
.B(n_629),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_554),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_592),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_636),
.B(n_510),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_592),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_560),
.B(n_252),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_554),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_592),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_636),
.B(n_532),
.C(n_531),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_572),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_592),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_555),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_589),
.B(n_436),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_621),
.B(n_438),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_592),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_621),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_591),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_592),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_567),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_573),
.B(n_434),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_592),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_567),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_567),
.Y(n_788)
);

INVx5_ASAP7_75t_L g789 ( 
.A(n_594),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_594),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_555),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_642),
.B(n_465),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_642),
.B(n_469),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_571),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_591),
.Y(n_795)
);

OR2x6_ASAP7_75t_L g796 ( 
.A(n_634),
.B(n_284),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_594),
.Y(n_797)
);

INVxp67_ASAP7_75t_SL g798 ( 
.A(n_567),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_795),
.B(n_511),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_683),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_657),
.B(n_649),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_769),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_683),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_657),
.B(n_594),
.Y(n_804)
);

INVxp33_ASAP7_75t_L g805 ( 
.A(n_660),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_739),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_675),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_738),
.B(n_782),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_738),
.B(n_594),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_739),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_681),
.B(n_594),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_655),
.B(n_594),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_658),
.B(n_598),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_782),
.B(n_598),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_692),
.Y(n_815)
);

AND2x6_ASAP7_75t_SL g816 ( 
.A(n_643),
.B(n_385),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_778),
.B(n_524),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_740),
.B(n_758),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_742),
.B(n_634),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_742),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_664),
.B(n_598),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_740),
.B(n_598),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_688),
.B(n_536),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_706),
.B(n_598),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_722),
.B(n_598),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_692),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_741),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_733),
.B(n_539),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_741),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_776),
.Y(n_830)
);

INVx8_ASAP7_75t_L g831 ( 
.A(n_713),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_749),
.B(n_598),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_750),
.B(n_616),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_754),
.B(n_616),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_644),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_696),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_765),
.B(n_540),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_696),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_701),
.B(n_616),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_740),
.B(n_616),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_703),
.A2(n_573),
.B(n_604),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_701),
.B(n_616),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_675),
.B(n_713),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_784),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_742),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_693),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_693),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_644),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_713),
.B(n_616),
.Y(n_849)
);

NAND3xp33_ASAP7_75t_L g850 ( 
.A(n_691),
.B(n_571),
.C(n_634),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_644),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_695),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_794),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_695),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_713),
.B(n_798),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_666),
.A2(n_642),
.B1(n_634),
.B2(n_604),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_713),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_740),
.B(n_616),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_SL g859 ( 
.A(n_662),
.B(n_285),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_666),
.B(n_618),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_666),
.B(n_618),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_666),
.B(n_618),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_752),
.B(n_753),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_752),
.B(n_618),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_753),
.B(n_618),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_648),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_767),
.B(n_772),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_671),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_781),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_758),
.B(n_618),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_758),
.B(n_618),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_767),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_758),
.B(n_763),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_716),
.A2(n_642),
.B1(n_617),
.B2(n_604),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_772),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_777),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_777),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_660),
.B(n_627),
.Y(n_878)
);

O2A1O1Ixp5_ASAP7_75t_L g879 ( 
.A1(n_703),
.A2(n_604),
.B(n_617),
.C(n_593),
.Y(n_879)
);

NAND2xp33_ASAP7_75t_L g880 ( 
.A(n_707),
.B(n_284),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_791),
.B(n_573),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_796),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_791),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_705),
.B(n_617),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_763),
.B(n_624),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_705),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_720),
.B(n_617),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_796),
.A2(n_707),
.B1(n_645),
.B2(n_652),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_720),
.B(n_593),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_671),
.B(n_627),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_646),
.B(n_571),
.Y(n_891)
);

NAND2xp33_ASAP7_75t_L g892 ( 
.A(n_707),
.B(n_287),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_724),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_724),
.B(n_593),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_690),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_648),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_763),
.B(n_725),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_796),
.A2(n_593),
.B1(n_287),
.B2(n_298),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_648),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_728),
.B(n_556),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_717),
.B(n_571),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_728),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_729),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_650),
.B(n_238),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_792),
.A2(n_365),
.B1(n_366),
.B2(n_357),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_729),
.B(n_556),
.Y(n_906)
);

NAND2xp33_ASAP7_75t_L g907 ( 
.A(n_707),
.B(n_290),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_763),
.B(n_624),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_737),
.B(n_561),
.Y(n_909)
);

INVxp33_ASAP7_75t_L g910 ( 
.A(n_723),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_654),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_751),
.B(n_561),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_784),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_785),
.B(n_569),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_654),
.Y(n_915)
);

NOR3xp33_ASAP7_75t_L g916 ( 
.A(n_735),
.B(n_793),
.C(n_779),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_697),
.B(n_624),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_784),
.B(n_569),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_787),
.B(n_570),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_697),
.B(n_624),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_787),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_756),
.B(n_630),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_654),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_766),
.A2(n_371),
.B1(n_381),
.B2(n_367),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_796),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_787),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_661),
.Y(n_927)
);

AOI221xp5_ASAP7_75t_L g928 ( 
.A1(n_735),
.A2(n_761),
.B1(n_346),
.B2(n_354),
.C(n_339),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_788),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_788),
.B(n_570),
.Y(n_930)
);

BUFx10_ASAP7_75t_L g931 ( 
.A(n_707),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_690),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_788),
.B(n_580),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_645),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_723),
.B(n_630),
.Y(n_935)
);

AND2x2_ASAP7_75t_SL g936 ( 
.A(n_694),
.B(n_290),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_686),
.B(n_239),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_708),
.B(n_710),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_697),
.B(n_624),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_699),
.B(n_624),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_796),
.A2(n_639),
.B(n_641),
.C(n_633),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_709),
.B(n_247),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_708),
.B(n_580),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_682),
.B(n_633),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_651),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_774),
.A2(n_298),
.B1(n_307),
.B2(n_302),
.Y(n_946)
);

INVx8_ASAP7_75t_L g947 ( 
.A(n_707),
.Y(n_947)
);

NAND2xp33_ASAP7_75t_L g948 ( 
.A(n_707),
.B(n_302),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_651),
.A2(n_641),
.B(n_639),
.C(n_652),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_771),
.B(n_248),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_710),
.B(n_584),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_776),
.B(n_584),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_707),
.A2(n_384),
.B1(n_386),
.B2(n_382),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_776),
.B(n_585),
.Y(n_954)
);

NAND3xp33_ASAP7_75t_L g955 ( 
.A(n_711),
.B(n_257),
.C(n_249),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_653),
.A2(n_307),
.B1(n_341),
.B2(n_310),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_699),
.B(n_624),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_776),
.B(n_585),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_699),
.B(n_628),
.Y(n_959)
);

NAND2x1p5_ASAP7_75t_L g960 ( 
.A(n_680),
.B(n_310),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_718),
.B(n_258),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_680),
.B(n_263),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_661),
.Y(n_963)
);

BUFx12f_ASAP7_75t_SL g964 ( 
.A(n_730),
.Y(n_964)
);

BUFx8_ASAP7_75t_L g965 ( 
.A(n_702),
.Y(n_965)
);

NOR2xp67_ASAP7_75t_L g966 ( 
.A(n_669),
.B(n_637),
.Y(n_966)
);

OAI22xp33_ASAP7_75t_L g967 ( 
.A1(n_653),
.A2(n_347),
.B1(n_360),
.B2(n_359),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_775),
.A2(n_626),
.B(n_623),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_702),
.B(n_628),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_661),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_835),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_802),
.B(n_656),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_800),
.A2(n_700),
.B(n_680),
.Y(n_973)
);

AO21x1_ASAP7_75t_L g974 ( 
.A1(n_801),
.A2(n_811),
.B(n_812),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_868),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_SL g976 ( 
.A1(n_801),
.A2(n_347),
.B(n_349),
.C(n_341),
.Y(n_976)
);

AO21x1_ASAP7_75t_L g977 ( 
.A1(n_813),
.A2(n_359),
.B(n_349),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_886),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_852),
.A2(n_393),
.B(n_394),
.C(n_360),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_890),
.B(n_517),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_852),
.A2(n_704),
.B1(n_712),
.B2(n_702),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_800),
.A2(n_700),
.B(n_680),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_843),
.A2(n_712),
.B1(n_715),
.B2(n_704),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_909),
.B(n_656),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_859),
.A2(n_394),
.B(n_403),
.C(n_393),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_832),
.B(n_704),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_912),
.B(n_659),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_922),
.B(n_659),
.Y(n_988)
);

OAI21xp33_ASAP7_75t_L g989 ( 
.A1(n_942),
.A2(n_273),
.B(n_265),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_935),
.B(n_518),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_859),
.A2(n_404),
.B(n_410),
.C(n_403),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_882),
.A2(n_410),
.B1(n_413),
.B2(n_404),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_820),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_882),
.A2(n_925),
.B1(n_804),
.B2(n_856),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_807),
.A2(n_414),
.B(n_417),
.C(n_413),
.Y(n_995)
);

OAI21xp33_ASAP7_75t_L g996 ( 
.A1(n_805),
.A2(n_276),
.B(n_274),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_800),
.A2(n_734),
.B(n_700),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_803),
.A2(n_734),
.B(n_700),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_807),
.B(n_663),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_835),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_805),
.B(n_799),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_803),
.A2(n_748),
.B(n_734),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_824),
.A2(n_757),
.B(n_748),
.Y(n_1003)
);

AND2x2_ASAP7_75t_SL g1004 ( 
.A(n_936),
.B(n_414),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_872),
.B(n_663),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_846),
.A2(n_668),
.B(n_673),
.C(n_667),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_825),
.A2(n_757),
.B(n_748),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_833),
.A2(n_834),
.B(n_821),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_848),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_849),
.A2(n_757),
.B(n_797),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_855),
.A2(n_757),
.B(n_797),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_822),
.A2(n_715),
.B(n_712),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_820),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_869),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_925),
.A2(n_429),
.B1(n_430),
.B2(n_417),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_819),
.B(n_715),
.Y(n_1016)
);

NOR2x1_ASAP7_75t_L g1017 ( 
.A(n_850),
.B(n_320),
.Y(n_1017)
);

NOR3xp33_ASAP7_75t_L g1018 ( 
.A(n_837),
.B(n_332),
.C(n_275),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_847),
.A2(n_668),
.B(n_673),
.C(n_667),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_822),
.A2(n_797),
.B(n_721),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_964),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_879),
.A2(n_679),
.B(n_677),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_875),
.B(n_677),
.Y(n_1023)
);

CKINVDCx10_ASAP7_75t_R g1024 ( 
.A(n_816),
.Y(n_1024)
);

INVx2_ASAP7_75t_SL g1025 ( 
.A(n_878),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_876),
.B(n_679),
.Y(n_1026)
);

NAND2xp33_ASAP7_75t_L g1027 ( 
.A(n_831),
.B(n_719),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_874),
.A2(n_430),
.B1(n_429),
.B2(n_719),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_877),
.B(n_883),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_840),
.A2(n_721),
.B(n_719),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_840),
.A2(n_790),
.B(n_726),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_820),
.Y(n_1032)
);

NOR2xp67_ASAP7_75t_L g1033 ( 
.A(n_891),
.B(n_689),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_848),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_858),
.A2(n_790),
.B(n_726),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_857),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_888),
.A2(n_726),
.B1(n_732),
.B2(n_721),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_858),
.A2(n_790),
.B(n_746),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_944),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_914),
.B(n_863),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_870),
.A2(n_746),
.B(n_732),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_819),
.B(n_732),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_870),
.A2(n_755),
.B(n_746),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_851),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_893),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_867),
.B(n_689),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_820),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_819),
.B(n_755),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_845),
.B(n_755),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_854),
.A2(n_764),
.B1(n_768),
.B2(n_760),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_871),
.A2(n_764),
.B(n_760),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_964),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_823),
.B(n_683),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_857),
.B(n_518),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_950),
.A2(n_764),
.B(n_768),
.C(n_760),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_853),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_828),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_910),
.B(n_407),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_871),
.A2(n_770),
.B(n_768),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_860),
.A2(n_773),
.B(n_770),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_817),
.B(n_519),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_861),
.A2(n_773),
.B(n_770),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_808),
.B(n_773),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_862),
.A2(n_908),
.B(n_885),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_808),
.Y(n_1065)
);

BUFx4f_ASAP7_75t_L g1066 ( 
.A(n_845),
.Y(n_1066)
);

AND2x2_ASAP7_75t_SL g1067 ( 
.A(n_936),
.B(n_916),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_902),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_946),
.A2(n_814),
.B(n_892),
.C(n_880),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_904),
.A2(n_780),
.B(n_786),
.C(n_783),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_885),
.A2(n_783),
.B(n_780),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_908),
.A2(n_783),
.B(n_780),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_815),
.B(n_786),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_884),
.A2(n_674),
.B(n_672),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_841),
.A2(n_786),
.B(n_731),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_826),
.B(n_672),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_809),
.A2(n_731),
.B(n_730),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_845),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_809),
.A2(n_731),
.B(n_730),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_903),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_845),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_938),
.A2(n_731),
.B(n_730),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_887),
.A2(n_674),
.B(n_672),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_910),
.B(n_519),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_937),
.A2(n_678),
.B(n_684),
.C(n_687),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_836),
.B(n_674),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_921),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_851),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_838),
.A2(n_898),
.B1(n_844),
.B2(n_814),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_L g1090 ( 
.A(n_928),
.B(n_283),
.C(n_277),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_866),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_941),
.A2(n_684),
.B(n_687),
.C(n_678),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_921),
.Y(n_1093)
);

OAI21xp33_ASAP7_75t_L g1094 ( 
.A1(n_961),
.A2(n_293),
.B(n_286),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_897),
.A2(n_731),
.B(n_730),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_897),
.A2(n_731),
.B(n_730),
.Y(n_1096)
);

OAI21xp33_ASAP7_75t_L g1097 ( 
.A1(n_905),
.A2(n_305),
.B(n_296),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_921),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_901),
.B(n_520),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_SL g1100 ( 
.A(n_965),
.B(n_411),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_913),
.B(n_678),
.Y(n_1101)
);

AND2x2_ASAP7_75t_SL g1102 ( 
.A(n_880),
.B(n_391),
.Y(n_1102)
);

NAND3xp33_ASAP7_75t_L g1103 ( 
.A(n_955),
.B(n_312),
.C(n_308),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_895),
.B(n_520),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_892),
.A2(n_684),
.B(n_687),
.C(n_596),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_864),
.A2(n_865),
.B(n_842),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_934),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_818),
.A2(n_744),
.B(n_736),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_866),
.Y(n_1109)
);

OAI321xp33_ASAP7_75t_L g1110 ( 
.A1(n_967),
.A2(n_422),
.A3(n_426),
.B1(n_433),
.B2(n_391),
.C(n_427),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_945),
.Y(n_1111)
);

CKINVDCx8_ASAP7_75t_R g1112 ( 
.A(n_921),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_818),
.A2(n_744),
.B(n_736),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_962),
.B(n_523),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_844),
.B(n_669),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_806),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_873),
.A2(n_744),
.B(n_736),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_844),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_806),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_873),
.A2(n_744),
.B(n_736),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_895),
.B(n_647),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_924),
.B(n_683),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_839),
.A2(n_744),
.B(n_736),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_SL g1124 ( 
.A1(n_831),
.A2(n_422),
.B1(n_427),
.B2(n_409),
.Y(n_1124)
);

AO21x1_ASAP7_75t_L g1125 ( 
.A1(n_960),
.A2(n_426),
.B(n_409),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_889),
.A2(n_744),
.B(n_736),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_931),
.B(n_714),
.Y(n_1127)
);

INVx11_ASAP7_75t_L g1128 ( 
.A(n_965),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_949),
.A2(n_670),
.B(n_762),
.C(n_759),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_810),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_926),
.B(n_929),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_894),
.A2(n_670),
.B(n_665),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_830),
.A2(n_747),
.B(n_685),
.Y(n_1133)
);

NOR3xp33_ASAP7_75t_L g1134 ( 
.A(n_907),
.B(n_323),
.C(n_313),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_965),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_918),
.A2(n_747),
.B(n_685),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_932),
.B(n_647),
.Y(n_1137)
);

BUFx8_ASAP7_75t_L g1138 ( 
.A(n_932),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_907),
.A2(n_587),
.B(n_596),
.C(n_600),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_827),
.B(n_647),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_919),
.B(n_523),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_896),
.A2(n_670),
.B(n_665),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_930),
.A2(n_747),
.B(n_685),
.Y(n_1143)
);

AO21x1_ASAP7_75t_L g1144 ( 
.A1(n_960),
.A2(n_433),
.B(n_587),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_827),
.Y(n_1145)
);

BUFx2_ASAP7_75t_SL g1146 ( 
.A(n_966),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_933),
.A2(n_747),
.B(n_685),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_947),
.A2(n_747),
.B(n_685),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_829),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_831),
.Y(n_1150)
);

NOR2xp67_ASAP7_75t_L g1151 ( 
.A(n_943),
.B(n_535),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_948),
.A2(n_611),
.B(n_600),
.C(n_605),
.Y(n_1152)
);

AO21x1_ASAP7_75t_L g1153 ( 
.A1(n_917),
.A2(n_606),
.B(n_605),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_931),
.B(n_714),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_896),
.B(n_665),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_831),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_899),
.B(n_676),
.Y(n_1157)
);

NOR3xp33_ASAP7_75t_L g1158 ( 
.A(n_948),
.B(n_326),
.C(n_324),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_951),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_899),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1008),
.A2(n_947),
.B(n_952),
.Y(n_1161)
);

OAI22x1_ASAP7_75t_L g1162 ( 
.A1(n_1057),
.A2(n_375),
.B1(n_328),
.B2(n_333),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1039),
.B(n_881),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1058),
.B(n_900),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1040),
.B(n_906),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1058),
.B(n_953),
.Y(n_1166)
);

INVx6_ASAP7_75t_L g1167 ( 
.A(n_1138),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1061),
.B(n_980),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1114),
.B(n_911),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_971),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_990),
.B(n_535),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1067),
.A2(n_428),
.B1(n_421),
.B2(n_387),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1004),
.A2(n_956),
.B1(n_947),
.B2(n_970),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_1036),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1014),
.Y(n_1175)
);

AND2x6_ASAP7_75t_L g1176 ( 
.A(n_1150),
.B(n_911),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1018),
.A2(n_947),
.B(n_954),
.C(n_958),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_988),
.B(n_915),
.Y(n_1178)
);

AND3x1_ASAP7_75t_SL g1179 ( 
.A(n_1024),
.B(n_541),
.C(n_537),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1099),
.B(n_931),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1004),
.A2(n_970),
.B1(n_963),
.B2(n_927),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_1025),
.B(n_915),
.Y(n_1182)
);

O2A1O1Ixp5_ASAP7_75t_L g1183 ( 
.A1(n_977),
.A2(n_1053),
.B(n_974),
.C(n_1122),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_972),
.B(n_923),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_SL g1185 ( 
.A1(n_1056),
.A2(n_361),
.B1(n_327),
.B2(n_334),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_975),
.B(n_1001),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1000),
.Y(n_1187)
);

AO21x1_ASAP7_75t_L g1188 ( 
.A1(n_1018),
.A2(n_939),
.B(n_920),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1112),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1067),
.B(n_714),
.Y(n_1190)
);

AOI21x1_ASAP7_75t_L g1191 ( 
.A1(n_986),
.A2(n_940),
.B(n_939),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1064),
.A2(n_927),
.B(n_923),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_975),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1107),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1111),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1009),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1084),
.B(n_537),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1102),
.A2(n_963),
.B1(n_351),
.B2(n_432),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1159),
.B(n_541),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_985),
.A2(n_969),
.B(n_959),
.C(n_957),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_984),
.B(n_968),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1102),
.A2(n_338),
.B1(n_431),
.B2(n_423),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_978),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_987),
.A2(n_335),
.B1(n_420),
.B2(n_342),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1138),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1104),
.B(n_543),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1021),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1034),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1141),
.B(n_676),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1017),
.A2(n_419),
.B1(n_390),
.B2(n_395),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1141),
.B(n_676),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1036),
.Y(n_1212)
);

NOR2xp67_ASAP7_75t_L g1213 ( 
.A(n_1103),
.B(n_388),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_991),
.A2(n_969),
.B(n_959),
.C(n_543),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1104),
.B(n_544),
.Y(n_1215)
);

AO32x1_ASAP7_75t_L g1216 ( 
.A1(n_992),
.A2(n_547),
.A3(n_545),
.B1(n_544),
.B2(n_498),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1045),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1124),
.A2(n_350),
.B1(n_358),
.B2(n_362),
.Y(n_1218)
);

NOR3xp33_ASAP7_75t_L g1219 ( 
.A(n_1090),
.B(n_416),
.C(n_415),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1036),
.Y(n_1220)
);

NOR2x1_ASAP7_75t_L g1221 ( 
.A(n_1033),
.B(n_676),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1029),
.B(n_698),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1068),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1021),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1065),
.B(n_698),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1127),
.A2(n_747),
.B(n_685),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_989),
.B(n_1094),
.Y(n_1227)
);

O2A1O1Ixp5_ASAP7_75t_L g1228 ( 
.A1(n_1144),
.A2(n_698),
.B(n_762),
.C(n_759),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1127),
.A2(n_789),
.B(n_714),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1080),
.B(n_698),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_1134),
.A2(n_762),
.B(n_759),
.C(n_745),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_R g1232 ( 
.A(n_1100),
.B(n_397),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1052),
.B(n_545),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1154),
.A2(n_789),
.B(n_762),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1154),
.A2(n_789),
.B(n_759),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1116),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1097),
.B(n_364),
.Y(n_1237)
);

NAND3xp33_ASAP7_75t_SL g1238 ( 
.A(n_1134),
.B(n_389),
.C(n_383),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_986),
.A2(n_612),
.B(n_606),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1054),
.B(n_398),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1046),
.B(n_727),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1124),
.A2(n_368),
.B1(n_370),
.B2(n_372),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1003),
.A2(n_789),
.B(n_745),
.Y(n_1243)
);

AOI221x1_ASAP7_75t_L g1244 ( 
.A1(n_1070),
.A2(n_547),
.B1(n_615),
.B2(n_614),
.C(n_612),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1119),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1015),
.A2(n_614),
.B(n_608),
.C(n_611),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1044),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_996),
.B(n_373),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_995),
.A2(n_615),
.B(n_607),
.C(n_608),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1007),
.A2(n_789),
.B(n_745),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1027),
.A2(n_789),
.B(n_745),
.Y(n_1251)
);

NAND2x1p5_ASAP7_75t_L g1252 ( 
.A(n_1150),
.B(n_727),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_973),
.A2(n_727),
.B(n_628),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1036),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1088),
.Y(n_1255)
);

O2A1O1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_979),
.A2(n_607),
.B(n_637),
.C(n_498),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1055),
.A2(n_727),
.B(n_626),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1052),
.B(n_374),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_976),
.A2(n_637),
.B(n_501),
.C(n_503),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1110),
.A2(n_637),
.B(n_501),
.C(n_503),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_1054),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1091),
.Y(n_1262)
);

NOR3xp33_ASAP7_75t_L g1263 ( 
.A(n_994),
.B(n_408),
.C(n_418),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_982),
.A2(n_628),
.B(n_626),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1078),
.B(n_399),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_999),
.A2(n_502),
.B(n_635),
.C(n_631),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_997),
.A2(n_628),
.B(n_743),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1069),
.A2(n_1019),
.B(n_1006),
.C(n_1089),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_998),
.A2(n_628),
.B(n_743),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1158),
.A2(n_412),
.B1(n_261),
.B2(n_252),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1128),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1078),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1130),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1093),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1151),
.B(n_631),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1158),
.A2(n_412),
.B1(n_261),
.B2(n_405),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_R g1277 ( 
.A(n_1135),
.B(n_400),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1002),
.A2(n_743),
.B(n_638),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1145),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_L g1280 ( 
.A(n_1078),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_R g1281 ( 
.A(n_993),
.B(n_379),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1069),
.A2(n_396),
.B1(n_392),
.B2(n_502),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1118),
.B(n_261),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1109),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1160),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1093),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1106),
.A2(n_743),
.B(n_638),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1093),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1131),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1149),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1085),
.A2(n_638),
.B(n_635),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1150),
.B(n_635),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1005),
.B(n_640),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1078),
.B(n_412),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1081),
.B(n_640),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1150),
.B(n_91),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1155),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1023),
.B(n_640),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1081),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1081),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1074),
.A2(n_640),
.B(n_219),
.Y(n_1301)
);

INVx6_ASAP7_75t_L g1302 ( 
.A(n_1081),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1026),
.B(n_640),
.Y(n_1303)
);

INVxp67_ASAP7_75t_L g1304 ( 
.A(n_1146),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1076),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_1093),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1063),
.B(n_993),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1101),
.B(n_640),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1013),
.B(n_640),
.Y(n_1309)
);

NOR3xp33_ASAP7_75t_SL g1310 ( 
.A(n_1016),
.B(n_12),
.C(n_14),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1013),
.B(n_12),
.Y(n_1311)
);

HAxp5_ASAP7_75t_L g1312 ( 
.A(n_1125),
.B(n_14),
.CON(n_1312),
.SN(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1157),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1006),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1028),
.A2(n_1019),
.B(n_1092),
.C(n_1129),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_981),
.A2(n_15),
.B1(n_17),
.B2(n_19),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1098),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1032),
.B(n_20),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1156),
.B(n_212),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1060),
.A2(n_21),
.B(n_24),
.C(n_28),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1126),
.A2(n_206),
.B(n_205),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1050),
.A2(n_21),
.B1(n_29),
.B2(n_32),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1192),
.A2(n_1072),
.B(n_1071),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_1306),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1166),
.A2(n_1011),
.B(n_1101),
.C(n_1062),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1161),
.A2(n_1132),
.B(n_1010),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1199),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_SL g1328 ( 
.A1(n_1188),
.A2(n_1153),
.B(n_1113),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1268),
.A2(n_1037),
.A3(n_1075),
.B(n_1108),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_SL g1330 ( 
.A1(n_1315),
.A2(n_1301),
.B(n_1321),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1201),
.A2(n_1083),
.B(n_1148),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1192),
.A2(n_1253),
.B(n_1264),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1261),
.B(n_1189),
.Y(n_1333)
);

CKINVDCx20_ASAP7_75t_R g1334 ( 
.A(n_1271),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1201),
.A2(n_1117),
.B(n_1120),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1194),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1195),
.Y(n_1337)
);

AO31x2_ASAP7_75t_L g1338 ( 
.A1(n_1244),
.A2(n_1095),
.A3(n_1096),
.B(n_1041),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1165),
.A2(n_1022),
.B(n_1123),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1191),
.A2(n_1038),
.B(n_1012),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1203),
.Y(n_1341)
);

NOR2x1_ASAP7_75t_L g1342 ( 
.A(n_1174),
.B(n_1087),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1177),
.A2(n_1082),
.B(n_1142),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1217),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1168),
.B(n_1032),
.Y(n_1345)
);

NAND2x1p5_ASAP7_75t_L g1346 ( 
.A(n_1174),
.B(n_1156),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1164),
.B(n_1047),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1215),
.B(n_1047),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1301),
.A2(n_1115),
.B(n_1016),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1186),
.B(n_1087),
.Y(n_1350)
);

AOI221xp5_ASAP7_75t_L g1351 ( 
.A1(n_1218),
.A2(n_1152),
.B1(n_1139),
.B2(n_1086),
.C(n_1105),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1183),
.A2(n_1105),
.B(n_1020),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1163),
.B(n_1042),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1193),
.B(n_1042),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1197),
.B(n_1048),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1169),
.A2(n_1048),
.B(n_1137),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1171),
.B(n_1073),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1227),
.A2(n_1098),
.B1(n_1156),
.B2(n_1121),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1308),
.A2(n_1049),
.B(n_1136),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1308),
.A2(n_1049),
.B(n_1147),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1312),
.A2(n_1152),
.B(n_1139),
.C(n_1035),
.Y(n_1361)
);

AOI221xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1322),
.A2(n_1031),
.B1(n_1043),
.B2(n_1051),
.C(n_1059),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1180),
.A2(n_1143),
.B(n_1077),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1305),
.B(n_1098),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1173),
.A2(n_1079),
.B(n_1133),
.Y(n_1365)
);

INVxp67_ASAP7_75t_SL g1366 ( 
.A(n_1289),
.Y(n_1366)
);

A2O1A1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1237),
.A2(n_1030),
.B(n_983),
.C(n_1140),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1189),
.B(n_1098),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1228),
.A2(n_201),
.B(n_197),
.Y(n_1369)
);

NOR4xp25_ASAP7_75t_L g1370 ( 
.A(n_1314),
.B(n_29),
.C(n_32),
.D(n_35),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1205),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1223),
.Y(n_1372)
);

AO31x2_ASAP7_75t_L g1373 ( 
.A1(n_1181),
.A2(n_36),
.A3(n_37),
.B(n_38),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_1182),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1206),
.B(n_36),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1173),
.A2(n_1241),
.B(n_1293),
.Y(n_1376)
);

AND2x6_ASAP7_75t_L g1377 ( 
.A(n_1296),
.B(n_191),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1189),
.B(n_189),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1184),
.B(n_37),
.Y(n_1379)
);

INVx6_ASAP7_75t_L g1380 ( 
.A(n_1167),
.Y(n_1380)
);

AOI221x1_ASAP7_75t_L g1381 ( 
.A1(n_1263),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.C(n_44),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1287),
.A2(n_188),
.B(n_184),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1190),
.A2(n_1239),
.B(n_1298),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1291),
.A2(n_182),
.B(n_178),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1167),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1243),
.A2(n_173),
.B(n_161),
.Y(n_1386)
);

AOI221xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1322),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.C(n_53),
.Y(n_1387)
);

AO31x2_ASAP7_75t_L g1388 ( 
.A1(n_1320),
.A2(n_46),
.A3(n_53),
.B(n_55),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1241),
.A2(n_152),
.B(n_147),
.Y(n_1389)
);

AOI221xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1316),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.C(n_61),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1298),
.A2(n_144),
.B(n_130),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1248),
.B(n_57),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1236),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1250),
.A2(n_129),
.B(n_122),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1257),
.A2(n_107),
.B(n_103),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1175),
.B(n_58),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1257),
.A2(n_1267),
.B(n_1269),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1224),
.B(n_59),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1291),
.A2(n_1303),
.B(n_1200),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_SL g1400 ( 
.A1(n_1316),
.A2(n_61),
.B(n_62),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1234),
.A2(n_62),
.B(n_63),
.Y(n_1401)
);

AOI31xp67_ASAP7_75t_L g1402 ( 
.A1(n_1303),
.A2(n_64),
.A3(n_68),
.B(n_71),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_1270),
.B(n_64),
.C(n_71),
.Y(n_1403)
);

AO31x2_ASAP7_75t_L g1404 ( 
.A1(n_1307),
.A2(n_73),
.A3(n_78),
.B(n_79),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1258),
.B(n_78),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1235),
.A2(n_79),
.B(n_80),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1278),
.A2(n_80),
.B(n_81),
.Y(n_1407)
);

AO31x2_ASAP7_75t_L g1408 ( 
.A1(n_1282),
.A2(n_81),
.A3(n_84),
.B(n_86),
.Y(n_1408)
);

A2O1A1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1219),
.A2(n_84),
.B(n_86),
.C(n_1283),
.Y(n_1409)
);

O2A1O1Ixp5_ASAP7_75t_L g1410 ( 
.A1(n_1294),
.A2(n_1265),
.B(n_1231),
.C(n_1318),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1245),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1170),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1178),
.A2(n_1229),
.B(n_1222),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1178),
.A2(n_1290),
.B1(n_1279),
.B2(n_1273),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1187),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1196),
.Y(n_1416)
);

INVxp33_ASAP7_75t_SL g1417 ( 
.A(n_1277),
.Y(n_1417)
);

AOI21x1_ASAP7_75t_SL g1418 ( 
.A1(n_1296),
.A2(n_1319),
.B(n_1292),
.Y(n_1418)
);

OAI221xp5_ASAP7_75t_L g1419 ( 
.A1(n_1276),
.A2(n_1185),
.B1(n_1172),
.B2(n_1218),
.C(n_1242),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1297),
.B(n_1313),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1242),
.A2(n_1202),
.B(n_1238),
.C(n_1204),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1207),
.Y(n_1422)
);

AOI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1226),
.A2(n_1251),
.B(n_1295),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1233),
.B(n_1204),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1209),
.A2(n_1211),
.B1(n_1304),
.B2(n_1208),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1247),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1202),
.A2(n_1240),
.B(n_1282),
.C(n_1198),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1214),
.A2(n_1210),
.B(n_1311),
.C(n_1213),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1198),
.A2(n_1310),
.B(n_1275),
.C(n_1233),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1221),
.A2(n_1230),
.B(n_1225),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1211),
.A2(n_1256),
.B(n_1285),
.C(n_1284),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1255),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1309),
.A2(n_1292),
.B(n_1319),
.Y(n_1433)
);

AOI221xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1260),
.A2(n_1162),
.B1(n_1246),
.B2(n_1249),
.C(n_1266),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1288),
.A2(n_1252),
.B(n_1216),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1262),
.A2(n_1259),
.B(n_1286),
.C(n_1274),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1300),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1252),
.A2(n_1216),
.B(n_1286),
.Y(n_1438)
);

NOR2xp67_ASAP7_75t_L g1439 ( 
.A(n_1280),
.B(n_1274),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1281),
.B(n_1232),
.Y(n_1440)
);

AO32x2_ASAP7_75t_L g1441 ( 
.A1(n_1216),
.A2(n_1176),
.A3(n_1179),
.B1(n_1317),
.B2(n_1302),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1272),
.A2(n_1299),
.B(n_1212),
.Y(n_1442)
);

AO21x1_ASAP7_75t_L g1443 ( 
.A1(n_1176),
.A2(n_1272),
.B(n_1299),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1272),
.Y(n_1444)
);

AO21x1_ASAP7_75t_L g1445 ( 
.A1(n_1176),
.A2(n_1299),
.B(n_1302),
.Y(n_1445)
);

AND2x6_ASAP7_75t_L g1446 ( 
.A(n_1212),
.B(n_1220),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1176),
.A2(n_1220),
.B(n_1254),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1254),
.A2(n_803),
.B(n_800),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1254),
.A2(n_1166),
.B1(n_1067),
.B2(n_1018),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1212),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1192),
.A2(n_1253),
.B(n_1264),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1168),
.B(n_802),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1271),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1192),
.A2(n_1253),
.B(n_1264),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_SL g1455 ( 
.A1(n_1268),
.A2(n_991),
.B(n_985),
.C(n_801),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1268),
.A2(n_1301),
.B(n_1315),
.Y(n_1456)
);

O2A1O1Ixp5_ASAP7_75t_L g1457 ( 
.A1(n_1301),
.A2(n_1183),
.B(n_1227),
.C(n_1188),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1193),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1161),
.A2(n_803),
.B(n_800),
.Y(n_1459)
);

INVxp67_ASAP7_75t_SL g1460 ( 
.A(n_1289),
.Y(n_1460)
);

AO31x2_ASAP7_75t_L g1461 ( 
.A1(n_1188),
.A2(n_1268),
.A3(n_1244),
.B(n_977),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1192),
.A2(n_1253),
.B(n_1264),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_SL g1463 ( 
.A1(n_1268),
.A2(n_991),
.B(n_985),
.C(n_801),
.Y(n_1463)
);

AOI221x1_ASAP7_75t_L g1464 ( 
.A1(n_1263),
.A2(n_1018),
.B1(n_1301),
.B2(n_916),
.C(n_1268),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1161),
.A2(n_803),
.B(n_800),
.Y(n_1465)
);

INVx6_ASAP7_75t_SL g1466 ( 
.A(n_1233),
.Y(n_1466)
);

NOR2xp67_ASAP7_75t_L g1467 ( 
.A(n_1304),
.B(n_1056),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1192),
.A2(n_1253),
.B(n_1264),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1168),
.B(n_718),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1161),
.A2(n_803),
.B(n_800),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1192),
.A2(n_1253),
.B(n_1264),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_SL g1472 ( 
.A1(n_1268),
.A2(n_991),
.B(n_985),
.C(n_801),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1194),
.Y(n_1473)
);

O2A1O1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1312),
.A2(n_802),
.B(n_1018),
.C(n_916),
.Y(n_1474)
);

A2O1A1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1166),
.A2(n_1227),
.B(n_1237),
.C(n_1301),
.Y(n_1475)
);

AO31x2_ASAP7_75t_L g1476 ( 
.A1(n_1188),
.A2(n_1268),
.A3(n_1244),
.B(n_977),
.Y(n_1476)
);

NAND3xp33_ASAP7_75t_L g1477 ( 
.A(n_1166),
.B(n_1018),
.C(n_802),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1268),
.A2(n_1301),
.B(n_1315),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1192),
.A2(n_1253),
.B(n_1264),
.Y(n_1479)
);

INVxp67_ASAP7_75t_SL g1480 ( 
.A(n_1289),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1161),
.A2(n_803),
.B(n_800),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1194),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1168),
.B(n_802),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1168),
.B(n_802),
.Y(n_1484)
);

OR2x6_ASAP7_75t_L g1485 ( 
.A(n_1189),
.B(n_1280),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1186),
.Y(n_1486)
);

AO21x2_ASAP7_75t_L g1487 ( 
.A1(n_1301),
.A2(n_1268),
.B(n_1177),
.Y(n_1487)
);

AO31x2_ASAP7_75t_L g1488 ( 
.A1(n_1188),
.A2(n_1268),
.A3(n_1244),
.B(n_977),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1168),
.B(n_802),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1268),
.A2(n_1301),
.B(n_1315),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1165),
.A2(n_802),
.B1(n_1040),
.B2(n_1057),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1161),
.A2(n_803),
.B(n_800),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1268),
.A2(n_1301),
.B(n_1315),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_SL g1494 ( 
.A(n_1271),
.B(n_1004),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1419),
.A2(n_1477),
.B1(n_1403),
.B2(n_1405),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1494),
.A2(n_1493),
.B1(n_1456),
.B2(n_1478),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1494),
.A2(n_1493),
.B1(n_1456),
.B2(n_1478),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1477),
.A2(n_1403),
.B1(n_1490),
.B2(n_1392),
.Y(n_1498)
);

BUFx12f_ASAP7_75t_L g1499 ( 
.A(n_1453),
.Y(n_1499)
);

BUFx8_ASAP7_75t_SL g1500 ( 
.A(n_1334),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1490),
.A2(n_1400),
.B1(n_1449),
.B2(n_1491),
.Y(n_1501)
);

INVx6_ASAP7_75t_L g1502 ( 
.A(n_1485),
.Y(n_1502)
);

OAI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1381),
.A2(n_1327),
.B1(n_1486),
.B2(n_1464),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1487),
.A2(n_1330),
.B1(n_1377),
.B2(n_1353),
.Y(n_1504)
);

BUFx12f_ASAP7_75t_L g1505 ( 
.A(n_1385),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1324),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1487),
.A2(n_1377),
.B1(n_1327),
.B2(n_1355),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1475),
.A2(n_1489),
.B1(n_1484),
.B2(n_1483),
.Y(n_1508)
);

CKINVDCx11_ASAP7_75t_R g1509 ( 
.A(n_1485),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1377),
.A2(n_1424),
.B1(n_1357),
.B2(n_1351),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1466),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1377),
.A2(n_1382),
.B1(n_1440),
.B2(n_1390),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1379),
.A2(n_1396),
.B1(n_1382),
.B2(n_1375),
.Y(n_1513)
);

CKINVDCx6p67_ASAP7_75t_R g1514 ( 
.A(n_1485),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1399),
.A2(n_1398),
.B1(n_1374),
.B2(n_1452),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1422),
.Y(n_1516)
);

CKINVDCx11_ASAP7_75t_R g1517 ( 
.A(n_1422),
.Y(n_1517)
);

BUFx8_ASAP7_75t_L g1518 ( 
.A(n_1333),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1390),
.A2(n_1387),
.B1(n_1417),
.B2(n_1366),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1399),
.A2(n_1350),
.B1(n_1482),
.B2(n_1372),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1467),
.A2(n_1333),
.B1(n_1409),
.B2(n_1469),
.Y(n_1521)
);

OAI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1460),
.A2(n_1480),
.B1(n_1347),
.B2(n_1420),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1474),
.A2(n_1421),
.B1(n_1354),
.B2(n_1427),
.Y(n_1523)
);

BUFx4f_ASAP7_75t_L g1524 ( 
.A(n_1380),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1412),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1371),
.Y(n_1526)
);

CKINVDCx6p67_ASAP7_75t_R g1527 ( 
.A(n_1378),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1380),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1345),
.A2(n_1428),
.B1(n_1433),
.B2(n_1458),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1416),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1348),
.A2(n_1344),
.B1(n_1473),
.B2(n_1341),
.Y(n_1531)
);

OAI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1337),
.A2(n_1393),
.B1(n_1411),
.B2(n_1414),
.Y(n_1532)
);

OAI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1364),
.A2(n_1415),
.B1(n_1432),
.B2(n_1387),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1426),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1378),
.A2(n_1425),
.B1(n_1384),
.B2(n_1376),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1466),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1346),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1373),
.Y(n_1538)
);

INVx3_ASAP7_75t_SL g1539 ( 
.A(n_1368),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1384),
.A2(n_1370),
.B1(n_1407),
.B2(n_1352),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1429),
.A2(n_1437),
.B1(n_1325),
.B2(n_1439),
.Y(n_1541)
);

CKINVDCx11_ASAP7_75t_R g1542 ( 
.A(n_1444),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1450),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_SL g1544 ( 
.A(n_1446),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1446),
.Y(n_1545)
);

BUFx12f_ASAP7_75t_L g1546 ( 
.A(n_1346),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1370),
.B(n_1388),
.Y(n_1547)
);

BUFx10_ASAP7_75t_L g1548 ( 
.A(n_1402),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1342),
.Y(n_1549)
);

BUFx2_ASAP7_75t_SL g1550 ( 
.A(n_1445),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1447),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1389),
.A2(n_1407),
.B1(n_1391),
.B2(n_1349),
.Y(n_1552)
);

CKINVDCx6p67_ASAP7_75t_R g1553 ( 
.A(n_1418),
.Y(n_1553)
);

INVx6_ASAP7_75t_L g1554 ( 
.A(n_1443),
.Y(n_1554)
);

INVx4_ASAP7_75t_L g1555 ( 
.A(n_1369),
.Y(n_1555)
);

BUFx2_ASAP7_75t_SL g1556 ( 
.A(n_1442),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1401),
.Y(n_1557)
);

BUFx8_ASAP7_75t_L g1558 ( 
.A(n_1441),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1404),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1358),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1352),
.A2(n_1395),
.B1(n_1369),
.B2(n_1406),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1339),
.A2(n_1356),
.B1(n_1365),
.B2(n_1328),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1326),
.A2(n_1492),
.B(n_1481),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_SL g1564 ( 
.A1(n_1408),
.A2(n_1457),
.B1(n_1455),
.B2(n_1463),
.Y(n_1564)
);

BUFx10_ASAP7_75t_L g1565 ( 
.A(n_1408),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1436),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1410),
.A2(n_1361),
.B(n_1367),
.Y(n_1567)
);

CKINVDCx11_ASAP7_75t_R g1568 ( 
.A(n_1408),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_1438),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1343),
.A2(n_1331),
.B1(n_1413),
.B2(n_1360),
.Y(n_1570)
);

CKINVDCx11_ASAP7_75t_R g1571 ( 
.A(n_1388),
.Y(n_1571)
);

NAND2x1p5_ASAP7_75t_L g1572 ( 
.A(n_1386),
.B(n_1394),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1388),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1359),
.A2(n_1335),
.B1(n_1435),
.B2(n_1397),
.Y(n_1574)
);

INVx6_ASAP7_75t_L g1575 ( 
.A(n_1431),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1441),
.Y(n_1576)
);

CKINVDCx11_ASAP7_75t_R g1577 ( 
.A(n_1472),
.Y(n_1577)
);

CKINVDCx11_ASAP7_75t_R g1578 ( 
.A(n_1434),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1363),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_SL g1580 ( 
.A1(n_1441),
.A2(n_1434),
.B1(n_1479),
.B2(n_1332),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_SL g1581 ( 
.A1(n_1451),
.A2(n_1454),
.B1(n_1471),
.B2(n_1468),
.Y(n_1581)
);

CKINVDCx11_ASAP7_75t_R g1582 ( 
.A(n_1362),
.Y(n_1582)
);

BUFx4_ASAP7_75t_R g1583 ( 
.A(n_1461),
.Y(n_1583)
);

OAI21xp33_ASAP7_75t_L g1584 ( 
.A1(n_1383),
.A2(n_1430),
.B(n_1323),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1462),
.A2(n_1340),
.B1(n_1470),
.B2(n_1465),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1459),
.A2(n_1448),
.B1(n_1476),
.B2(n_1461),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1329),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1476),
.A2(n_1488),
.B1(n_1362),
.B2(n_1329),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1338),
.A2(n_1419),
.B1(n_1477),
.B2(n_1403),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1423),
.A2(n_1475),
.B1(n_1477),
.B2(n_1057),
.Y(n_1590)
);

BUFx8_ASAP7_75t_L g1591 ( 
.A(n_1338),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1338),
.Y(n_1592)
);

INVx6_ASAP7_75t_L g1593 ( 
.A(n_1485),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1494),
.A2(n_735),
.B1(n_1004),
.B2(n_1405),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1422),
.Y(n_1595)
);

INVx4_ASAP7_75t_L g1596 ( 
.A(n_1485),
.Y(n_1596)
);

BUFx8_ASAP7_75t_SL g1597 ( 
.A(n_1334),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1475),
.A2(n_1477),
.B1(n_1057),
.B2(n_802),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1475),
.A2(n_1477),
.B1(n_1057),
.B2(n_802),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1494),
.A2(n_735),
.B1(n_1004),
.B2(n_1405),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1419),
.A2(n_1477),
.B1(n_1403),
.B2(n_1405),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1327),
.B(n_1486),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1327),
.B(n_1486),
.Y(n_1603)
);

BUFx12f_ASAP7_75t_L g1604 ( 
.A(n_1453),
.Y(n_1604)
);

BUFx12f_ASAP7_75t_L g1605 ( 
.A(n_1453),
.Y(n_1605)
);

BUFx10_ASAP7_75t_L g1606 ( 
.A(n_1453),
.Y(n_1606)
);

INVx4_ASAP7_75t_L g1607 ( 
.A(n_1485),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1324),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1336),
.Y(n_1609)
);

INVx6_ASAP7_75t_L g1610 ( 
.A(n_1485),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1419),
.A2(n_1477),
.B1(n_1403),
.B2(n_1405),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1419),
.A2(n_1477),
.B1(n_1403),
.B2(n_1405),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1336),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1446),
.Y(n_1614)
);

INVx3_ASAP7_75t_SL g1615 ( 
.A(n_1453),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1336),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_1446),
.Y(n_1617)
);

INVx8_ASAP7_75t_L g1618 ( 
.A(n_1446),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1419),
.A2(n_1477),
.B1(n_1403),
.B2(n_1405),
.Y(n_1619)
);

NAND2x1p5_ASAP7_75t_L g1620 ( 
.A(n_1447),
.B(n_1066),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1453),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1336),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1422),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1419),
.A2(n_1477),
.B1(n_1403),
.B2(n_1405),
.Y(n_1624)
);

CKINVDCx11_ASAP7_75t_R g1625 ( 
.A(n_1324),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1494),
.A2(n_735),
.B1(n_1004),
.B2(n_1405),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1336),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1336),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1446),
.Y(n_1629)
);

CKINVDCx10_ASAP7_75t_R g1630 ( 
.A(n_1485),
.Y(n_1630)
);

NAND2x1p5_ASAP7_75t_L g1631 ( 
.A(n_1447),
.B(n_1066),
.Y(n_1631)
);

CKINVDCx6p67_ASAP7_75t_R g1632 ( 
.A(n_1485),
.Y(n_1632)
);

BUFx2_ASAP7_75t_SL g1633 ( 
.A(n_1324),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1422),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1334),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1475),
.A2(n_1477),
.B1(n_1057),
.B2(n_802),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1336),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1324),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1336),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1422),
.Y(n_1640)
);

INVx8_ASAP7_75t_L g1641 ( 
.A(n_1446),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1324),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1419),
.A2(n_1477),
.B1(n_1403),
.B2(n_1405),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1419),
.A2(n_1477),
.B1(n_1403),
.B2(n_1405),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1475),
.A2(n_1477),
.B1(n_1057),
.B2(n_802),
.Y(n_1645)
);

NAND2x1p5_ASAP7_75t_L g1646 ( 
.A(n_1447),
.B(n_1066),
.Y(n_1646)
);

INVx5_ASAP7_75t_L g1647 ( 
.A(n_1446),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1419),
.A2(n_1477),
.B1(n_1403),
.B2(n_1405),
.Y(n_1648)
);

OAI22x1_ASAP7_75t_SL g1649 ( 
.A1(n_1417),
.A2(n_1385),
.B1(n_575),
.B2(n_1271),
.Y(n_1649)
);

BUFx8_ASAP7_75t_L g1650 ( 
.A(n_1440),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1336),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1475),
.A2(n_1478),
.B(n_1456),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1446),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1587),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1551),
.B(n_1579),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1516),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1559),
.Y(n_1657)
);

INVx4_ASAP7_75t_L g1658 ( 
.A(n_1647),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1573),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1538),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1567),
.B(n_1652),
.Y(n_1661)
);

INVx5_ASAP7_75t_L g1662 ( 
.A(n_1575),
.Y(n_1662)
);

O2A1O1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1598),
.A2(n_1599),
.B(n_1636),
.C(n_1645),
.Y(n_1663)
);

OAI21x1_ASAP7_75t_L g1664 ( 
.A1(n_1563),
.A2(n_1572),
.B(n_1585),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1547),
.B(n_1496),
.Y(n_1665)
);

BUFx2_ASAP7_75t_L g1666 ( 
.A(n_1591),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1508),
.B(n_1515),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1496),
.B(n_1497),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1565),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1592),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1495),
.A2(n_1611),
.B(n_1601),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1565),
.Y(n_1672)
);

AO21x2_ASAP7_75t_L g1673 ( 
.A1(n_1584),
.A2(n_1533),
.B(n_1557),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1595),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1497),
.B(n_1576),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_1554),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1623),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1576),
.B(n_1582),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1591),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1634),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1555),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1640),
.Y(n_1682)
);

AOI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1590),
.A2(n_1523),
.B(n_1541),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1613),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1502),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1576),
.B(n_1589),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1576),
.B(n_1589),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1502),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1572),
.A2(n_1585),
.B(n_1574),
.Y(n_1689)
);

OAI21x1_ASAP7_75t_L g1690 ( 
.A1(n_1574),
.A2(n_1570),
.B(n_1562),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1588),
.B(n_1504),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1583),
.Y(n_1692)
);

BUFx3_ASAP7_75t_L g1693 ( 
.A(n_1502),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1602),
.Y(n_1694)
);

AO21x2_ASAP7_75t_L g1695 ( 
.A1(n_1533),
.A2(n_1532),
.B(n_1503),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1588),
.B(n_1504),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1593),
.Y(n_1697)
);

INVx4_ASAP7_75t_L g1698 ( 
.A(n_1647),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1569),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1548),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1532),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1548),
.Y(n_1702)
);

OA21x2_ASAP7_75t_L g1703 ( 
.A1(n_1570),
.A2(n_1562),
.B(n_1586),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1616),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1580),
.B(n_1498),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1622),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1552),
.A2(n_1586),
.B(n_1631),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1628),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1517),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1495),
.A2(n_1619),
.B1(n_1648),
.B2(n_1644),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1637),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1515),
.B(n_1601),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1651),
.Y(n_1713)
);

BUFx12f_ASAP7_75t_L g1714 ( 
.A(n_1625),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1575),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1593),
.Y(n_1716)
);

AO21x2_ASAP7_75t_L g1717 ( 
.A1(n_1503),
.A2(n_1529),
.B(n_1522),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1558),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1575),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1520),
.B(n_1522),
.Y(n_1720)
);

NAND2x1p5_ASAP7_75t_L g1721 ( 
.A(n_1566),
.B(n_1647),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_SL g1722 ( 
.A1(n_1558),
.A2(n_1566),
.B1(n_1593),
.B2(n_1610),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1564),
.Y(n_1723)
);

BUFx3_ASAP7_75t_L g1724 ( 
.A(n_1610),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1552),
.A2(n_1535),
.B(n_1510),
.Y(n_1725)
);

OAI21x1_ASAP7_75t_L g1726 ( 
.A1(n_1620),
.A2(n_1646),
.B(n_1631),
.Y(n_1726)
);

AOI21x1_ASAP7_75t_L g1727 ( 
.A1(n_1531),
.A2(n_1549),
.B(n_1545),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1554),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1580),
.B(n_1498),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1620),
.Y(n_1730)
);

OA21x2_ASAP7_75t_L g1731 ( 
.A1(n_1535),
.A2(n_1520),
.B(n_1510),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_1577),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1564),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1609),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1610),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1627),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1646),
.A2(n_1507),
.B(n_1501),
.Y(n_1737)
);

OA21x2_ASAP7_75t_L g1738 ( 
.A1(n_1507),
.A2(n_1501),
.B(n_1648),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1639),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1611),
.A2(n_1612),
.B1(n_1619),
.B2(n_1643),
.Y(n_1740)
);

BUFx2_ASAP7_75t_SL g1741 ( 
.A(n_1647),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1596),
.B(n_1607),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1560),
.B(n_1603),
.Y(n_1743)
);

AOI21x1_ASAP7_75t_L g1744 ( 
.A1(n_1534),
.A2(n_1530),
.B(n_1525),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1612),
.B(n_1624),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1571),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1539),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1568),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1550),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1578),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_L g1751 ( 
.A(n_1624),
.B(n_1643),
.C(n_1644),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1556),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1581),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1539),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1581),
.Y(n_1755)
);

BUFx12f_ASAP7_75t_L g1756 ( 
.A(n_1509),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1594),
.A2(n_1600),
.B1(n_1626),
.B2(n_1521),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1540),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1540),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1543),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1561),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1618),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1537),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1561),
.Y(n_1764)
);

NAND2x1_ASAP7_75t_L g1765 ( 
.A(n_1614),
.B(n_1653),
.Y(n_1765)
);

OAI21x1_ASAP7_75t_L g1766 ( 
.A1(n_1513),
.A2(n_1553),
.B(n_1544),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1513),
.B(n_1519),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1512),
.B(n_1519),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1512),
.Y(n_1769)
);

OAI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1594),
.A2(n_1600),
.B(n_1626),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1544),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1607),
.B(n_1653),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1617),
.Y(n_1773)
);

BUFx4f_ASAP7_75t_SL g1774 ( 
.A(n_1635),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1506),
.B(n_1608),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1617),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1629),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_SL g1778 ( 
.A1(n_1633),
.A2(n_1518),
.B1(n_1641),
.B2(n_1638),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1694),
.B(n_1642),
.Y(n_1779)
);

AO32x2_ASAP7_75t_L g1780 ( 
.A1(n_1757),
.A2(n_1632),
.A3(n_1514),
.B1(n_1542),
.B2(n_1630),
.Y(n_1780)
);

OAI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1751),
.A2(n_1536),
.B(n_1524),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1661),
.B(n_1527),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1661),
.B(n_1518),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1725),
.A2(n_1641),
.B(n_1629),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1661),
.B(n_1653),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1660),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1743),
.B(n_1615),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1693),
.B(n_1511),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1710),
.A2(n_1649),
.B1(n_1650),
.B2(n_1615),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1678),
.B(n_1748),
.Y(n_1790)
);

INVxp33_ASAP7_75t_L g1791 ( 
.A(n_1656),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1697),
.B(n_1528),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1678),
.B(n_1606),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1748),
.B(n_1606),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1743),
.B(n_1526),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1748),
.B(n_1524),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1675),
.B(n_1621),
.Y(n_1797)
);

A2O1A1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1671),
.A2(n_1546),
.B(n_1650),
.C(n_1597),
.Y(n_1798)
);

NOR2x1_ASAP7_75t_SL g1799 ( 
.A(n_1662),
.B(n_1499),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1697),
.B(n_1505),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1659),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1740),
.A2(n_1604),
.B1(n_1605),
.B2(n_1500),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1774),
.Y(n_1803)
);

INVx5_ASAP7_75t_L g1804 ( 
.A(n_1662),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1745),
.B(n_1663),
.Y(n_1805)
);

O2A1O1Ixp33_ASAP7_75t_SL g1806 ( 
.A1(n_1750),
.A2(n_1770),
.B(n_1712),
.C(n_1767),
.Y(n_1806)
);

O2A1O1Ixp33_ASAP7_75t_SL g1807 ( 
.A1(n_1750),
.A2(n_1767),
.B(n_1667),
.C(n_1765),
.Y(n_1807)
);

NOR2x1_ASAP7_75t_SL g1808 ( 
.A(n_1662),
.B(n_1717),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1668),
.A2(n_1750),
.B1(n_1768),
.B2(n_1662),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1697),
.B(n_1724),
.Y(n_1810)
);

AO32x2_ASAP7_75t_L g1811 ( 
.A1(n_1685),
.A2(n_1716),
.A3(n_1688),
.B1(n_1698),
.B2(n_1658),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1746),
.B(n_1665),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_1714),
.Y(n_1813)
);

OAI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1668),
.A2(n_1768),
.B1(n_1662),
.B2(n_1769),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1661),
.B(n_1701),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1692),
.B(n_1718),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1657),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1714),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1718),
.B(n_1686),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1724),
.B(n_1735),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1699),
.B(n_1686),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1662),
.A2(n_1720),
.B1(n_1732),
.B2(n_1738),
.Y(n_1822)
);

OA21x2_ASAP7_75t_L g1823 ( 
.A1(n_1707),
.A2(n_1689),
.B(n_1690),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1687),
.B(n_1655),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1687),
.B(n_1655),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1683),
.B(n_1720),
.Y(n_1826)
);

OA21x2_ASAP7_75t_L g1827 ( 
.A1(n_1707),
.A2(n_1737),
.B(n_1664),
.Y(n_1827)
);

AOI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1717),
.A2(n_1705),
.B1(n_1729),
.B2(n_1701),
.C(n_1695),
.Y(n_1828)
);

INVxp67_ASAP7_75t_L g1829 ( 
.A(n_1749),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1735),
.B(n_1679),
.Y(n_1830)
);

A2O1A1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1705),
.A2(n_1729),
.B(n_1737),
.C(n_1766),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1747),
.Y(n_1832)
);

AO32x2_ASAP7_75t_L g1833 ( 
.A1(n_1685),
.A2(n_1716),
.A3(n_1688),
.B1(n_1698),
.B2(n_1658),
.Y(n_1833)
);

NOR2x1_ASAP7_75t_L g1834 ( 
.A(n_1752),
.B(n_1749),
.Y(n_1834)
);

OAI21x1_ASAP7_75t_L g1835 ( 
.A1(n_1726),
.A2(n_1744),
.B(n_1683),
.Y(n_1835)
);

A2O1A1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1766),
.A2(n_1733),
.B(n_1723),
.C(n_1719),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1666),
.B(n_1674),
.Y(n_1837)
);

INVx2_ASAP7_75t_SL g1838 ( 
.A(n_1756),
.Y(n_1838)
);

NOR2x1_ASAP7_75t_SL g1839 ( 
.A(n_1727),
.B(n_1741),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1758),
.B(n_1759),
.Y(n_1840)
);

BUFx3_ASAP7_75t_L g1841 ( 
.A(n_1756),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1719),
.B(n_1715),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1742),
.B(n_1730),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1677),
.B(n_1680),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1682),
.B(n_1763),
.Y(n_1845)
);

A2O1A1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1723),
.A2(n_1733),
.B(n_1715),
.C(n_1759),
.Y(n_1846)
);

AND2x4_ASAP7_75t_SL g1847 ( 
.A(n_1732),
.B(n_1762),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1704),
.B(n_1706),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1684),
.B(n_1704),
.Y(n_1849)
);

AO21x1_ASAP7_75t_L g1850 ( 
.A1(n_1721),
.A2(n_1773),
.B(n_1776),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1732),
.A2(n_1738),
.B1(n_1722),
.B2(n_1715),
.Y(n_1851)
);

NOR3xp33_ASAP7_75t_SL g1852 ( 
.A(n_1775),
.B(n_1702),
.C(n_1672),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1754),
.B(n_1728),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1738),
.A2(n_1731),
.B1(n_1778),
.B2(n_1695),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1742),
.B(n_1730),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1823),
.B(n_1753),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1786),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1815),
.B(n_1761),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1815),
.B(n_1761),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1823),
.B(n_1753),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1786),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1812),
.B(n_1755),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1824),
.B(n_1764),
.Y(n_1863)
);

INVx4_ASAP7_75t_L g1864 ( 
.A(n_1804),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1827),
.B(n_1764),
.Y(n_1865)
);

INVx1_ASAP7_75t_SL g1866 ( 
.A(n_1832),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1801),
.Y(n_1867)
);

NOR2x1_ASAP7_75t_L g1868 ( 
.A(n_1834),
.B(n_1695),
.Y(n_1868)
);

NOR2xp67_ASAP7_75t_L g1869 ( 
.A(n_1804),
.B(n_1702),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1828),
.B(n_1691),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1805),
.A2(n_1731),
.B1(n_1691),
.B2(n_1696),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1817),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1825),
.B(n_1696),
.Y(n_1873)
);

NOR3xp33_ASAP7_75t_L g1874 ( 
.A(n_1805),
.B(n_1728),
.C(n_1752),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1827),
.B(n_1703),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1831),
.B(n_1703),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1828),
.B(n_1670),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1829),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1831),
.B(n_1703),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1848),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1848),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1806),
.A2(n_1731),
.B1(n_1732),
.B2(n_1771),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1809),
.A2(n_1771),
.B1(n_1676),
.B2(n_1742),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1849),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1821),
.B(n_1681),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1826),
.B(n_1670),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1826),
.B(n_1840),
.Y(n_1887)
);

AOI21xp33_ASAP7_75t_L g1888 ( 
.A1(n_1854),
.A2(n_1752),
.B(n_1700),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1811),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1819),
.B(n_1681),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1811),
.B(n_1654),
.Y(n_1891)
);

INVxp67_ASAP7_75t_L g1892 ( 
.A(n_1853),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1811),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1816),
.B(n_1669),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1811),
.B(n_1669),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1808),
.B(n_1673),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1845),
.B(n_1846),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1822),
.B(n_1673),
.Y(n_1898)
);

INVx2_ASAP7_75t_SL g1899 ( 
.A(n_1878),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1892),
.B(n_1844),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1870),
.A2(n_1809),
.B1(n_1851),
.B2(n_1822),
.Y(n_1901)
);

OAI211xp5_ASAP7_75t_L g1902 ( 
.A1(n_1870),
.A2(n_1806),
.B(n_1836),
.C(n_1781),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1891),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1858),
.B(n_1791),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1891),
.Y(n_1905)
);

OAI221xp5_ASAP7_75t_L g1906 ( 
.A1(n_1871),
.A2(n_1789),
.B1(n_1802),
.B2(n_1781),
.C(n_1798),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1878),
.Y(n_1907)
);

OAI211xp5_ASAP7_75t_L g1908 ( 
.A1(n_1882),
.A2(n_1836),
.B(n_1846),
.C(n_1807),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1857),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1882),
.A2(n_1852),
.B(n_1807),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1873),
.B(n_1790),
.Y(n_1911)
);

INVxp67_ASAP7_75t_SL g1912 ( 
.A(n_1868),
.Y(n_1912)
);

AOI211xp5_ASAP7_75t_L g1913 ( 
.A1(n_1888),
.A2(n_1802),
.B(n_1798),
.C(n_1851),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1891),
.B(n_1843),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1873),
.B(n_1837),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1867),
.Y(n_1916)
);

BUFx3_ASAP7_75t_L g1917 ( 
.A(n_1866),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1863),
.B(n_1833),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1863),
.B(n_1833),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1858),
.B(n_1791),
.Y(n_1920)
);

INVx3_ASAP7_75t_L g1921 ( 
.A(n_1864),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1892),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1890),
.B(n_1833),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1887),
.B(n_1853),
.Y(n_1924)
);

NAND3xp33_ASAP7_75t_L g1925 ( 
.A(n_1868),
.B(n_1852),
.C(n_1814),
.Y(n_1925)
);

OAI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1883),
.A2(n_1784),
.B1(n_1721),
.B2(n_1783),
.Y(n_1926)
);

AOI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1876),
.A2(n_1814),
.B1(n_1879),
.B2(n_1784),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1867),
.Y(n_1928)
);

OAI211xp5_ASAP7_75t_L g1929 ( 
.A1(n_1877),
.A2(n_1842),
.B(n_1783),
.C(n_1760),
.Y(n_1929)
);

INVx4_ASAP7_75t_L g1930 ( 
.A(n_1864),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1859),
.B(n_1779),
.Y(n_1931)
);

BUFx2_ASAP7_75t_L g1932 ( 
.A(n_1889),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1857),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1866),
.A2(n_1721),
.B1(n_1732),
.B2(n_1782),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1861),
.Y(n_1935)
);

AOI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1876),
.A2(n_1782),
.B1(n_1787),
.B2(n_1794),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1890),
.B(n_1839),
.Y(n_1937)
);

AOI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1876),
.A2(n_1830),
.B1(n_1785),
.B2(n_1788),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1862),
.B(n_1797),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1879),
.A2(n_1830),
.B1(n_1785),
.B2(n_1788),
.Y(n_1940)
);

AO21x2_ASAP7_75t_L g1941 ( 
.A1(n_1896),
.A2(n_1850),
.B(n_1835),
.Y(n_1941)
);

AOI221xp5_ASAP7_75t_L g1942 ( 
.A1(n_1879),
.A2(n_1842),
.B1(n_1711),
.B2(n_1713),
.C(n_1708),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1859),
.B(n_1673),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1887),
.B(n_1672),
.Y(n_1944)
);

OR2x6_ASAP7_75t_L g1945 ( 
.A(n_1864),
.B(n_1898),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1862),
.B(n_1855),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1864),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1874),
.A2(n_1838),
.B1(n_1810),
.B2(n_1820),
.Y(n_1948)
);

OAI221xp5_ASAP7_75t_L g1949 ( 
.A1(n_1877),
.A2(n_1709),
.B1(n_1795),
.B2(n_1818),
.C(n_1841),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1897),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1897),
.B(n_1885),
.Y(n_1951)
);

OAI33xp33_ASAP7_75t_L g1952 ( 
.A1(n_1886),
.A2(n_1713),
.A3(n_1736),
.B1(n_1739),
.B2(n_1734),
.B3(n_1773),
.Y(n_1952)
);

XOR2xp5_ASAP7_75t_L g1953 ( 
.A(n_1894),
.B(n_1813),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1872),
.Y(n_1954)
);

INVxp67_ASAP7_75t_L g1955 ( 
.A(n_1884),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1872),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1950),
.B(n_1880),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1903),
.B(n_1889),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1907),
.Y(n_1959)
);

NOR2xp67_ASAP7_75t_L g1960 ( 
.A(n_1925),
.B(n_1893),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1903),
.B(n_1893),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1916),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1949),
.B(n_1796),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1932),
.B(n_1898),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1905),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1916),
.Y(n_1966)
);

NOR3xp33_ASAP7_75t_L g1967 ( 
.A(n_1906),
.B(n_1902),
.C(n_1908),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1928),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1899),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1928),
.Y(n_1970)
);

AND2x2_ASAP7_75t_SL g1971 ( 
.A(n_1901),
.B(n_1874),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1918),
.B(n_1896),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1925),
.A2(n_1910),
.B1(n_1927),
.B2(n_1888),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_SL g1974 ( 
.A(n_1910),
.B(n_1804),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1954),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1913),
.B(n_1804),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1918),
.B(n_1875),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1954),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1932),
.B(n_1865),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1921),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1919),
.B(n_1875),
.Y(n_1981)
);

INVx1_ASAP7_75t_SL g1982 ( 
.A(n_1941),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1921),
.B(n_1869),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1919),
.B(n_1875),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1921),
.B(n_1869),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1955),
.B(n_1881),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1956),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1909),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1941),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1923),
.B(n_1895),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1943),
.B(n_1865),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1941),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1923),
.B(n_1895),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1909),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1914),
.B(n_1856),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1914),
.B(n_1856),
.Y(n_1996)
);

NOR2xp67_ASAP7_75t_L g1997 ( 
.A(n_1927),
.B(n_1856),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1933),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1914),
.B(n_1860),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1933),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1914),
.B(n_1860),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1922),
.B(n_1881),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1899),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1935),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1945),
.B(n_1860),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1964),
.B(n_1943),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1988),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1988),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1964),
.B(n_1944),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1961),
.Y(n_2010)
);

AND2x4_ASAP7_75t_L g2011 ( 
.A(n_1983),
.B(n_1945),
.Y(n_2011)
);

OAI22xp5_ASAP7_75t_L g2012 ( 
.A1(n_1973),
.A2(n_1913),
.B1(n_1953),
.B2(n_1948),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1971),
.B(n_1911),
.Y(n_2013)
);

INVx1_ASAP7_75t_SL g2014 ( 
.A(n_1976),
.Y(n_2014)
);

INVx3_ASAP7_75t_L g2015 ( 
.A(n_1980),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1988),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1994),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1957),
.B(n_1951),
.Y(n_2018)
);

AOI21xp33_ASAP7_75t_L g2019 ( 
.A1(n_1973),
.A2(n_1929),
.B(n_1934),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1997),
.B(n_1937),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1971),
.B(n_1911),
.Y(n_2021)
);

AO22x1_ASAP7_75t_L g2022 ( 
.A1(n_1967),
.A2(n_1917),
.B1(n_1912),
.B2(n_1793),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1994),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1994),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2000),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1957),
.B(n_1904),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1997),
.B(n_1937),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1964),
.B(n_1944),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2000),
.Y(n_2029)
);

OAI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_1971),
.A2(n_1953),
.B1(n_1938),
.B2(n_1940),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1967),
.B(n_1931),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1971),
.B(n_1915),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2000),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1997),
.B(n_1945),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1961),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2004),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1961),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1971),
.B(n_1915),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1963),
.B(n_1939),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1990),
.B(n_1945),
.Y(n_2040)
);

OAI21xp33_ASAP7_75t_L g2041 ( 
.A1(n_1976),
.A2(n_1936),
.B(n_1945),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2004),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2004),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1963),
.B(n_1939),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1998),
.Y(n_2045)
);

OR2x2_ASAP7_75t_L g2046 ( 
.A(n_1964),
.B(n_1904),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1998),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1961),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1998),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1974),
.B(n_1917),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1990),
.B(n_1946),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_1991),
.B(n_1920),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1998),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_1991),
.B(n_1920),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1990),
.B(n_1946),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1986),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_2031),
.B(n_2014),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2007),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2008),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2015),
.Y(n_2060)
);

OAI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_2012),
.A2(n_1974),
.B1(n_1960),
.B2(n_1732),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_2013),
.B(n_1931),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2016),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2051),
.B(n_1995),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_2051),
.B(n_1960),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2017),
.Y(n_2066)
);

INVx2_ASAP7_75t_SL g2067 ( 
.A(n_2011),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2023),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2031),
.B(n_1960),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_SL g2070 ( 
.A(n_2019),
.B(n_1974),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_2021),
.B(n_1924),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2024),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2039),
.B(n_2002),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2025),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2055),
.B(n_2040),
.Y(n_2075)
);

AOI22xp5_ASAP7_75t_L g2076 ( 
.A1(n_2030),
.A2(n_1926),
.B1(n_2005),
.B2(n_1952),
.Y(n_2076)
);

AOI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_2041),
.A2(n_2005),
.B1(n_1983),
.B2(n_1985),
.Y(n_2077)
);

INVx3_ASAP7_75t_SL g2078 ( 
.A(n_2050),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2044),
.B(n_2002),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2055),
.B(n_1995),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2040),
.B(n_1995),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2029),
.Y(n_2082)
);

INVxp67_ASAP7_75t_L g2083 ( 
.A(n_2032),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_2038),
.B(n_1959),
.Y(n_2084)
);

OR2x6_ASAP7_75t_L g2085 ( 
.A(n_2050),
.B(n_1741),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2033),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2036),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2034),
.B(n_2005),
.Y(n_2088)
);

NOR2x1_ASAP7_75t_L g2089 ( 
.A(n_2034),
.B(n_1980),
.Y(n_2089)
);

NAND2x1p5_ASAP7_75t_L g2090 ( 
.A(n_2011),
.B(n_1930),
.Y(n_2090)
);

OR2x2_ASAP7_75t_L g2091 ( 
.A(n_2018),
.B(n_1959),
.Y(n_2091)
);

OAI21xp33_ASAP7_75t_L g2092 ( 
.A1(n_2056),
.A2(n_2005),
.B(n_1991),
.Y(n_2092)
);

NOR4xp75_ASAP7_75t_L g2093 ( 
.A(n_2020),
.B(n_2027),
.C(n_2015),
.D(n_1980),
.Y(n_2093)
);

INVxp33_ASAP7_75t_L g2094 ( 
.A(n_2046),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2042),
.Y(n_2095)
);

NOR3xp33_ASAP7_75t_L g2096 ( 
.A(n_2022),
.B(n_1982),
.C(n_1989),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2065),
.Y(n_2097)
);

OAI221xp5_ASAP7_75t_L g2098 ( 
.A1(n_2070),
.A2(n_2046),
.B1(n_2026),
.B2(n_2052),
.C(n_2054),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_2057),
.B(n_1803),
.Y(n_2099)
);

INVx2_ASAP7_75t_SL g2100 ( 
.A(n_2089),
.Y(n_2100)
);

AOI21xp5_ASAP7_75t_L g2101 ( 
.A1(n_2070),
.A2(n_1982),
.B(n_2011),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2069),
.B(n_2020),
.Y(n_2102)
);

INVxp67_ASAP7_75t_L g2103 ( 
.A(n_2067),
.Y(n_2103)
);

OAI32xp33_ASAP7_75t_L g2104 ( 
.A1(n_2096),
.A2(n_1982),
.A3(n_1979),
.B1(n_1992),
.B2(n_1989),
.Y(n_2104)
);

INVx2_ASAP7_75t_SL g2105 ( 
.A(n_2090),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2078),
.B(n_2027),
.Y(n_2106)
);

OAI21xp33_ASAP7_75t_L g2107 ( 
.A1(n_2076),
.A2(n_1992),
.B(n_1989),
.Y(n_2107)
);

AOI32xp33_ASAP7_75t_L g2108 ( 
.A1(n_2061),
.A2(n_2096),
.A3(n_2094),
.B1(n_2065),
.B2(n_2078),
.Y(n_2108)
);

INVxp67_ASAP7_75t_L g2109 ( 
.A(n_2067),
.Y(n_2109)
);

AOI321xp33_ASAP7_75t_L g2110 ( 
.A1(n_2061),
.A2(n_1989),
.A3(n_1992),
.B1(n_2054),
.B2(n_2052),
.C(n_2006),
.Y(n_2110)
);

OAI21xp5_ASAP7_75t_SL g2111 ( 
.A1(n_2077),
.A2(n_1800),
.B(n_1847),
.Y(n_2111)
);

OAI31xp33_ASAP7_75t_L g2112 ( 
.A1(n_2094),
.A2(n_2028),
.A3(n_2009),
.B(n_1985),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2075),
.B(n_1995),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2083),
.B(n_2009),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2085),
.B(n_1996),
.Y(n_2115)
);

O2A1O1Ixp33_ASAP7_75t_L g2116 ( 
.A1(n_2083),
.A2(n_1992),
.B(n_2028),
.C(n_1979),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2071),
.B(n_1990),
.Y(n_2117)
);

AOI222xp33_ASAP7_75t_L g2118 ( 
.A1(n_2092),
.A2(n_1942),
.B1(n_1865),
.B2(n_1993),
.C1(n_1972),
.C2(n_1981),
.Y(n_2118)
);

OA21x2_ASAP7_75t_L g2119 ( 
.A1(n_2060),
.A2(n_2059),
.B(n_2058),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2063),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2088),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2085),
.B(n_1996),
.Y(n_2122)
);

AOI21xp33_ASAP7_75t_L g2123 ( 
.A1(n_2085),
.A2(n_2006),
.B(n_2043),
.Y(n_2123)
);

INVxp67_ASAP7_75t_SL g2124 ( 
.A(n_2090),
.Y(n_2124)
);

AOI322xp5_ASAP7_75t_L g2125 ( 
.A1(n_2073),
.A2(n_1993),
.A3(n_1981),
.B1(n_1977),
.B2(n_1984),
.C1(n_1972),
.C2(n_1958),
.Y(n_2125)
);

AND2x4_ASAP7_75t_L g2126 ( 
.A(n_2100),
.B(n_2093),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_2107),
.A2(n_2079),
.B(n_2084),
.Y(n_2127)
);

OAI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_2107),
.A2(n_2091),
.B(n_2062),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2120),
.Y(n_2129)
);

AOI321xp33_ASAP7_75t_SL g2130 ( 
.A1(n_2110),
.A2(n_2088),
.A3(n_2095),
.B1(n_2087),
.B2(n_2086),
.C(n_2082),
.Y(n_2130)
);

OAI22xp33_ASAP7_75t_L g2131 ( 
.A1(n_2098),
.A2(n_1979),
.B1(n_1780),
.B2(n_2003),
.Y(n_2131)
);

AOI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_2108),
.A2(n_2068),
.B(n_2066),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2103),
.B(n_2064),
.Y(n_2133)
);

OAI21xp5_ASAP7_75t_L g2134 ( 
.A1(n_2101),
.A2(n_2074),
.B(n_2072),
.Y(n_2134)
);

AOI21xp33_ASAP7_75t_L g2135 ( 
.A1(n_2108),
.A2(n_2060),
.B(n_2081),
.Y(n_2135)
);

OAI21xp33_ASAP7_75t_L g2136 ( 
.A1(n_2102),
.A2(n_2080),
.B(n_2047),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2106),
.B(n_1996),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_2112),
.B(n_1983),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2109),
.B(n_1993),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2120),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2119),
.Y(n_2141)
);

AOI221xp5_ASAP7_75t_L g2142 ( 
.A1(n_2104),
.A2(n_2053),
.B1(n_2049),
.B2(n_2045),
.C(n_2015),
.Y(n_2142)
);

AOI21xp5_ASAP7_75t_SL g2143 ( 
.A1(n_2124),
.A2(n_1800),
.B(n_1983),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2106),
.B(n_1996),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2097),
.B(n_2121),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_2100),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2097),
.B(n_1993),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2121),
.B(n_1999),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2099),
.B(n_1999),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2146),
.B(n_2114),
.Y(n_2150)
);

HAxp5_ASAP7_75t_SL g2151 ( 
.A(n_2130),
.B(n_2111),
.CON(n_2151),
.SN(n_2151)
);

INVxp33_ASAP7_75t_L g2152 ( 
.A(n_2133),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2146),
.B(n_2105),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2132),
.B(n_2105),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2145),
.B(n_2113),
.Y(n_2155)
);

XOR2x2_ASAP7_75t_L g2156 ( 
.A(n_2149),
.B(n_1792),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2141),
.Y(n_2157)
);

OR2x2_ASAP7_75t_L g2158 ( 
.A(n_2139),
.B(n_2117),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2129),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2137),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2140),
.B(n_2125),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2147),
.Y(n_2162)
);

OAI221xp5_ASAP7_75t_L g2163 ( 
.A1(n_2128),
.A2(n_2123),
.B1(n_2118),
.B2(n_2116),
.C(n_2122),
.Y(n_2163)
);

A2O1A1Ixp33_ASAP7_75t_L g2164 ( 
.A1(n_2127),
.A2(n_2104),
.B(n_2122),
.C(n_2115),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2160),
.B(n_2144),
.Y(n_2165)
);

NAND3xp33_ASAP7_75t_SL g2166 ( 
.A(n_2164),
.B(n_2134),
.C(n_2138),
.Y(n_2166)
);

AOI211xp5_ASAP7_75t_L g2167 ( 
.A1(n_2163),
.A2(n_2131),
.B(n_2154),
.C(n_2135),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2157),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2156),
.Y(n_2169)
);

HB1xp67_ASAP7_75t_L g2170 ( 
.A(n_2153),
.Y(n_2170)
);

OAI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_2161),
.A2(n_2131),
.B1(n_2152),
.B2(n_2126),
.Y(n_2171)
);

NOR3x1_ASAP7_75t_L g2172 ( 
.A(n_2150),
.B(n_2138),
.C(n_2148),
.Y(n_2172)
);

HB1xp67_ASAP7_75t_L g2173 ( 
.A(n_2150),
.Y(n_2173)
);

AOI211xp5_ASAP7_75t_SL g2174 ( 
.A1(n_2161),
.A2(n_2143),
.B(n_2151),
.C(n_2159),
.Y(n_2174)
);

NAND3xp33_ASAP7_75t_L g2175 ( 
.A(n_2162),
.B(n_2126),
.C(n_2136),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_2155),
.B(n_2126),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2170),
.B(n_2158),
.Y(n_2177)
);

OAI21xp5_ASAP7_75t_L g2178 ( 
.A1(n_2166),
.A2(n_2119),
.B(n_2115),
.Y(n_2178)
);

A2O1A1Ixp33_ASAP7_75t_SL g2179 ( 
.A1(n_2174),
.A2(n_2113),
.B(n_1980),
.C(n_2119),
.Y(n_2179)
);

OAI221xp5_ASAP7_75t_SL g2180 ( 
.A1(n_2167),
.A2(n_2175),
.B1(n_2169),
.B2(n_2173),
.C(n_2165),
.Y(n_2180)
);

OAI211xp5_ASAP7_75t_SL g2181 ( 
.A1(n_2174),
.A2(n_2176),
.B(n_2171),
.C(n_2168),
.Y(n_2181)
);

NAND3xp33_ASAP7_75t_L g2182 ( 
.A(n_2172),
.B(n_2142),
.C(n_2119),
.Y(n_2182)
);

AOI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_2166),
.A2(n_1983),
.B1(n_1985),
.B2(n_1980),
.Y(n_2183)
);

AOI21xp33_ASAP7_75t_SL g2184 ( 
.A1(n_2177),
.A2(n_1792),
.B(n_1983),
.Y(n_2184)
);

AOI221xp5_ASAP7_75t_L g2185 ( 
.A1(n_2181),
.A2(n_1980),
.B1(n_1983),
.B2(n_1985),
.C(n_1969),
.Y(n_2185)
);

AOI21x1_ASAP7_75t_L g2186 ( 
.A1(n_2182),
.A2(n_2003),
.B(n_1969),
.Y(n_2186)
);

OR3x1_ASAP7_75t_L g2187 ( 
.A(n_2180),
.B(n_1780),
.C(n_1777),
.Y(n_2187)
);

NOR3xp33_ASAP7_75t_SL g2188 ( 
.A(n_2178),
.B(n_1900),
.C(n_1986),
.Y(n_2188)
);

AOI22xp5_ASAP7_75t_L g2189 ( 
.A1(n_2183),
.A2(n_1985),
.B1(n_1930),
.B2(n_2035),
.Y(n_2189)
);

NOR5xp2_ASAP7_75t_L g2190 ( 
.A(n_2179),
.B(n_1962),
.C(n_1970),
.D(n_1975),
.E(n_1978),
.Y(n_2190)
);

AND3x1_ASAP7_75t_L g2191 ( 
.A(n_2188),
.B(n_1947),
.C(n_2010),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2186),
.Y(n_2192)
);

AOI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_2187),
.A2(n_1985),
.B1(n_2037),
.B2(n_2035),
.Y(n_2193)
);

NAND4xp75_ASAP7_75t_L g2194 ( 
.A(n_2185),
.B(n_2001),
.C(n_1999),
.D(n_1972),
.Y(n_2194)
);

XNOR2xp5_ASAP7_75t_L g2195 ( 
.A(n_2189),
.B(n_2184),
.Y(n_2195)
);

AOI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2194),
.A2(n_1985),
.B1(n_2190),
.B2(n_2037),
.Y(n_2196)
);

INVx2_ASAP7_75t_SL g2197 ( 
.A(n_2195),
.Y(n_2197)
);

NOR2xp67_ASAP7_75t_L g2198 ( 
.A(n_2192),
.B(n_2010),
.Y(n_2198)
);

OAI22xp5_ASAP7_75t_SL g2199 ( 
.A1(n_2197),
.A2(n_2191),
.B1(n_2193),
.B2(n_2048),
.Y(n_2199)
);

AOI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_2199),
.A2(n_2198),
.B1(n_2196),
.B2(n_2048),
.Y(n_2200)
);

AOI211x1_ASAP7_75t_L g2201 ( 
.A1(n_2200),
.A2(n_1972),
.B(n_1962),
.C(n_1987),
.Y(n_2201)
);

AO211x2_ASAP7_75t_L g2202 ( 
.A1(n_2200),
.A2(n_1970),
.B(n_1962),
.C(n_1987),
.Y(n_2202)
);

OAI22xp5_ASAP7_75t_SL g2203 ( 
.A1(n_2201),
.A2(n_1979),
.B1(n_1930),
.B2(n_1991),
.Y(n_2203)
);

OAI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_2202),
.A2(n_1965),
.B1(n_1968),
.B2(n_1966),
.Y(n_2204)
);

OAI21x1_ASAP7_75t_SL g2205 ( 
.A1(n_2204),
.A2(n_1799),
.B(n_1966),
.Y(n_2205)
);

OAI21xp5_ASAP7_75t_L g2206 ( 
.A1(n_2203),
.A2(n_2001),
.B(n_1999),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2205),
.B(n_1966),
.Y(n_2207)
);

OAI21xp5_ASAP7_75t_L g2208 ( 
.A1(n_2207),
.A2(n_2206),
.B(n_2001),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2208),
.Y(n_2209)
);

AOI221xp5_ASAP7_75t_L g2210 ( 
.A1(n_2209),
.A2(n_1970),
.B1(n_1987),
.B2(n_1975),
.C(n_1978),
.Y(n_2210)
);

AOI211xp5_ASAP7_75t_L g2211 ( 
.A1(n_2210),
.A2(n_1762),
.B(n_1947),
.C(n_1772),
.Y(n_2211)
);


endmodule