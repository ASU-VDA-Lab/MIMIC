module fake_jpeg_4369_n_224 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_224);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_18),
.B1(n_14),
.B2(n_22),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_22),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_R g54 ( 
.A(n_36),
.B(n_25),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_30),
.B1(n_28),
.B2(n_27),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_50),
.B1(n_39),
.B2(n_48),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_13),
.B1(n_18),
.B2(n_14),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_13),
.B1(n_18),
.B2(n_14),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

AO22x1_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_30),
.B1(n_28),
.B2(n_27),
.Y(n_50)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_40),
.A3(n_42),
.B1(n_28),
.B2(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_58),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_13),
.B1(n_18),
.B2(n_14),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_59),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_44),
.B1(n_36),
.B2(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_72),
.B1(n_46),
.B2(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_73),
.Y(n_91)
);

OA21x2_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_43),
.B(n_55),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_28),
.B1(n_45),
.B2(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_46),
.B1(n_57),
.B2(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_38),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_85),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_84),
.B1(n_87),
.B2(n_95),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_54),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_64),
.C(n_76),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_83),
.A2(n_35),
.B1(n_14),
.B2(n_26),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_61),
.B1(n_52),
.B2(n_46),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_56),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_92),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_45),
.B1(n_56),
.B2(n_35),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_94),
.Y(n_111)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_73),
.B1(n_75),
.B2(n_69),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_56),
.B(n_17),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_63),
.B(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_105),
.B(n_114),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_104),
.C(n_83),
.Y(n_118)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_116),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_83),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_79),
.B(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_72),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_34),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_92),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_96),
.Y(n_124)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_71),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_25),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_77),
.B1(n_60),
.B2(n_27),
.Y(n_135)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_82),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_118),
.C(n_119),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_84),
.C(n_81),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_121),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_105),
.B(n_99),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_88),
.Y(n_126)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_130),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_90),
.B1(n_91),
.B2(n_85),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_115),
.B1(n_114),
.B2(n_99),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_96),
.C(n_95),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_134),
.C(n_114),
.Y(n_150)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

AOI221xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_85),
.B1(n_91),
.B2(n_87),
.C(n_90),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_31),
.A3(n_23),
.B1(n_33),
.B2(n_26),
.C1(n_27),
.C2(n_32),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_133),
.B(n_123),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_42),
.C(n_29),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_103),
.B1(n_98),
.B2(n_108),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_98),
.B(n_101),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_109),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_134),
.A2(n_109),
.B1(n_113),
.B2(n_103),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_148),
.B1(n_122),
.B2(n_133),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_99),
.Y(n_146)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_141),
.Y(n_163)
);

AO22x1_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_111),
.B1(n_25),
.B2(n_116),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_126),
.B(n_42),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_121),
.B1(n_120),
.B2(n_119),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_125),
.A2(n_32),
.B(n_25),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_15),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_118),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_20),
.B(n_24),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_167),
.C(n_170),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_156),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_124),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_166),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_122),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_123),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_38),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_169),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_31),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_23),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_175),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_20),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_145),
.B1(n_148),
.B2(n_143),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_182),
.B1(n_167),
.B2(n_161),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_146),
.B(n_151),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_156),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_151),
.B1(n_142),
.B2(n_140),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_144),
.B1(n_26),
.B2(n_13),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_186),
.A2(n_188),
.B1(n_17),
.B2(n_27),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_33),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_163),
.C(n_161),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_170),
.C(n_160),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_33),
.C(n_26),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_187),
.B(n_20),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_195),
.B(n_198),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_19),
.Y(n_196)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_17),
.C(n_19),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_19),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_184),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_19),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_176),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_194),
.B(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_202),
.B(n_203),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_179),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_190),
.A2(n_24),
.B1(n_21),
.B2(n_177),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_197),
.A3(n_193),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_205),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_206),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_207),
.B(n_204),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_212),
.C(n_213),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_201),
.B(n_8),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_210),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_216),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_9),
.B(n_4),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_218),
.A2(n_219),
.B(n_10),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_10),
.C(n_11),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_221),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_0),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_0),
.Y(n_224)
);


endmodule