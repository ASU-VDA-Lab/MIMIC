module real_jpeg_27180_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_0),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_64),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_0),
.A2(n_47),
.B1(n_50),
.B2(n_64),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_1),
.A2(n_27),
.B1(n_83),
.B2(n_106),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_1),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_1),
.A2(n_27),
.B1(n_47),
.B2(n_50),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_3),
.A2(n_47),
.B1(n_50),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_3),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_5),
.A2(n_38),
.B1(n_47),
.B2(n_50),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_6),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_51),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_8),
.A2(n_47),
.B1(n_50),
.B2(n_66),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_9),
.B(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_9),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_SL g82 ( 
.A1(n_9),
.A2(n_26),
.B(n_43),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_9),
.A2(n_71),
.B1(n_83),
.B2(n_106),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_9),
.A2(n_34),
.B(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_9),
.B(n_34),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_9),
.B(n_39),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_9),
.A2(n_74),
.B1(n_76),
.B2(n_146),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_9),
.A2(n_25),
.B(n_161),
.Y(n_160)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_11),
.A2(n_47),
.B1(n_50),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_15),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_113),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_111),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_19),
.B(n_78),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_56),
.C(n_67),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_20),
.A2(n_21),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_40),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_41),
.C(n_45),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_37),
.B2(n_39),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_24),
.A2(n_29),
.B1(n_33),
.B2(n_160),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_30),
.Y(n_32)
);

AO22x1_ASAP7_75t_L g42 ( 
.A1(n_25),
.A2(n_26),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

OAI32xp33_ASAP7_75t_L g69 ( 
.A1(n_25),
.A2(n_30),
.A3(n_35),
.B1(n_70),
.B2(n_72),
.Y(n_69)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_26),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_29),
.A2(n_33),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_35),
.B1(n_59),
.B2(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_34),
.B(n_36),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_34),
.A2(n_50),
.A3(n_59),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_37),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_42),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_42),
.A2(n_43),
.B(n_106),
.C(n_107),
.Y(n_105)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_43),
.B(n_106),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_71),
.B(n_82),
.C(n_83),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_52),
.B2(n_54),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_46),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_54),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_46),
.A2(n_86),
.B1(n_139),
.B2(n_141),
.Y(n_138)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_50),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_47),
.B(n_60),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_47),
.B(n_151),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_49),
.Y(n_77)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_56),
.A2(n_67),
.B1(n_68),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_56),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_62),
.B2(n_65),
.Y(n_56)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_57),
.A2(n_58),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_57),
.A2(n_58),
.B1(n_122),
.B2(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_58),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_58),
.B(n_71),
.Y(n_147)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_63),
.A2(n_101),
.B1(n_103),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_65),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_69),
.B(n_73),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_70),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_71),
.B(n_76),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_74),
.A2(n_76),
.B1(n_140),
.B2(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_92),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_170),
.B(n_176),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_155),
.B(n_169),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_136),
.B(n_154),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_127),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_117),
.B(n_127),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_123),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_119),
.B1(n_123),
.B2(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_132),
.C(n_134),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_133),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_143),
.B(n_153),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_138),
.B(n_142),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_148),
.B(n_152),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_145),
.B(n_147),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_156),
.B(n_157),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_159),
.Y(n_165)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_165),
.C(n_168),
.Y(n_171)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);


endmodule