module fake_jpeg_11347_n_36 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_36);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_0),
.C(n_2),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_18),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_0),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.C(n_21),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_17),
.B(n_16),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_12),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_26),
.C(n_27),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_13),
.Y(n_27)
);

AOI221xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_16),
.B1(n_3),
.B2(n_1),
.C(n_13),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_31),
.C(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_13),
.C(n_5),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_29),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_SL g35 ( 
.A1(n_34),
.A2(n_33),
.B(n_9),
.C(n_10),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_35),
.B(n_7),
.Y(n_36)
);


endmodule