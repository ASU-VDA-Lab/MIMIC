module fake_jpeg_6748_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_43),
.A2(n_21),
.B1(n_40),
.B2(n_37),
.Y(n_74)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_46),
.B(n_49),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_50),
.Y(n_75)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_18),
.B(n_9),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_59),
.Y(n_79)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_18),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_53),
.A2(n_24),
.B1(n_36),
.B2(n_39),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_SL g57 ( 
.A1(n_19),
.A2(n_1),
.B(n_2),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_22),
.Y(n_68)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_64),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_41),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_66),
.A2(n_108),
.B1(n_28),
.B2(n_31),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_80),
.Y(n_115)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_88),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_20),
.B1(n_40),
.B2(n_37),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_73),
.A2(n_90),
.B1(n_95),
.B2(n_103),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_76),
.B1(n_97),
.B2(n_32),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_23),
.B1(n_35),
.B2(n_26),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_30),
.B1(n_7),
.B2(n_8),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_35),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_5),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_25),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_21),
.Y(n_89)
);

NAND4xp25_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_88),
.C(n_97),
.D(n_79),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_21),
.B1(n_40),
.B2(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_96),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_46),
.A2(n_24),
.B1(n_37),
.B2(n_36),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_97)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_102),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_27),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_44),
.A2(n_36),
.B1(n_39),
.B2(n_41),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_32),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_65),
.A2(n_39),
.B1(n_28),
.B2(n_31),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_112),
.A2(n_122),
.B(n_86),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_130),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_116),
.B(n_140),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_66),
.A2(n_30),
.B1(n_8),
.B2(n_9),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_142),
.B1(n_113),
.B2(n_114),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_66),
.A2(n_16),
.B(n_10),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_15),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_88),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

FAx1_ASAP7_75t_L g131 ( 
.A(n_66),
.B(n_5),
.CI(n_12),
.CON(n_131),
.SN(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_72),
.B(n_70),
.C(n_86),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_89),
.A2(n_85),
.B1(n_81),
.B2(n_83),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_133),
.A2(n_136),
.B1(n_83),
.B2(n_105),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_68),
.A2(n_13),
.B1(n_14),
.B2(n_89),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_134),
.A2(n_122),
.B1(n_116),
.B2(n_110),
.Y(n_175)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_137),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_85),
.A2(n_13),
.B1(n_14),
.B2(n_81),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_138),
.B(n_145),
.Y(n_179)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_87),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_82),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_68),
.A2(n_77),
.B1(n_104),
.B2(n_99),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_124),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_91),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_149),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_107),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_152),
.A2(n_162),
.B(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_121),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_160),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_155),
.A2(n_169),
.B1(n_148),
.B2(n_161),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_98),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_163),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_102),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_157),
.A2(n_144),
.B(n_119),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_93),
.Y(n_159)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_94),
.B(n_92),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_135),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_70),
.Y(n_165)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_118),
.Y(n_166)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_86),
.B(n_67),
.C(n_87),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_175),
.B1(n_128),
.B2(n_141),
.Y(n_185)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_115),
.A2(n_67),
.A3(n_87),
.B1(n_131),
.B2(n_125),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_67),
.Y(n_173)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_178),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_140),
.Y(n_178)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_143),
.A3(n_134),
.B1(n_110),
.B2(n_114),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_131),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_182),
.B(n_201),
.Y(n_231)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_193),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_185),
.A2(n_204),
.B1(n_206),
.B2(n_203),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_128),
.B1(n_141),
.B2(n_119),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_126),
.B(n_124),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_205),
.B(n_164),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_144),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_147),
.B(n_126),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_210),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_169),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_159),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_162),
.B(n_150),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_119),
.B1(n_148),
.B2(n_175),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_149),
.A2(n_156),
.B(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_153),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_157),
.B(n_166),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_211),
.B(n_160),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_212),
.A2(n_170),
.B1(n_167),
.B2(n_157),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_171),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_214),
.B(n_224),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_197),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_225),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_155),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_219),
.C(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_188),
.C(n_206),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_220),
.A2(n_207),
.B(n_187),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_221),
.A2(n_170),
.B1(n_200),
.B2(n_157),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_222),
.A2(n_190),
.B1(n_202),
.B2(n_211),
.Y(n_256)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_228),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_179),
.C(n_178),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_183),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_232),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_188),
.A2(n_146),
.B(n_161),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_236),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_196),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_200),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_238),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_179),
.C(n_165),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_237),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_180),
.C(n_172),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_185),
.B1(n_186),
.B2(n_182),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_240),
.A2(n_232),
.B1(n_223),
.B2(n_208),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_222),
.B(n_194),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_218),
.C(n_238),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_244),
.A2(n_181),
.B1(n_184),
.B2(n_193),
.Y(n_275)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_250),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_186),
.B1(n_209),
.B2(n_202),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_256),
.B1(n_231),
.B2(n_207),
.Y(n_266)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

OAI322xp33_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_213),
.A3(n_219),
.B1(n_230),
.B2(n_227),
.C1(n_167),
.C2(n_224),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_187),
.Y(n_269)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_216),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_254),
.Y(n_271)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

NOR3xp33_ASAP7_75t_SL g257 ( 
.A(n_213),
.B(n_167),
.C(n_189),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_257),
.B(n_214),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_189),
.Y(n_258)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_236),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_269),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_229),
.B1(n_217),
.B2(n_221),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_262),
.A2(n_266),
.B1(n_268),
.B2(n_272),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_242),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_247),
.Y(n_277)
);

OA22x2_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_220),
.B1(n_231),
.B2(n_215),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_226),
.C(n_228),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_251),
.C(n_274),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_250),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_223),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_251),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_248),
.B1(n_265),
.B2(n_259),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_278),
.Y(n_292)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_282),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_284),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_283),
.B(n_285),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_270),
.B(n_243),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_263),
.Y(n_286)
);

OAI31xp33_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_262),
.A3(n_255),
.B(n_243),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_246),
.B(n_239),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_268),
.Y(n_289)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_282),
.B(n_268),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_241),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_295),
.A2(n_296),
.B(n_258),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_271),
.B(n_241),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_266),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_301),
.C(n_302),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_239),
.Y(n_300)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_283),
.C(n_260),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_291),
.C(n_276),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_254),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_304),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_289),
.B1(n_255),
.B2(n_297),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_301),
.C(n_312),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_244),
.B1(n_292),
.B2(n_181),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_269),
.B(n_276),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_302),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_314),
.B(n_311),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_307),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_SL g319 ( 
.A(n_318),
.B(n_308),
.C(n_317),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_311),
.Y(n_320)
);


endmodule