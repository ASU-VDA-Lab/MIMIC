module fake_jpeg_2984_n_57 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_57);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2x1_ASAP7_75t_R g23 ( 
.A(n_20),
.B(n_0),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NAND2x1_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_1),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_16),
.B1(n_21),
.B2(n_20),
.Y(n_28)
);

NOR4xp25_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_23),
.C(n_25),
.D(n_4),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_17),
.B1(n_21),
.B2(n_16),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_19),
.B(n_3),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_34),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_17),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_2),
.C(n_5),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_19),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_39),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_45),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_10),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_39),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_50),
.B1(n_44),
.B2(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_6),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_44),
.B1(n_42),
.B2(n_7),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

NOR2xp67_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_45),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_53),
.A2(n_47),
.B(n_12),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_55),
.A2(n_11),
.B(n_14),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_54),
.Y(n_57)
);


endmodule