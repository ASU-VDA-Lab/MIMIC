module fake_jpeg_22065_n_132 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_17),
.A2(n_14),
.B1(n_25),
.B2(n_24),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_19),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_21),
.B1(n_26),
.B2(n_22),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_19),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_7),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_15),
.Y(n_44)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_53),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_61),
.B1(n_28),
.B2(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_18),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_24),
.B1(n_26),
.B2(n_22),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_59),
.B1(n_20),
.B2(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_57),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_21),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_32),
.A2(n_24),
.B1(n_20),
.B2(n_28),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_35),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_SL g93 ( 
.A(n_66),
.B(n_61),
.C(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_62),
.B1(n_43),
.B2(n_61),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_32),
.C(n_29),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_66),
.C(n_56),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_55),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_20),
.B1(n_32),
.B2(n_13),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_75),
.B1(n_77),
.B2(n_45),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_20),
.B1(n_32),
.B2(n_9),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_10),
.B(n_52),
.C(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_89),
.C(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_64),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_88),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_90),
.B1(n_91),
.B2(n_77),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_59),
.C(n_60),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_96),
.C(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_47),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_79),
.B(n_74),
.Y(n_89)
);

OA21x2_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_61),
.B(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_44),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_99),
.B1(n_43),
.B2(n_81),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_67),
.B1(n_71),
.B2(n_64),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_104),
.B1(n_96),
.B2(n_87),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_106),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_57),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_88),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_112),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_98),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_94),
.C(n_92),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_115),
.C(n_101),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_82),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_118),
.B(n_111),
.Y(n_123)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_120),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_101),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_102),
.C(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_121),
.B(n_115),
.Y(n_124)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_120),
.C(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_118),
.B1(n_113),
.B2(n_62),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_127),
.C(n_49),
.Y(n_129)
);

OAI21x1_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_81),
.B(n_82),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_10),
.C(n_76),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_78),
.Y(n_132)
);


endmodule