module fake_jpeg_17128_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_3),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_19),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

AND2x4_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_17),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_19),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_30),
.B(n_21),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_49),
.B(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_24),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_34),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_30),
.C(n_33),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_80),
.C(n_54),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_74),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_70),
.Y(n_85)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_64),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_66),
.B(n_73),
.Y(n_92)
);

CKINVDCx9p33_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_15),
.B1(n_35),
.B2(n_37),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_57),
.B1(n_69),
.B2(n_38),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_37),
.B1(n_35),
.B2(n_21),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_83),
.B1(n_37),
.B2(n_38),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_23),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_75),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_21),
.B(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_40),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_79),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_39),
.C(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_42),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_37),
.B1(n_15),
.B2(n_34),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_86),
.A2(n_90),
.B1(n_106),
.B2(n_28),
.Y(n_138)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_38),
.B1(n_32),
.B2(n_34),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_98),
.B1(n_75),
.B2(n_76),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_38),
.B1(n_32),
.B2(n_34),
.Y(n_98)
);

HAxp5_ASAP7_75t_SL g135 ( 
.A(n_99),
.B(n_17),
.CON(n_135),
.SN(n_135)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_74),
.B1(n_56),
.B2(n_58),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_108),
.B1(n_112),
.B2(n_42),
.Y(n_128)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_102),
.B(n_103),
.CI(n_104),
.CON(n_118),
.SN(n_118)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_51),
.C(n_33),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_16),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_61),
.A2(n_27),
.B(n_24),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_56),
.A2(n_52),
.B1(n_32),
.B2(n_34),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_80),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_32),
.B1(n_15),
.B2(n_28),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_113),
.B(n_117),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_116),
.B1(n_130),
.B2(n_89),
.Y(n_152)
);

OAI22x1_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_90),
.B1(n_87),
.B2(n_99),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_125),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

CKINVDCx11_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_122),
.B(n_123),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_83),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_41),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_128),
.B(n_33),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_65),
.B1(n_60),
.B2(n_28),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_41),
.Y(n_131)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_85),
.B(n_26),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_133),
.B(n_26),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_29),
.B(n_31),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_54),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_95),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_138),
.A2(n_103),
.B1(n_100),
.B2(n_112),
.Y(n_140)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_152),
.B1(n_166),
.B2(n_124),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_104),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_153),
.C(n_155),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_86),
.B1(n_102),
.B2(n_93),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_144),
.A2(n_145),
.B1(n_149),
.B2(n_161),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_125),
.B1(n_134),
.B2(n_119),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_98),
.B(n_108),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_121),
.B1(n_129),
.B2(n_139),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_95),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_154),
.B(n_156),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_95),
.C(n_84),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_46),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_169),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_62),
.B(n_1),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_39),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_115),
.A2(n_91),
.B1(n_28),
.B2(n_33),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_54),
.B1(n_62),
.B2(n_22),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_39),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_39),
.Y(n_165)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_128),
.A2(n_91),
.B1(n_39),
.B2(n_27),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_129),
.B1(n_120),
.B2(n_127),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_16),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_120),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_171),
.B(n_29),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_172),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_173),
.B(n_171),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_142),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_178),
.A2(n_181),
.B(n_183),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_179),
.B(n_180),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_132),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_182),
.B(n_184),
.Y(n_220)
);

AND2x6_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_14),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_94),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_188),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_94),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_187),
.B(n_195),
.Y(n_222)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_27),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_191),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_109),
.B1(n_31),
.B2(n_23),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_192),
.B1(n_196),
.B2(n_151),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_41),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_144),
.A2(n_77),
.B1(n_54),
.B2(n_62),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_150),
.B1(n_160),
.B2(n_151),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_25),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_143),
.A2(n_149),
.B1(n_145),
.B2(n_148),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_200),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_143),
.B(n_25),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_18),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_18),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_161),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_0),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_206),
.B1(n_227),
.B2(n_229),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_204),
.B1(n_198),
.B2(n_177),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_141),
.C(n_158),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_217),
.C(n_224),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_211),
.B(n_173),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_189),
.B(n_169),
.Y(n_212)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_140),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_225),
.B(n_203),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_168),
.C(n_136),
.Y(n_217)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_136),
.C(n_25),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_136),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_228),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_177),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_18),
.Y(n_228)
);

OAI22x1_ASAP7_75t_SL g229 ( 
.A1(n_196),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_175),
.B1(n_193),
.B2(n_192),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_218),
.B1(n_213),
.B2(n_227),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_226),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_206),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_241),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_186),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_237),
.B(n_245),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_205),
.B1(n_219),
.B2(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_174),
.B1(n_178),
.B2(n_183),
.Y(n_243)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_224),
.B(n_200),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_182),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_213),
.Y(n_265)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_175),
.B(n_181),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_SL g266 ( 
.A1(n_248),
.A2(n_188),
.B(n_222),
.C(n_223),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_207),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_265),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_207),
.C(n_214),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_263),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_235),
.A2(n_240),
.B1(n_231),
.B2(n_249),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_208),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_248),
.B(n_230),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_233),
.C(n_237),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_269),
.C(n_271),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_245),
.C(n_246),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_241),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_230),
.C(n_236),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_278),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_276),
.Y(n_288)
);

AO21x2_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_238),
.B(n_185),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_277),
.A2(n_272),
.B1(n_275),
.B2(n_271),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_262),
.B(n_250),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_212),
.C(n_201),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_266),
.Y(n_283)
);

OAI21x1_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_211),
.B(n_8),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_280),
.A2(n_252),
.B1(n_256),
.B2(n_254),
.Y(n_281)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_253),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_284),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_269),
.C(n_267),
.Y(n_297)
);

A2O1A1Ixp33_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_266),
.B(n_8),
.C(n_9),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_8),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_292),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_13),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_279),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_12),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_286),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_267),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_297),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_22),
.C(n_12),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_300),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_1),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_301),
.A2(n_284),
.B(n_289),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_304),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_306),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_291),
.B1(n_288),
.B2(n_3),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_11),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_301),
.C(n_298),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_302),
.B(n_293),
.Y(n_311)
);

AOI332xp33_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_310),
.A3(n_306),
.B1(n_296),
.B2(n_308),
.B3(n_9),
.C1(n_10),
.C2(n_6),
.Y(n_312)
);

NOR3xp33_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_10),
.C(n_9),
.Y(n_313)
);

OAI321xp33_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_1),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_314),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_315)
);

AOI21x1_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_4),
.B(n_7),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_4),
.B1(n_7),
.B2(n_280),
.Y(n_317)
);


endmodule