module fake_netlist_1_12738_n_33 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
NAND2x1p5_ASAP7_75t_L g13 ( .A(n_0), .B(n_10), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
NOR2xp67_ASAP7_75t_L g15 ( .A(n_8), .B(n_9), .Y(n_15) );
BUFx4f_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
NOR2xp67_ASAP7_75t_L g17 ( .A(n_12), .B(n_1), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_16), .B(n_14), .Y(n_19) );
INVx2_ASAP7_75t_SL g20 ( .A(n_19), .Y(n_20) );
OAI222xp33_ASAP7_75t_L g21 ( .A1(n_18), .A2(n_13), .B1(n_14), .B2(n_12), .C1(n_11), .C2(n_17), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_13), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
AOI31xp33_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_13), .A3(n_20), .B(n_21), .Y(n_24) );
AOI222xp33_ASAP7_75t_L g25 ( .A1(n_22), .A2(n_21), .B1(n_11), .B2(n_14), .C1(n_15), .C2(n_5), .Y(n_25) );
NOR3xp33_ASAP7_75t_L g26 ( .A(n_24), .B(n_22), .C(n_15), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_24), .B(n_23), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
OR2x2_ASAP7_75t_L g29 ( .A(n_26), .B(n_23), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_25), .B1(n_2), .B2(n_3), .Y(n_30) );
OAI22x1_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_31) );
OAI311xp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_5), .A3(n_6), .B1(n_7), .C1(n_8), .Y(n_32) );
AOI22x1_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_31), .B1(n_6), .B2(n_7), .Y(n_33) );
endmodule