module fake_jpeg_8370_n_106 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_6),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_68),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_3),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_74),
.B1(n_75),
.B2(n_61),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_57),
.B1(n_11),
.B2(n_12),
.Y(n_78)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_73),
.Y(n_83)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_81),
.B1(n_84),
.B2(n_49),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_82),
.B1(n_47),
.B2(n_13),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_75),
.A2(n_66),
.B1(n_64),
.B2(n_56),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_46),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_54),
.B1(n_52),
.B2(n_50),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_89),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_9),
.B1(n_14),
.B2(n_18),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_93),
.A2(n_91),
.B1(n_90),
.B2(n_86),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_85),
.C(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_95),
.B(n_85),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_96),
.Y(n_97)
);

OAI211xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_92),
.B(n_20),
.C(n_24),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_19),
.B(n_26),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_27),
.C(n_28),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_30),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_31),
.B1(n_35),
.B2(n_37),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_38),
.B(n_41),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_42),
.B(n_43),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_45),
.Y(n_106)
);


endmodule