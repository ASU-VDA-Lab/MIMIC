module fake_jpeg_19743_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_17),
.B(n_19),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_22),
.B1(n_15),
.B2(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_14),
.B(n_1),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

AOI21xp33_ASAP7_75t_SL g21 ( 
.A1(n_15),
.A2(n_2),
.B(n_4),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_20),
.B(n_8),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_33),
.B(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.C(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_11),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_28),
.C(n_27),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_12),
.C(n_10),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_33),
.B(n_29),
.C(n_27),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_36),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_42),
.C(n_6),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_37),
.B1(n_38),
.B2(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_48),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_53),
.A2(n_51),
.B(n_10),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_10),
.Y(n_55)
);


endmodule