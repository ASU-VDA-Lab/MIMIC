module real_jpeg_23831_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx3_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_1),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_1),
.B(n_61),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_1),
.B(n_43),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_1),
.B(n_36),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_1),
.B(n_40),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_1),
.B(n_50),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_1),
.B(n_133),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_1),
.B(n_210),
.Y(n_378)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_2),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_2),
.B(n_43),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_2),
.B(n_40),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_2),
.B(n_50),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_2),
.B(n_303),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_3),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_3),
.B(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_3),
.B(n_43),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_3),
.B(n_36),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_3),
.B(n_40),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_3),
.B(n_50),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_3),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_3),
.B(n_303),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_6),
.B(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_6),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_6),
.B(n_43),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_6),
.B(n_36),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_6),
.B(n_40),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_6),
.B(n_50),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_6),
.B(n_133),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_6),
.B(n_210),
.Y(n_365)
);

INVx8_ASAP7_75t_SL g135 ( 
.A(n_7),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_8),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_43),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_8),
.B(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_8),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_8),
.B(n_50),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_8),
.B(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_8),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_9),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_9),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_9),
.B(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_9),
.B(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_9),
.B(n_40),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_9),
.B(n_50),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_9),
.B(n_133),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_9),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_10),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_10),
.B(n_36),
.Y(n_92)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_10),
.B(n_61),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_10),
.B(n_133),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_12),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_12),
.B(n_61),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_12),
.B(n_43),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_12),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_12),
.B(n_50),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_12),
.B(n_133),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_12),
.B(n_210),
.Y(n_331)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_13),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_14),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_14),
.B(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_14),
.B(n_36),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_14),
.B(n_40),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_14),
.B(n_50),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_14),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_14),
.B(n_229),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_16),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_16),
.B(n_61),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_16),
.B(n_43),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_16),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_16),
.B(n_40),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_16),
.B(n_50),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_16),
.B(n_229),
.Y(n_350)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_17),
.Y(n_108)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_384),
.B(n_385),
.C(n_389),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_374),
.C(n_383),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_359),
.C(n_360),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_337),
.C(n_338),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_307),
.C(n_308),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_281),
.C(n_282),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_249),
.C(n_250),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_212),
.C(n_213),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_175),
.C(n_176),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_142),
.C(n_143),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_113),
.C(n_114),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_72),
.C(n_85),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_53),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_45),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_33),
.B(n_45),
.C(n_53),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.C(n_41),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_34),
.A2(n_35),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_36),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_40),
.Y(n_222)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_46),
.B(n_48),
.C(n_49),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_63),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_54),
.B(n_64),
.C(n_65),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_61),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_67),
.B(n_71),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.C(n_84),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_77),
.B1(n_84),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_83),
.B(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_109),
.C(n_110),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_94),
.C(n_99),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_92),
.C(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.C(n_104),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_102),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_108),
.B(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_128),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_129),
.C(n_141),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_124),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_123),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_123),
.C(n_124),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_118),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_122),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_124),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_126),
.CI(n_127),
.CON(n_124),
.SN(n_124)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_126),
.C(n_127),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_141),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_139),
.B2(n_140),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_132),
.Y(n_138)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_134),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_134),
.B(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_134),
.B(n_219),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_134),
.B(n_234),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_138),
.C(n_140),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_158),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_147),
.C(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_154),
.C(n_157),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_149),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_151),
.CI(n_152),
.CON(n_149),
.SN(n_149)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_151),
.C(n_152),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_165),
.C(n_173),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_165),
.B1(n_173),
.B2(n_174),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_161),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_163),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_164),
.B(n_201),
.C(n_202),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_165),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_171),
.C(n_172),
.Y(n_196)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx11_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_169),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_197),
.B2(n_211),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_198),
.C(n_199),
.Y(n_212)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_181),
.C(n_190),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_190),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_186),
.C(n_189),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_184),
.B(n_234),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_188),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_195),
.C(n_196),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_194),
.Y(n_195)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_209),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_207),
.C(n_209),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_206),
.B(n_234),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_247),
.B2(n_248),
.Y(n_213)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_238),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_238),
.C(n_247),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_225),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_226),
.C(n_227),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_218),
.B(n_221),
.C(n_223),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_230),
.B1(n_231),
.B2(n_237),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_228),
.Y(n_237)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_233),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_236),
.C(n_237),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_232),
.B(n_256),
.C(n_259),
.Y(n_305)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_245),
.C(n_246),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_253),
.C(n_280),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_267),
.B2(n_280),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_262),
.C(n_263),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_259),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_259),
.A2(n_260),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_SL g322 ( 
.A(n_259),
.B(n_286),
.C(n_289),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g391 ( 
.A(n_263),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_265),
.CI(n_266),
.CON(n_263),
.SN(n_263)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_265),
.C(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_270),
.C(n_271),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_279),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_275),
.C(n_277),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_274),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_275),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_276),
.A2(n_277),
.B1(n_302),
.B2(n_304),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_277),
.B(n_304),
.C(n_305),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_306),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_296),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_296),
.C(n_306),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_291),
.C(n_292),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_288),
.A2(n_289),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_SL g348 ( 
.A(n_289),
.B(n_315),
.C(n_317),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g394 ( 
.A(n_292),
.Y(n_394)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.CI(n_295),
.CON(n_292),
.SN(n_292)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_294),
.C(n_295),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_299),
.C(n_300),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_305),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_302),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_311),
.C(n_324),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_323),
.B2(n_324),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_319),
.B2(n_320),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_321),
.C(n_322),
.Y(n_340)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_317),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_317),
.A2(n_318),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_317),
.B(n_353),
.C(n_354),
.Y(n_366)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_327),
.C(n_330),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_330),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_333),
.C(n_336),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_335),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_339),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.Y(n_338)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_339),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_341),
.C(n_358),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_347),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_348),
.C(n_349),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_363),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_343),
.B(n_361),
.C(n_363),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_345),
.CI(n_346),
.CON(n_343),
.SN(n_343)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_351),
.B1(n_354),
.B2(n_355),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_350),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_351),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_352),
.A2(n_353),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_370),
.C(n_373),
.Y(n_376)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_356),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_366),
.C(n_367),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_372),
.B2(n_373),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_370),
.A2(n_371),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_SL g390 ( 
.A(n_371),
.B(n_378),
.C(n_381),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_372),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_382),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_377),
.C(n_382),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_380),
.A2(n_381),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_381),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_390),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_388),
.Y(n_389)
);


endmodule