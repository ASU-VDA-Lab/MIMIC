module fake_jpeg_31057_n_305 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_305);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_288;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_5),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_52),
.Y(n_66)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_26),
.B(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_41),
.Y(n_67)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_35),
.Y(n_70)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_56),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_58),
.Y(n_92)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_61),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_SL g64 ( 
.A1(n_53),
.A2(n_25),
.B(n_32),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_64),
.B(n_32),
.C(n_34),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_67),
.B(n_79),
.Y(n_110)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_70),
.B(n_75),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_28),
.B1(n_27),
.B2(n_39),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_39),
.B1(n_31),
.B2(n_30),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_46),
.B(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_35),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_80),
.B(n_83),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_81),
.A2(n_32),
.B1(n_34),
.B2(n_4),
.Y(n_132)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_20),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_84),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_19),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_86),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_22),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_87),
.Y(n_137)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_43),
.A2(n_28),
.B1(n_32),
.B2(n_42),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_43),
.B(n_40),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_43),
.B(n_40),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_58),
.B(n_24),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_24),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_23),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_51),
.B(n_23),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_52),
.B(n_22),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_98),
.Y(n_109)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_111),
.A2(n_71),
.B1(n_82),
.B2(n_97),
.Y(n_148)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_122),
.A2(n_124),
.B1(n_131),
.B2(n_76),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_64),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_73),
.C(n_72),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_65),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_134),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_68),
.A2(n_32),
.B1(n_34),
.B2(n_4),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_78),
.B1(n_89),
.B2(n_88),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_2),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_90),
.A2(n_34),
.B1(n_4),
.B2(n_5),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_79),
.B(n_108),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_129),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_144),
.B(n_151),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_124),
.B1(n_122),
.B2(n_118),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_173),
.B1(n_109),
.B2(n_139),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_148),
.B(n_77),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_149),
.B(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_85),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_161),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_66),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_115),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_152),
.B(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_110),
.B(n_102),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_90),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_154),
.A2(n_156),
.B(n_103),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_102),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_71),
.B(n_97),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_72),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_158),
.Y(n_188)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_90),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_71),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_170),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_119),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_3),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_113),
.C(n_121),
.Y(n_186)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_126),
.B(n_78),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_92),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_121),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_138),
.B1(n_77),
.B2(n_107),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_177),
.A2(n_182),
.B1(n_194),
.B2(n_160),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_172),
.A2(n_116),
.B1(n_119),
.B2(n_117),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_180),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_161),
.A2(n_117),
.B1(n_109),
.B2(n_139),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_133),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_183),
.C(n_186),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_105),
.B1(n_141),
.B2(n_114),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_150),
.B(n_92),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_185),
.B(n_198),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_114),
.C(n_92),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_201),
.C(n_147),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_174),
.B(n_163),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_105),
.B1(n_96),
.B2(n_95),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_200),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_76),
.B1(n_107),
.B2(n_93),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_154),
.A2(n_96),
.B1(n_95),
.B2(n_73),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_138),
.C(n_112),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_103),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_157),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_148),
.B(n_156),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_210),
.B(n_213),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_149),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_211),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_169),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_217),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_188),
.B(n_171),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_218),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_223),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_180),
.B1(n_179),
.B2(n_192),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_204),
.B(n_194),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_227),
.Y(n_236)
);

AOI221xp5_ASAP7_75t_L g226 ( 
.A1(n_176),
.A2(n_159),
.B1(n_157),
.B2(n_173),
.C(n_162),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_184),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_178),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_238),
.B1(n_241),
.B2(n_215),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_220),
.C(n_186),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_233),
.C(n_242),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_237),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_201),
.C(n_183),
.Y(n_233)
);

OAI321xp33_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_176),
.A3(n_184),
.B1(n_185),
.B2(n_181),
.C(n_202),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_204),
.B1(n_177),
.B2(n_182),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_189),
.C(n_187),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_187),
.C(n_162),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_246),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_160),
.C(n_195),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_213),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_227),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_250),
.Y(n_267)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_251),
.B(n_252),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_240),
.A2(n_222),
.B(n_208),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_211),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_260),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_226),
.B1(n_214),
.B2(n_218),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_205),
.B1(n_219),
.B2(n_209),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_219),
.B1(n_209),
.B2(n_217),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_261),
.B1(n_255),
.B2(n_239),
.Y(n_266)
);

AOI321xp33_ASAP7_75t_L g260 ( 
.A1(n_242),
.A2(n_216),
.A3(n_207),
.B1(n_224),
.B2(n_225),
.C(n_164),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_207),
.B1(n_195),
.B2(n_165),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_230),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_264),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_229),
.C(n_230),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_269),
.C(n_270),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_146),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_245),
.C(n_246),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_232),
.C(n_234),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_234),
.C(n_244),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_259),
.C(n_257),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_279),
.Y(n_289)
);

NAND2xp33_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_249),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_277),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_260),
.Y(n_278)
);

AOI31xp33_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_270),
.A3(n_268),
.B(n_273),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_272),
.A2(n_261),
.B1(n_252),
.B2(n_165),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_281),
.B(n_283),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_263),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_271),
.B(n_3),
.Y(n_282)
);

OAI221xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_146),
.C(n_164),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_285),
.A2(n_287),
.B(n_274),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_275),
.A2(n_146),
.B1(n_93),
.B2(n_262),
.Y(n_287)
);

AOI31xp33_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_164),
.A3(n_6),
.B(n_7),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_283),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_10),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_291),
.B(n_296),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_293),
.B(n_11),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_287),
.A2(n_276),
.B(n_9),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_295),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_8),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_284),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_298),
.B(n_299),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_11),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_297),
.B(n_12),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_303),
.A2(n_301),
.B(n_13),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_11),
.Y(n_305)
);


endmodule