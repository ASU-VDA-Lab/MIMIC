module fake_jpeg_12908_n_291 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_45),
.Y(n_109)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_61),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_51),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_63),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_21),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_67),
.Y(n_90)
);

INVx2_ASAP7_75t_R g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_108),
.B1(n_86),
.B2(n_89),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_80),
.B(n_5),
.Y(n_127)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_85),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_68),
.A2(n_39),
.B1(n_33),
.B2(n_29),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_86),
.A2(n_89),
.B(n_95),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_29),
.B1(n_41),
.B2(n_35),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_27),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_91),
.B(n_97),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_27),
.B1(n_35),
.B2(n_34),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_94),
.B1(n_110),
.B2(n_4),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_43),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_48),
.A2(n_23),
.B1(n_25),
.B2(n_28),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_31),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_54),
.B(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_98),
.B(n_99),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_28),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_55),
.B(n_25),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_100),
.B(n_10),
.Y(n_145)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_56),
.B(n_0),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_104),
.Y(n_113)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_60),
.A2(n_23),
.B1(n_36),
.B2(n_4),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_47),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_17),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_112),
.B(n_118),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_SL g156 ( 
.A(n_113),
.B(n_74),
.C(n_103),
.Y(n_156)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_115),
.B(n_140),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_134),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_15),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g172 ( 
.A(n_119),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_119),
.B1(n_125),
.B2(n_113),
.Y(n_165)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_1),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_124),
.A2(n_140),
.B1(n_144),
.B2(n_141),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_142),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_129),
.A2(n_77),
.B1(n_83),
.B2(n_96),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_131),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_76),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_15),
.B(n_8),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_93),
.B(n_84),
.Y(n_166)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_141),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_102),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_87),
.B(n_6),
.C(n_9),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_79),
.B(n_6),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_9),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_74),
.A2(n_9),
.B(n_10),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_121),
.B(n_124),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_11),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_74),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_79),
.B(n_11),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_84),
.B(n_72),
.C(n_93),
.Y(n_160)
);

OR2x4_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_12),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_166),
.B(n_123),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_173),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_159),
.B(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_135),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_162),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_72),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_165),
.A2(n_167),
.B1(n_157),
.B2(n_161),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_114),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_169),
.Y(n_194)
);

AOI32xp33_ASAP7_75t_L g170 ( 
.A1(n_116),
.A2(n_77),
.A3(n_83),
.B1(n_96),
.B2(n_147),
.Y(n_170)
);

AOI32xp33_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_125),
.A3(n_123),
.B1(n_137),
.B2(n_134),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_115),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

NOR2x1_ASAP7_75t_R g173 ( 
.A(n_144),
.B(n_136),
.Y(n_173)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_175),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_172),
.B1(n_160),
.B2(n_148),
.Y(n_210)
);

AO22x1_ASAP7_75t_SL g181 ( 
.A1(n_178),
.A2(n_122),
.B1(n_135),
.B2(n_117),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_185),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_201),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_184),
.A2(n_188),
.B(n_167),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_143),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_143),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_190),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_117),
.B(n_120),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_194),
.B(n_183),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_120),
.B(n_126),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_132),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_168),
.Y(n_191)
);

A2O1A1O1Ixp25_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_192),
.B(n_204),
.C(n_172),
.D(n_149),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_157),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_158),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_172),
.Y(n_216)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_178),
.A2(n_151),
.B1(n_173),
.B2(n_170),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_182),
.B1(n_179),
.B2(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_174),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_152),
.B(n_162),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_156),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_211),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_223),
.B1(n_181),
.B2(n_205),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_192),
.B(n_154),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_217),
.Y(n_234)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_149),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_216),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_169),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_196),
.B(n_189),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_219),
.B(n_226),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_175),
.B(n_153),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_175),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_220),
.B(n_198),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_194),
.A2(n_153),
.B1(n_174),
.B2(n_202),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_240),
.B1(n_243),
.B2(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

BUFx12_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_238),
.Y(n_244)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_237),
.A2(n_239),
.B1(n_208),
.B2(n_218),
.Y(n_245)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_221),
.Y(n_239)
);

NAND5xp2_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_199),
.C(n_195),
.D(n_180),
.E(n_181),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_212),
.B(n_225),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_222),
.A2(n_188),
.B1(n_181),
.B2(n_199),
.Y(n_243)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_206),
.C(n_220),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_253),
.C(n_254),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_247),
.A2(n_255),
.B1(n_241),
.B2(n_237),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_208),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_234),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_234),
.B(n_211),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_223),
.B1(n_225),
.B2(n_207),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_229),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_262),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_230),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_260),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_197),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_244),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_255),
.Y(n_267)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_248),
.B1(n_249),
.B2(n_235),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_259),
.C(n_246),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_267),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_269),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_252),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_254),
.C(n_233),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_257),
.B(n_228),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_272),
.B(n_261),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_256),
.A2(n_233),
.B1(n_241),
.B2(n_226),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_263),
.B1(n_240),
.B2(n_256),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_278),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_271),
.C(n_199),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_261),
.C(n_264),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_268),
.B1(n_270),
.B2(n_273),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_282),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_R g283 ( 
.A(n_277),
.B(n_267),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_280),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_285),
.B(n_275),
.Y(n_287)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_284),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_287),
.C(n_274),
.Y(n_288)
);

NOR3xp33_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_193),
.C(n_231),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_289),
.A2(n_197),
.B1(n_238),
.B2(n_200),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_188),
.Y(n_291)
);


endmodule