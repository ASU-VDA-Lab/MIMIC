module fake_jpeg_5291_n_210 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_210);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_8),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_42),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_8),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_19),
.B(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_25),
.B1(n_27),
.B2(n_15),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_48),
.A2(n_57),
.B1(n_61),
.B2(n_64),
.Y(n_112)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_52),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_25),
.B1(n_34),
.B2(n_44),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_50),
.A2(n_28),
.B1(n_29),
.B2(n_18),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_58),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_30),
.B1(n_31),
.B2(n_14),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_22),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_31),
.B1(n_14),
.B2(n_21),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_22),
.B1(n_21),
.B2(n_24),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_71),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_16),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_74),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_77),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_28),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_23),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_23),
.Y(n_83)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_35),
.B(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_28),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_28),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_114),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_85),
.B1(n_56),
.B2(n_51),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_67),
.B1(n_79),
.B2(n_87),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_111),
.B1(n_53),
.B2(n_84),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_83),
.B(n_62),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_54),
.C(n_47),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_107),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_82),
.B(n_79),
.C(n_67),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_28),
.B1(n_29),
.B2(n_18),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_76),
.B1(n_74),
.B2(n_55),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_29),
.B1(n_18),
.B2(n_2),
.Y(n_111)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_119),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_99),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_120),
.B(n_127),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_102),
.C(n_111),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_59),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_49),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_129),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_84),
.B1(n_51),
.B2(n_56),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_135),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_105),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_58),
.B1(n_78),
.B2(n_68),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_18),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_78),
.B(n_29),
.C(n_18),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_103),
.B(n_114),
.C(n_100),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_59),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_0),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_141),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_29),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_137),
.B(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_92),
.A2(n_59),
.B1(n_70),
.B2(n_4),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_1),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_94),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_9),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_1),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_88),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_149),
.C(n_151),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_152),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_110),
.C(n_90),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_90),
.C(n_88),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_160),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_108),
.C(n_113),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_120),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_161),
.B(n_131),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_108),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_164),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_120),
.A2(n_113),
.B(n_103),
.C(n_4),
.D(n_5),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_163),
.B(n_127),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_1),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_160),
.C(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_173),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_139),
.Y(n_173)
);

OAI321xp33_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_120),
.A3(n_133),
.B1(n_118),
.B2(n_128),
.C(n_141),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_144),
.B(n_149),
.C(n_163),
.D(n_164),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_154),
.B(n_137),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_131),
.A3(n_127),
.B1(n_137),
.B2(n_138),
.C1(n_136),
.C2(n_123),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_179),
.B(n_155),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_SL g178 ( 
.A1(n_158),
.A2(n_125),
.A3(n_119),
.B1(n_132),
.B2(n_6),
.C1(n_10),
.C2(n_11),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_SL g188 ( 
.A(n_178),
.B(n_12),
.C(n_13),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_2),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_180),
.B(n_184),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_151),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_186),
.C(n_166),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_148),
.B1(n_143),
.B2(n_159),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_143),
.B1(n_152),
.B2(n_153),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_189),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_173),
.A2(n_150),
.B1(n_91),
.B2(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_167),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_169),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_182),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_196),
.C(n_186),
.Y(n_199)
);

AOI322xp5_ASAP7_75t_L g196 ( 
.A1(n_187),
.A2(n_171),
.A3(n_170),
.B1(n_172),
.B2(n_179),
.C1(n_147),
.C2(n_100),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_187),
.C(n_180),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_199),
.C(n_200),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_183),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_197),
.C(n_185),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_202),
.A2(n_197),
.B(n_191),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_93),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_207),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_206),
.C(n_203),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_209),
.Y(n_210)
);


endmodule