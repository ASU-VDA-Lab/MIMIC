module fake_jpeg_22465_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

OR2x2_ASAP7_75t_L g9 ( 
.A(n_7),
.B(n_6),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_17),
.A2(n_14),
.B1(n_10),
.B2(n_13),
.Y(n_24)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx6p67_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

NOR2x1_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_22),
.B(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_21),
.B1(n_9),
.B2(n_15),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_22),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_19),
.B1(n_17),
.B2(n_20),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_37),
.B1(n_25),
.B2(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_21),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_18),
.B1(n_20),
.B2(n_14),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_32),
.B1(n_33),
.B2(n_28),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_1),
.B(n_2),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_25),
.C(n_10),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_39),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.C(n_44),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_39),
.C(n_25),
.Y(n_49)
);

AO21x1_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_4),
.B(n_5),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_4),
.C(n_7),
.Y(n_52)
);

BUFx24_ASAP7_75t_SL g53 ( 
.A(n_52),
.Y(n_53)
);


endmodule