module real_aes_7436_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g466 ( .A1(n_0), .A2(n_144), .B(n_467), .C(n_470), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_1), .B(n_461), .Y(n_472) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
INVx1_ASAP7_75t_L g182 ( .A(n_3), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_4), .B(n_145), .Y(n_544) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_5), .A2(n_123), .B1(n_124), .B2(n_430), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g430 ( .A(n_5), .Y(n_430) );
OAI22xp5_ASAP7_75t_SL g738 ( .A1(n_5), .A2(n_95), .B1(n_430), .B2(n_739), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_6), .A2(n_446), .B(n_493), .Y(n_492) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_7), .A2(n_151), .B(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_8), .A2(n_36), .B1(n_148), .B2(n_200), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_9), .B(n_151), .Y(n_168) );
AND2x6_ASAP7_75t_L g153 ( .A(n_10), .B(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_11), .A2(n_153), .B(n_449), .C(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_12), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_12), .B(n_38), .Y(n_435) );
INVx1_ASAP7_75t_L g135 ( .A(n_13), .Y(n_135) );
INVx1_ASAP7_75t_L g174 ( .A(n_14), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_15), .B(n_141), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_16), .B(n_145), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_17), .B(n_131), .Y(n_130) );
AO32x2_ASAP7_75t_L g211 ( .A1(n_18), .A2(n_151), .A3(n_152), .B1(n_171), .B2(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_19), .B(n_148), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_20), .B(n_131), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_21), .A2(n_54), .B1(n_148), .B2(n_200), .Y(n_214) );
AOI22xp33_ASAP7_75t_SL g208 ( .A1(n_22), .A2(n_80), .B1(n_141), .B2(n_148), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_23), .B(n_148), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_24), .A2(n_152), .B(n_449), .C(n_451), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_25), .A2(n_152), .B(n_449), .C(n_527), .Y(n_526) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_26), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_27), .A2(n_96), .B1(n_118), .B2(n_119), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_27), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_28), .B(n_190), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_29), .A2(n_446), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_30), .B(n_190), .Y(n_227) );
INVx2_ASAP7_75t_L g143 ( .A(n_31), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_32), .A2(n_481), .B(n_482), .C(n_486), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_33), .B(n_148), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_34), .B(n_190), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_35), .B(n_196), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_37), .Y(n_745) );
INVx1_ASAP7_75t_L g114 ( .A(n_38), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_39), .B(n_445), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_40), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_41), .B(n_145), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_42), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_43), .B(n_446), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_44), .A2(n_481), .B(n_486), .C(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_45), .B(n_148), .Y(n_161) );
INVx1_ASAP7_75t_L g468 ( .A(n_46), .Y(n_468) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_47), .A2(n_737), .B1(n_740), .B2(n_741), .Y(n_736) );
INVx1_ASAP7_75t_L g741 ( .A(n_47), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_48), .A2(n_89), .B1(n_200), .B2(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g507 ( .A(n_49), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_50), .B(n_148), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_51), .B(n_148), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_52), .B(n_446), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_53), .B(n_166), .Y(n_165) );
AOI22xp33_ASAP7_75t_SL g147 ( .A1(n_55), .A2(n_59), .B1(n_141), .B2(n_148), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_56), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_57), .B(n_148), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_58), .B(n_148), .Y(n_247) );
INVx1_ASAP7_75t_L g154 ( .A(n_60), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_61), .B(n_446), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_62), .B(n_461), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_63), .A2(n_166), .B(n_177), .C(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_64), .B(n_148), .Y(n_183) );
INVx1_ASAP7_75t_L g134 ( .A(n_65), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_66), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_67), .B(n_145), .Y(n_484) );
AO32x2_ASAP7_75t_L g204 ( .A1(n_68), .A2(n_151), .A3(n_152), .B1(n_205), .B2(n_209), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_69), .B(n_146), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_70), .A2(n_103), .B1(n_115), .B2(n_748), .Y(n_102) );
INVx1_ASAP7_75t_L g246 ( .A(n_71), .Y(n_246) );
INVx1_ASAP7_75t_L g222 ( .A(n_72), .Y(n_222) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_73), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_74), .B(n_453), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_75), .A2(n_449), .B(n_486), .C(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_76), .B(n_141), .Y(n_223) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_77), .Y(n_494) );
INVx1_ASAP7_75t_L g111 ( .A(n_78), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_79), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_81), .B(n_200), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_82), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_83), .B(n_141), .Y(n_226) );
INVx2_ASAP7_75t_L g132 ( .A(n_84), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_85), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_86), .B(n_138), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_87), .B(n_141), .Y(n_162) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_88), .B(n_108), .C(n_109), .Y(n_107) );
OR2x2_ASAP7_75t_L g433 ( .A(n_88), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g721 ( .A(n_88), .Y(n_721) );
OR2x2_ASAP7_75t_L g735 ( .A(n_88), .B(n_729), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g140 ( .A1(n_90), .A2(n_101), .B1(n_141), .B2(n_142), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_91), .B(n_446), .Y(n_479) );
INVx1_ASAP7_75t_L g483 ( .A(n_92), .Y(n_483) );
INVxp67_ASAP7_75t_L g497 ( .A(n_93), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_94), .B(n_141), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_95), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_96), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_97), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g514 ( .A(n_98), .Y(n_514) );
INVx1_ASAP7_75t_L g543 ( .A(n_99), .Y(n_543) );
AND2x2_ASAP7_75t_L g509 ( .A(n_100), .B(n_190), .Y(n_509) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx5_ASAP7_75t_SL g748 ( .A(n_105), .Y(n_748) );
AND2x2_ASAP7_75t_SL g105 ( .A(n_106), .B(n_112), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g434 ( .A(n_108), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AO221x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_730), .B1(n_733), .B2(n_742), .C(n_744), .Y(n_115) );
OAI222xp33_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_120), .B1(n_722), .B2(n_723), .C1(n_726), .C2(n_727), .Y(n_116) );
INVx1_ASAP7_75t_L g722 ( .A(n_117), .Y(n_722) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_431), .B1(n_436), .B2(n_718), .Y(n_121) );
INVx1_ASAP7_75t_L g725 ( .A(n_122), .Y(n_725) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
XNOR2xp5_ASAP7_75t_L g737 ( .A(n_124), .B(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_SL g124 ( .A(n_125), .B(n_364), .Y(n_124) );
NOR5xp2_ASAP7_75t_L g125 ( .A(n_126), .B(n_277), .C(n_323), .D(n_336), .E(n_348), .Y(n_125) );
OAI211xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_185), .B(n_231), .C(n_258), .Y(n_126) );
INVx1_ASAP7_75t_SL g359 ( .A(n_127), .Y(n_359) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_155), .Y(n_127) );
AND2x2_ASAP7_75t_L g283 ( .A(n_128), .B(n_156), .Y(n_283) );
AND2x2_ASAP7_75t_L g311 ( .A(n_128), .B(n_257), .Y(n_311) );
AND2x2_ASAP7_75t_L g319 ( .A(n_128), .B(n_262), .Y(n_319) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g249 ( .A(n_129), .B(n_157), .Y(n_249) );
INVx2_ASAP7_75t_L g261 ( .A(n_129), .Y(n_261) );
AND2x2_ASAP7_75t_L g386 ( .A(n_129), .B(n_328), .Y(n_386) );
OR2x2_ASAP7_75t_L g388 ( .A(n_129), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_136), .Y(n_129) );
INVx1_ASAP7_75t_L g255 ( .A(n_130), .Y(n_255) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_131), .Y(n_151) );
INVx1_ASAP7_75t_L g171 ( .A(n_131), .Y(n_171) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_132), .B(n_133), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
NAND3xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_150), .C(n_152), .Y(n_136) );
AO21x1_ASAP7_75t_L g254 ( .A1(n_137), .A2(n_150), .B(n_255), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_140), .B1(n_144), .B2(n_147), .Y(n_137) );
INVx2_ASAP7_75t_L g201 ( .A(n_138), .Y(n_201) );
OAI22xp5_ASAP7_75t_SL g205 ( .A1(n_138), .A2(n_146), .B1(n_206), .B2(n_208), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_138), .A2(n_144), .B1(n_213), .B2(n_214), .Y(n_212) );
INVx4_ASAP7_75t_L g469 ( .A(n_138), .Y(n_469) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx3_ASAP7_75t_L g146 ( .A(n_139), .Y(n_146) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_139), .Y(n_179) );
INVx1_ASAP7_75t_L g196 ( .A(n_139), .Y(n_196) );
AND2x2_ASAP7_75t_L g447 ( .A(n_139), .B(n_167), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_139), .Y(n_450) );
INVx2_ASAP7_75t_L g175 ( .A(n_141), .Y(n_175) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
INVx1_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_144), .A2(n_164), .B(n_165), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_L g180 ( .A1(n_144), .A2(n_181), .B(n_182), .C(n_183), .Y(n_180) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_145), .A2(n_161), .B(n_162), .Y(n_160) );
O2A1O1Ixp5_ASAP7_75t_SL g220 ( .A1(n_145), .A2(n_221), .B(n_222), .C(n_223), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_145), .A2(n_243), .B(n_244), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_145), .B(n_497), .Y(n_496) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g221 ( .A(n_148), .Y(n_221) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_148), .Y(n_545) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g200 ( .A(n_149), .Y(n_200) );
BUFx3_ASAP7_75t_L g207 ( .A(n_149), .Y(n_207) );
AND2x6_ASAP7_75t_L g449 ( .A(n_149), .B(n_450), .Y(n_449) );
INVx3_ASAP7_75t_L g461 ( .A(n_150), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_150), .B(n_488), .Y(n_487) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_150), .A2(n_513), .B(n_520), .Y(n_512) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_150), .A2(n_540), .B(n_547), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_150), .B(n_548), .Y(n_547) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_151), .A2(n_159), .B(n_168), .Y(n_158) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_151), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_151), .A2(n_525), .B(n_526), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_152), .A2(n_242), .B(n_245), .Y(n_241) );
BUFx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_153), .A2(n_160), .B(n_163), .Y(n_159) );
OAI21xp5_ASAP7_75t_L g172 ( .A1(n_153), .A2(n_173), .B(n_180), .Y(n_172) );
OAI21xp5_ASAP7_75t_L g191 ( .A1(n_153), .A2(n_192), .B(n_197), .Y(n_191) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_153), .A2(n_220), .B(n_224), .Y(n_219) );
AND2x4_ASAP7_75t_L g446 ( .A(n_153), .B(n_447), .Y(n_446) );
INVx4_ASAP7_75t_SL g471 ( .A(n_153), .Y(n_471) );
NAND2x1p5_ASAP7_75t_L g515 ( .A(n_153), .B(n_447), .Y(n_515) );
INVx2_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g299 ( .A(n_156), .B(n_271), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_156), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g413 ( .A(n_156), .B(n_253), .Y(n_413) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_169), .Y(n_156) );
AND2x2_ASAP7_75t_L g256 ( .A(n_157), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g303 ( .A(n_157), .Y(n_303) );
AND2x2_ASAP7_75t_L g328 ( .A(n_157), .B(n_240), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_157), .B(n_361), .Y(n_398) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g262 ( .A(n_158), .B(n_240), .Y(n_262) );
AND2x2_ASAP7_75t_L g276 ( .A(n_158), .B(n_239), .Y(n_276) );
AND2x2_ASAP7_75t_L g293 ( .A(n_158), .B(n_169), .Y(n_293) );
AND2x2_ASAP7_75t_L g350 ( .A(n_158), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_158), .B(n_257), .Y(n_363) );
AND2x2_ASAP7_75t_L g415 ( .A(n_158), .B(n_340), .Y(n_415) );
INVx2_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g238 ( .A(n_169), .B(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g257 ( .A(n_169), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_169), .B(n_240), .Y(n_334) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_172), .B(n_184), .Y(n_169) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_170), .A2(n_241), .B(n_248), .Y(n_240) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_171), .B(n_521), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_176), .C(n_177), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_175), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_175), .A2(n_528), .B(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_177), .A2(n_543), .B(n_544), .C(n_545), .Y(n_542) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_178), .A2(n_225), .B(n_226), .Y(n_224) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g453 ( .A(n_179), .Y(n_453) );
O2A1O1Ixp5_ASAP7_75t_L g245 ( .A1(n_181), .A2(n_201), .B(n_246), .C(n_247), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_181), .A2(n_452), .B(n_454), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_215), .B(n_228), .Y(n_185) );
INVx1_ASAP7_75t_SL g347 ( .A(n_186), .Y(n_347) );
AND2x4_ASAP7_75t_L g186 ( .A(n_187), .B(n_203), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_SL g235 ( .A(n_188), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g230 ( .A(n_189), .Y(n_230) );
INVx1_ASAP7_75t_L g267 ( .A(n_189), .Y(n_267) );
AND2x2_ASAP7_75t_L g288 ( .A(n_189), .B(n_210), .Y(n_288) );
AND2x2_ASAP7_75t_L g322 ( .A(n_189), .B(n_211), .Y(n_322) );
OR2x2_ASAP7_75t_L g341 ( .A(n_189), .B(n_217), .Y(n_341) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_189), .Y(n_355) );
AND2x2_ASAP7_75t_L g368 ( .A(n_189), .B(n_369), .Y(n_368) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_202), .Y(n_189) );
INVx2_ASAP7_75t_L g209 ( .A(n_190), .Y(n_209) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_190), .A2(n_219), .B(n_227), .Y(n_218) );
INVx1_ASAP7_75t_L g459 ( .A(n_190), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_190), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_190), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .Y(n_192) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_201), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_203), .A2(n_290), .B1(n_291), .B2(n_300), .Y(n_289) );
AND2x2_ASAP7_75t_L g373 ( .A(n_203), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_210), .Y(n_203) );
INVx1_ASAP7_75t_L g234 ( .A(n_204), .Y(n_234) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_204), .Y(n_271) );
INVx1_ASAP7_75t_L g282 ( .A(n_204), .Y(n_282) );
AND2x2_ASAP7_75t_L g297 ( .A(n_204), .B(n_211), .Y(n_297) );
INVx2_ASAP7_75t_L g470 ( .A(n_207), .Y(n_470) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_207), .Y(n_485) );
INVx1_ASAP7_75t_L g456 ( .A(n_209), .Y(n_456) );
OR2x2_ASAP7_75t_L g251 ( .A(n_210), .B(n_236), .Y(n_251) );
AND2x2_ASAP7_75t_L g281 ( .A(n_210), .B(n_282), .Y(n_281) );
NOR2xp67_ASAP7_75t_L g369 ( .A(n_210), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g229 ( .A(n_211), .B(n_230), .Y(n_229) );
BUFx2_ASAP7_75t_L g338 ( .A(n_211), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_215), .B(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g316 ( .A(n_216), .B(n_282), .Y(n_316) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g228 ( .A(n_217), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g287 ( .A(n_217), .Y(n_287) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g236 ( .A(n_218), .Y(n_236) );
OR2x2_ASAP7_75t_L g266 ( .A(n_218), .B(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_218), .Y(n_321) );
AOI32xp33_ASAP7_75t_L g358 ( .A1(n_228), .A2(n_288), .A3(n_359), .B1(n_360), .B2(n_362), .Y(n_358) );
AND2x2_ASAP7_75t_L g284 ( .A(n_229), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_229), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_229), .B(n_316), .Y(n_402) );
INVx1_ASAP7_75t_L g407 ( .A(n_229), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_237), .B1(n_250), .B2(n_252), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
AND2x2_ASAP7_75t_L g337 ( .A(n_233), .B(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_234), .B(n_236), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_235), .A2(n_259), .B1(n_263), .B2(n_273), .Y(n_258) );
AND2x2_ASAP7_75t_L g280 ( .A(n_235), .B(n_281), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_235), .A2(n_249), .B(n_297), .C(n_332), .Y(n_331) );
OAI332xp33_ASAP7_75t_L g336 ( .A1(n_235), .A2(n_337), .A3(n_339), .B1(n_341), .B2(n_342), .B3(n_344), .C1(n_345), .C2(n_347), .Y(n_336) );
INVx2_ASAP7_75t_L g377 ( .A(n_235), .Y(n_377) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_236), .Y(n_295) );
INVx1_ASAP7_75t_L g370 ( .A(n_236), .Y(n_370) );
AND2x2_ASAP7_75t_L g424 ( .A(n_236), .B(n_288), .Y(n_424) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_249), .Y(n_237) );
AND2x2_ASAP7_75t_L g304 ( .A(n_239), .B(n_254), .Y(n_304) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g253 ( .A(n_240), .B(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g352 ( .A(n_240), .B(n_254), .Y(n_352) );
INVx1_ASAP7_75t_L g361 ( .A(n_240), .Y(n_361) );
INVx1_ASAP7_75t_L g335 ( .A(n_249), .Y(n_335) );
INVxp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g419 ( .A(n_251), .B(n_271), .Y(n_419) );
INVx1_ASAP7_75t_SL g330 ( .A(n_252), .Y(n_330) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_256), .Y(n_252) );
AND2x2_ASAP7_75t_L g357 ( .A(n_253), .B(n_315), .Y(n_357) );
INVx1_ASAP7_75t_L g376 ( .A(n_253), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_253), .B(n_343), .Y(n_378) );
INVx1_ASAP7_75t_L g275 ( .A(n_254), .Y(n_275) );
AND2x2_ASAP7_75t_L g279 ( .A(n_256), .B(n_260), .Y(n_279) );
AND2x2_ASAP7_75t_L g346 ( .A(n_256), .B(n_304), .Y(n_346) );
INVx2_ASAP7_75t_L g389 ( .A(n_256), .Y(n_389) );
INVx2_ASAP7_75t_L g272 ( .A(n_257), .Y(n_272) );
AND2x2_ASAP7_75t_L g274 ( .A(n_257), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
INVx1_ASAP7_75t_L g290 ( .A(n_260), .Y(n_290) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_261), .B(n_334), .Y(n_340) );
OR2x2_ASAP7_75t_L g404 ( .A(n_261), .B(n_363), .Y(n_404) );
INVx1_ASAP7_75t_L g428 ( .A(n_261), .Y(n_428) );
INVx1_ASAP7_75t_L g384 ( .A(n_262), .Y(n_384) );
AND2x2_ASAP7_75t_L g429 ( .A(n_262), .B(n_272), .Y(n_429) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_266), .A2(n_292), .B1(n_294), .B2(n_298), .Y(n_291) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OAI322xp33_ASAP7_75t_SL g375 ( .A1(n_269), .A2(n_376), .A3(n_377), .B1(n_378), .B2(n_379), .C1(n_382), .C2(n_384), .Y(n_375) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
AND2x2_ASAP7_75t_L g372 ( .A(n_270), .B(n_288), .Y(n_372) );
OR2x2_ASAP7_75t_L g406 ( .A(n_270), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g409 ( .A(n_270), .B(n_341), .Y(n_409) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g354 ( .A(n_271), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g410 ( .A(n_271), .B(n_341), .Y(n_410) );
INVx3_ASAP7_75t_L g343 ( .A(n_272), .Y(n_343) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_L g399 ( .A(n_274), .Y(n_399) );
AOI222xp33_ASAP7_75t_L g278 ( .A1(n_276), .A2(n_279), .B1(n_280), .B2(n_283), .C1(n_284), .C2(n_286), .Y(n_278) );
INVx1_ASAP7_75t_L g309 ( .A(n_276), .Y(n_309) );
NAND3xp33_ASAP7_75t_SL g277 ( .A(n_278), .B(n_289), .C(n_306), .Y(n_277) );
AND2x2_ASAP7_75t_L g394 ( .A(n_281), .B(n_295), .Y(n_394) );
BUFx2_ASAP7_75t_L g285 ( .A(n_282), .Y(n_285) );
INVx1_ASAP7_75t_L g326 ( .A(n_282), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_283), .A2(n_319), .B1(n_372), .B2(n_373), .C(n_375), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_285), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
AND2x2_ASAP7_75t_L g325 ( .A(n_288), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_293), .B(n_304), .Y(n_305) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
OAI21xp33_ASAP7_75t_L g300 ( .A1(n_295), .A2(n_301), .B(n_305), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_295), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g392 ( .A(n_297), .B(n_374), .Y(n_392) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g315 ( .A(n_303), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_304), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g421 ( .A(n_304), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_312), .B1(n_313), .B2(n_316), .C(n_317), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_308), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g417 ( .A(n_316), .B(n_322), .Y(n_417) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
OAI31xp33_ASAP7_75t_SL g385 ( .A1(n_320), .A2(n_359), .A3(n_386), .B(n_387), .Y(n_385) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g374 ( .A(n_321), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_322), .B(n_326), .Y(n_425) );
OAI221xp5_ASAP7_75t_SL g323 ( .A1(n_324), .A2(n_327), .B1(n_329), .B2(n_330), .C(n_331), .Y(n_323) );
INVx1_ASAP7_75t_L g329 ( .A(n_325), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_328), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g344 ( .A(n_337), .Y(n_344) );
INVx2_ASAP7_75t_L g380 ( .A(n_338), .Y(n_380) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g366 ( .A(n_343), .B(n_352), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_L g416 ( .A1(n_343), .A2(n_360), .B(n_417), .C(n_418), .Y(n_416) );
OAI221xp5_ASAP7_75t_SL g348 ( .A1(n_344), .A2(n_349), .B1(n_353), .B2(n_356), .C(n_358), .Y(n_348) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
A2O1A1Ixp33_ASAP7_75t_L g411 ( .A1(n_347), .A2(n_412), .B(n_414), .C(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_350), .A2(n_401), .B1(n_403), .B2(n_405), .C(n_408), .Y(n_400) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
NOR4xp25_ASAP7_75t_L g364 ( .A(n_365), .B(n_390), .C(n_411), .D(n_422), .Y(n_364) );
OAI211xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B(n_371), .C(n_385), .Y(n_365) );
INVx1_ASAP7_75t_SL g420 ( .A(n_372), .Y(n_420) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_SL g383 ( .A(n_381), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_388), .A2(n_397), .B1(n_409), .B2(n_410), .Y(n_408) );
A2O1A1Ixp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B(n_395), .C(n_400), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI31xp33_ASAP7_75t_L g422 ( .A1(n_393), .A2(n_423), .A3(n_425), .B(n_426), .Y(n_422) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B(n_421), .Y(n_418) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_433), .A2(n_437), .B1(n_720), .B2(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g720 ( .A(n_434), .B(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g729 ( .A(n_434), .Y(n_729) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_SL g437 ( .A(n_438), .B(n_654), .Y(n_437) );
NOR5xp2_ASAP7_75t_L g438 ( .A(n_439), .B(n_585), .C(n_614), .D(n_634), .E(n_641), .Y(n_438) );
OAI211xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_473), .B(n_530), .C(n_572), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_441), .A2(n_657), .B1(n_659), .B2(n_660), .Y(n_656) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_460), .Y(n_441) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_442), .Y(n_533) );
AND2x4_ASAP7_75t_L g565 ( .A(n_442), .B(n_566), .Y(n_565) );
INVx5_ASAP7_75t_L g583 ( .A(n_442), .Y(n_583) );
AND2x2_ASAP7_75t_L g592 ( .A(n_442), .B(n_584), .Y(n_592) );
AND2x2_ASAP7_75t_L g604 ( .A(n_442), .B(n_477), .Y(n_604) );
AND2x2_ASAP7_75t_L g700 ( .A(n_442), .B(n_568), .Y(n_700) );
OR2x6_ASAP7_75t_L g442 ( .A(n_443), .B(n_457), .Y(n_442) );
AOI21xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_448), .B(n_456), .Y(n_443) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx5_ASAP7_75t_L g465 ( .A(n_449), .Y(n_465) );
INVx2_ASAP7_75t_L g455 ( .A(n_453), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_455), .A2(n_483), .B(n_484), .C(n_485), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_455), .A2(n_485), .B(n_507), .C(n_508), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx2_ASAP7_75t_L g566 ( .A(n_460), .Y(n_566) );
AND2x2_ASAP7_75t_L g584 ( .A(n_460), .B(n_539), .Y(n_584) );
AND2x2_ASAP7_75t_L g603 ( .A(n_460), .B(n_538), .Y(n_603) );
AND2x2_ASAP7_75t_L g643 ( .A(n_460), .B(n_583), .Y(n_643) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B(n_472), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_465), .B(n_466), .C(n_471), .Y(n_463) );
INVx2_ASAP7_75t_L g481 ( .A(n_465), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_465), .A2(n_471), .B(n_494), .C(n_495), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g486 ( .A(n_471), .Y(n_486) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_499), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AOI322xp5_ASAP7_75t_L g702 ( .A1(n_476), .A2(n_510), .A3(n_557), .B1(n_565), .B2(n_619), .C1(n_703), .C2(n_706), .Y(n_702) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_489), .Y(n_476) );
INVx5_ASAP7_75t_L g535 ( .A(n_477), .Y(n_535) );
AND2x2_ASAP7_75t_L g551 ( .A(n_477), .B(n_537), .Y(n_551) );
BUFx2_ASAP7_75t_L g629 ( .A(n_477), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_477), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g706 ( .A(n_477), .B(n_613), .Y(n_706) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_487), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_489), .B(n_501), .Y(n_560) );
INVx1_ASAP7_75t_L g587 ( .A(n_489), .Y(n_587) );
AND2x2_ASAP7_75t_L g600 ( .A(n_489), .B(n_522), .Y(n_600) );
AND2x2_ASAP7_75t_L g701 ( .A(n_489), .B(n_619), .Y(n_701) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g555 ( .A(n_490), .B(n_501), .Y(n_555) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_490), .Y(n_563) );
OR2x2_ASAP7_75t_L g570 ( .A(n_490), .B(n_522), .Y(n_570) );
AND2x2_ASAP7_75t_L g580 ( .A(n_490), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_490), .B(n_512), .Y(n_609) );
INVxp67_ASAP7_75t_L g633 ( .A(n_490), .Y(n_633) );
AND2x2_ASAP7_75t_L g640 ( .A(n_490), .B(n_510), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_490), .B(n_522), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_490), .B(n_511), .Y(n_666) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B(n_498), .Y(n_490) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_501), .B(n_523), .Y(n_610) );
OR2x2_ASAP7_75t_L g632 ( .A(n_501), .B(n_511), .Y(n_632) );
AND2x2_ASAP7_75t_L g645 ( .A(n_501), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_501), .B(n_600), .Y(n_651) );
OAI211xp5_ASAP7_75t_SL g655 ( .A1(n_501), .A2(n_656), .B(n_661), .C(n_670), .Y(n_655) );
AND2x2_ASAP7_75t_L g716 ( .A(n_501), .B(n_522), .Y(n_716) );
INVx5_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g569 ( .A(n_502), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_502), .B(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_502), .B(n_564), .Y(n_576) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_502), .Y(n_578) );
OR2x2_ASAP7_75t_L g589 ( .A(n_502), .B(n_511), .Y(n_589) );
AND2x2_ASAP7_75t_SL g594 ( .A(n_502), .B(n_580), .Y(n_594) );
AND2x2_ASAP7_75t_L g619 ( .A(n_502), .B(n_511), .Y(n_619) );
AND2x2_ASAP7_75t_L g639 ( .A(n_502), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g677 ( .A(n_502), .B(n_510), .Y(n_677) );
OR2x2_ASAP7_75t_L g680 ( .A(n_502), .B(n_666), .Y(n_680) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_509), .Y(n_502) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_522), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g623 ( .A1(n_511), .A2(n_624), .B(n_627), .C(n_633), .Y(n_623) );
INVx5_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_512), .B(n_522), .Y(n_554) );
AND2x2_ASAP7_75t_L g558 ( .A(n_512), .B(n_523), .Y(n_558) );
OR2x2_ASAP7_75t_L g564 ( .A(n_512), .B(n_522), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_516), .Y(n_513) );
INVx1_ASAP7_75t_SL g581 ( .A(n_522), .Y(n_581) );
OR2x2_ASAP7_75t_L g709 ( .A(n_522), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_549), .B(n_552), .C(n_561), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AOI31xp33_ASAP7_75t_L g634 ( .A1(n_532), .A2(n_635), .A3(n_637), .B(n_638), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_533), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_534), .B(n_565), .Y(n_571) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_535), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g591 ( .A(n_535), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g596 ( .A(n_535), .B(n_566), .Y(n_596) );
AND2x2_ASAP7_75t_L g606 ( .A(n_535), .B(n_565), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_535), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g626 ( .A(n_535), .B(n_583), .Y(n_626) );
AND2x2_ASAP7_75t_L g631 ( .A(n_535), .B(n_603), .Y(n_631) );
OR2x2_ASAP7_75t_L g650 ( .A(n_535), .B(n_537), .Y(n_650) );
OR2x2_ASAP7_75t_L g652 ( .A(n_535), .B(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_535), .Y(n_699) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g599 ( .A(n_537), .B(n_566), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_537), .B(n_583), .Y(n_622) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g568 ( .A(n_539), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_546), .Y(n_540) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g659 ( .A(n_551), .B(n_583), .Y(n_659) );
AOI322xp5_ASAP7_75t_L g661 ( .A1(n_551), .A2(n_565), .A3(n_603), .B1(n_662), .B2(n_663), .C1(n_664), .C2(n_667), .Y(n_661) );
INVx1_ASAP7_75t_L g669 ( .A(n_551), .Y(n_669) );
NAND2xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_556), .Y(n_552) );
INVx1_ASAP7_75t_SL g663 ( .A(n_553), .Y(n_663) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
OR2x2_ASAP7_75t_L g615 ( .A(n_554), .B(n_560), .Y(n_615) );
INVx1_ASAP7_75t_L g646 ( .A(n_554), .Y(n_646) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI32xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .A3(n_567), .B1(n_569), .B2(n_571), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
AOI21xp33_ASAP7_75t_SL g601 ( .A1(n_564), .A2(n_579), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_SL g616 ( .A(n_565), .Y(n_616) );
AND2x4_ASAP7_75t_L g613 ( .A(n_566), .B(n_583), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_566), .B(n_649), .Y(n_648) );
AOI322xp5_ASAP7_75t_L g678 ( .A1(n_567), .A2(n_594), .A3(n_613), .B1(n_646), .B2(n_679), .C1(n_681), .C2(n_682), .Y(n_678) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_567), .A2(n_644), .B1(n_708), .B2(n_709), .C(n_711), .Y(n_707) );
AND2x2_ASAP7_75t_L g595 ( .A(n_568), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_SL g575 ( .A(n_570), .Y(n_575) );
OR2x2_ASAP7_75t_L g647 ( .A(n_570), .B(n_632), .Y(n_647) );
OAI31xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_576), .A3(n_577), .B(n_582), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_573), .A2(n_606), .B1(n_607), .B2(n_611), .Y(n_605) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g618 ( .A(n_575), .B(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_577), .A2(n_618), .B1(n_671), .B2(n_674), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g660 ( .A(n_580), .B(n_629), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_580), .B(n_619), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_581), .B(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g694 ( .A(n_581), .B(n_632), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_582), .A2(n_677), .B1(n_690), .B2(n_693), .Y(n_689) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx2_ASAP7_75t_L g598 ( .A(n_583), .Y(n_598) );
AND2x2_ASAP7_75t_L g681 ( .A(n_583), .B(n_603), .Y(n_681) );
OR2x2_ASAP7_75t_L g683 ( .A(n_583), .B(n_650), .Y(n_683) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_583), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_584), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_584), .B(n_629), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_590), .B(n_593), .C(n_605), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B1(n_597), .B2(n_600), .C(n_601), .Y(n_593) );
INVxp67_ASAP7_75t_L g705 ( .A(n_596), .Y(n_705) );
INVx1_ASAP7_75t_L g672 ( .A(n_597), .Y(n_672) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g636 ( .A(n_598), .B(n_603), .Y(n_636) );
INVx1_ASAP7_75t_L g653 ( .A(n_599), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_599), .B(n_626), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g668 ( .A(n_603), .Y(n_668) );
AND2x2_ASAP7_75t_L g674 ( .A(n_603), .B(n_629), .Y(n_674) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_SL g662 ( .A(n_610), .Y(n_662) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_613), .B(n_649), .Y(n_673) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .B1(n_617), .B2(n_620), .C(n_623), .Y(n_614) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g710 ( .A(n_619), .Y(n_710) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g628 ( .A(n_622), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_626), .B(n_685), .Y(n_684) );
AOI21xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_630), .B(n_632), .Y(n_627) );
OAI211xp5_ASAP7_75t_SL g675 ( .A1(n_630), .A2(n_676), .B(n_678), .C(n_684), .Y(n_675) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g687 ( .A(n_632), .Y(n_687) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI222xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_644), .B1(n_647), .B2(n_648), .C1(n_651), .C2(n_652), .Y(n_641) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g717 ( .A(n_648), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_649), .B(n_692), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_649), .A2(n_696), .B1(n_698), .B2(n_701), .Y(n_695) );
INVx2_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
NOR4xp25_ASAP7_75t_L g654 ( .A(n_655), .B(n_675), .C(n_688), .D(n_707), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_657), .B(n_687), .Y(n_697) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g664 ( .A(n_662), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_665), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_695), .C(n_702), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx2_ASAP7_75t_L g704 ( .A(n_700), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
OAI21xp5_ASAP7_75t_SL g711 ( .A1(n_712), .A2(n_714), .B(n_717), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NOR2x2_ASAP7_75t_L g728 ( .A(n_721), .B(n_729), .Y(n_728) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
BUFx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_SL g743 ( .A(n_731), .Y(n_743) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g747 ( .A(n_735), .Y(n_747) );
INVx1_ASAP7_75t_L g740 ( .A(n_737), .Y(n_740) );
BUFx3_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
endmodule