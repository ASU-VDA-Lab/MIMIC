module fake_aes_2459_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx1_ASAP7_75t_L g11 ( .A(n_7), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_5), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_9), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_8), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_3), .B(n_6), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_2), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
NOR3xp33_ASAP7_75t_SL g19 ( .A(n_13), .B(n_0), .C(n_1), .Y(n_19) );
INVx5_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_16), .B(n_0), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_11), .Y(n_22) );
AND2x4_ASAP7_75t_L g23 ( .A(n_21), .B(n_14), .Y(n_23) );
AOI22xp33_ASAP7_75t_SL g24 ( .A1(n_21), .A2(n_12), .B1(n_15), .B2(n_1), .Y(n_24) );
AND2x4_ASAP7_75t_L g25 ( .A(n_20), .B(n_2), .Y(n_25) );
INVx4_ASAP7_75t_L g26 ( .A(n_20), .Y(n_26) );
NAND2xp33_ASAP7_75t_R g27 ( .A(n_23), .B(n_19), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_24), .B(n_18), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_23), .Y(n_31) );
INVxp67_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_30), .Y(n_33) );
AOI21xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_25), .B(n_20), .Y(n_34) );
OAI21xp33_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_19), .B(n_22), .Y(n_35) );
AOI21xp5_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_26), .B(n_18), .Y(n_36) );
NAND2xp5_ASAP7_75t_SL g37 ( .A(n_35), .B(n_27), .Y(n_37) );
CKINVDCx20_ASAP7_75t_R g38 ( .A(n_37), .Y(n_38) );
AOI22xp33_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_36), .B1(n_27), .B2(n_10), .Y(n_39) );
endmodule