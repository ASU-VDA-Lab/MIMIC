module fake_jpeg_22646_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_49),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_28),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_51),
.B(n_18),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_56),
.Y(n_95)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

INVx5_ASAP7_75t_SL g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_61),
.Y(n_85)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_35),
.B1(n_22),
.B2(n_30),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_42),
.B1(n_31),
.B2(n_17),
.Y(n_91)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_67),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_28),
.B(n_29),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_26),
.C(n_24),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_17),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_31),
.C(n_27),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_35),
.B1(n_29),
.B2(n_19),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_65),
.A2(n_73),
.B1(n_79),
.B2(n_81),
.Y(n_116)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_22),
.B1(n_18),
.B2(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_24),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_17),
.Y(n_97)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_32),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_22),
.B1(n_18),
.B2(n_25),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_31),
.Y(n_83)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_86),
.B(n_89),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_48),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_110),
.B1(n_59),
.B2(n_72),
.Y(n_125)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_94),
.Y(n_141)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_93),
.B(n_102),
.CI(n_38),
.CON(n_134),
.SN(n_134)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_96),
.B(n_99),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_105),
.Y(n_146)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_74),
.B(n_19),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_100),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_101),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_64),
.B(n_17),
.CI(n_36),
.CON(n_102),
.SN(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_103),
.B(n_107),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_36),
.B1(n_49),
.B2(n_37),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_60),
.B1(n_62),
.B2(n_53),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_19),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_53),
.A2(n_26),
.B1(n_24),
.B2(n_29),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_119),
.B1(n_20),
.B2(n_23),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_34),
.C(n_33),
.Y(n_127)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_33),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_122),
.A2(n_129),
.B(n_146),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_86),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_132),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_143),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_69),
.B1(n_68),
.B2(n_61),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_127),
.B(n_11),
.C(n_1),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_71),
.B1(n_67),
.B2(n_76),
.Y(n_128)
);

NAND2xp33_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_0),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_137),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_89),
.A2(n_48),
.A3(n_38),
.B1(n_20),
.B2(n_23),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_38),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_133),
.B(n_136),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_134),
.B(n_85),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_13),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_95),
.A2(n_37),
.B1(n_27),
.B2(n_34),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_147),
.B1(n_156),
.B2(n_117),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_20),
.A3(n_38),
.B1(n_23),
.B2(n_12),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_88),
.Y(n_158)
);

AOI22x1_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_20),
.B1(n_23),
.B2(n_2),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_144),
.B(n_149),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_121),
.A2(n_32),
.B1(n_37),
.B2(n_27),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_91),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_148),
.A2(n_150),
.B1(n_152),
.B2(n_119),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_90),
.B(n_14),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_92),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_96),
.A2(n_12),
.B1(n_11),
.B2(n_8),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_99),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_158),
.A2(n_166),
.B1(n_1),
.B2(n_2),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_111),
.B(n_113),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_129),
.B(n_127),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_155),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_161),
.B(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_169),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_98),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_178),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_164),
.A2(n_191),
.B(n_169),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_168),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_173),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_172),
.A2(n_184),
.B1(n_3),
.B2(n_4),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_106),
.Y(n_177)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_124),
.B(n_115),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_104),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_180),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_106),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_155),
.B(n_8),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_131),
.B(n_94),
.Y(n_183)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_122),
.A2(n_117),
.B1(n_114),
.B2(n_101),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_187),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_147),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_191),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_7),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_0),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_134),
.B1(n_142),
.B2(n_132),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_196),
.B1(n_202),
.B2(n_203),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_217),
.B(n_181),
.Y(n_226)
);

AO22x1_ASAP7_75t_SL g195 ( 
.A1(n_167),
.A2(n_134),
.B1(n_136),
.B2(n_109),
.Y(n_195)
);

AO22x1_ASAP7_75t_SL g232 ( 
.A1(n_195),
.A2(n_186),
.B1(n_160),
.B2(n_172),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_135),
.B1(n_123),
.B2(n_140),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_11),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_219),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_165),
.A2(n_135),
.B1(n_123),
.B2(n_154),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_189),
.A2(n_154),
.B1(n_138),
.B2(n_137),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_138),
.B1(n_112),
.B2(n_108),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_207),
.B1(n_215),
.B2(n_220),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_3),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_177),
.B(n_174),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_200),
.B1(n_159),
.B2(n_209),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_185),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_164),
.A2(n_6),
.B(n_7),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_221),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_171),
.A2(n_7),
.B1(n_174),
.B2(n_167),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_162),
.Y(n_227)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_225),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_242),
.B(n_213),
.Y(n_250)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

AO21x1_ASAP7_75t_L g267 ( 
.A1(n_226),
.A2(n_232),
.B(n_159),
.Y(n_267)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_178),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_234),
.C(n_237),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_194),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_230),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_195),
.A2(n_166),
.B1(n_186),
.B2(n_170),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_231),
.A2(n_210),
.B1(n_184),
.B2(n_199),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_201),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_179),
.Y(n_236)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_201),
.C(n_186),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_203),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_238),
.B(n_239),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_211),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_209),
.A2(n_161),
.B(n_168),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_190),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_217),
.Y(n_257)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_233),
.B1(n_235),
.B2(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_242),
.C(n_226),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_195),
.B1(n_196),
.B2(n_222),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_252),
.A2(n_254),
.B1(n_256),
.B2(n_265),
.Y(n_272)
);

AOI22x1_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_192),
.B1(n_210),
.B2(n_215),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_213),
.B(n_193),
.C(n_175),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_263),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_267),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_234),
.B(n_219),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_212),
.B1(n_216),
.B2(n_176),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_231),
.B(n_176),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_240),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_225),
.Y(n_268)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_270),
.A2(n_188),
.B(n_182),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_237),
.C(n_229),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_279),
.C(n_284),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_253),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_282),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_223),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_283),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_243),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_281),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_228),
.B1(n_227),
.B2(n_236),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_256),
.B1(n_257),
.B2(n_261),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_224),
.C(n_240),
.Y(n_279)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_259),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_216),
.C(n_182),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_188),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_282),
.B1(n_269),
.B2(n_264),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_275),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_298),
.Y(n_303)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_272),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_250),
.B(n_255),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_295),
.Y(n_305)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_255),
.C(n_260),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_267),
.B(n_252),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_280),
.Y(n_300)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_270),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_307),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_281),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_299),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_306),
.A2(n_293),
.B1(n_289),
.B2(n_290),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_316),
.B(n_302),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_305),
.B(n_291),
.Y(n_311)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_295),
.C(n_292),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_317),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_318),
.Y(n_324)
);

NOR2x1_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_308),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_320),
.C(n_312),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_309),
.B(n_301),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_314),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_325),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_324),
.A2(n_321),
.B(n_319),
.Y(n_327)
);

AOI321xp33_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_326),
.A3(n_310),
.B1(n_300),
.B2(n_303),
.C(n_298),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_292),
.B(n_279),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_286),
.B(n_294),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_294),
.B1(n_278),
.B2(n_182),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_278),
.Y(n_332)
);


endmodule