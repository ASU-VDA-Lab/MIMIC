module fake_jpeg_17723_n_209 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_209);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_43),
.Y(n_65)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_45),
.B(n_52),
.Y(n_78)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_62),
.Y(n_100)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_5),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_59),
.Y(n_67)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

CKINVDCx6p67_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx6p67_ASAP7_75t_R g99 ( 
.A(n_56),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_92)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_63),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_10),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_31),
.C(n_37),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_76),
.Y(n_106)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_36),
.Y(n_71)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_25),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_35),
.B(n_27),
.C(n_23),
.Y(n_77)
);

NOR2x1_ASAP7_75t_R g131 ( 
.A(n_77),
.B(n_64),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_32),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_0),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_60),
.A2(n_38),
.B1(n_20),
.B2(n_29),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_92),
.B1(n_96),
.B2(n_12),
.Y(n_113)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_35),
.B1(n_23),
.B2(n_27),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_4),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_46),
.A2(n_32),
.B1(n_37),
.B2(n_31),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_12),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_16),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_16),
.Y(n_93)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_5),
.B1(n_2),
.B2(n_3),
.Y(n_96)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_41),
.B(n_16),
.Y(n_98)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_119),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_3),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_68),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_72),
.B1(n_66),
.B2(n_82),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_78),
.B(n_4),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_120),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_SL g146 ( 
.A(n_113),
.B(n_121),
.C(n_131),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_13),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_98),
.B(n_73),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_70),
.B(n_65),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_126),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_124),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_74),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_100),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_67),
.B(n_74),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_127),
.B(n_130),
.Y(n_156)
);

INVxp67_ASAP7_75t_SL g129 ( 
.A(n_89),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_92),
.B(n_88),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_125),
.B1(n_102),
.B2(n_128),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_95),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_91),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_115),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_121),
.B(n_119),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_87),
.B(n_99),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_91),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_84),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_107),
.B(n_123),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_113),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_165),
.C(n_166),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_153),
.A2(n_110),
.B1(n_86),
.B2(n_97),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_169),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_110),
.B1(n_128),
.B2(n_102),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_87),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_175),
.C(n_140),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_86),
.B1(n_117),
.B2(n_75),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_132),
.A2(n_117),
.B1(n_99),
.B2(n_87),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_171),
.A2(n_157),
.B(n_144),
.C(n_151),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_116),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_135),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_87),
.B1(n_99),
.B2(n_124),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_172),
.B1(n_158),
.B2(n_174),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_156),
.C(n_146),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_177),
.B(n_185),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_135),
.C(n_140),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_160),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_167),
.B(n_135),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_183),
.B1(n_170),
.B2(n_149),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_136),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_175),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_R g185 ( 
.A(n_168),
.B(n_134),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_186),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_191),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_194),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_159),
.B(n_162),
.C(n_166),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_176),
.C(n_177),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_176),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_199),
.Y(n_202)
);

AOI31xp67_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_191),
.A3(n_192),
.B(n_187),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_189),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_201),
.B(n_138),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_181),
.C(n_154),
.Y(n_206)
);

NAND4xp25_ASAP7_75t_SL g205 ( 
.A(n_203),
.B(n_133),
.C(n_152),
.D(n_143),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_205),
.B(n_206),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_154),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_202),
.Y(n_209)
);


endmodule