module real_jpeg_22790_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_267;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_0),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_0),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_0),
.B(n_71),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_0),
.B(n_54),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_0),
.B(n_59),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_0),
.B(n_28),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_0),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_0),
.B(n_45),
.Y(n_239)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_5),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_5),
.B(n_45),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_5),
.B(n_68),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_5),
.B(n_71),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_5),
.B(n_28),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_5),
.B(n_59),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_5),
.B(n_201),
.Y(n_200)
);

INVx8_ASAP7_75t_SL g52 ( 
.A(n_6),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_7),
.B(n_59),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_7),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_7),
.B(n_45),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_7),
.B(n_28),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_7),
.B(n_17),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_9),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_9),
.B(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_9),
.B(n_54),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_9),
.B(n_17),
.Y(n_144)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_11),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_11),
.B(n_50),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_11),
.B(n_54),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_11),
.B(n_59),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_11),
.B(n_71),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_11),
.B(n_28),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_11),
.B(n_17),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_12),
.B(n_54),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_12),
.B(n_45),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_12),
.B(n_71),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_12),
.B(n_28),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_12),
.B(n_50),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_13),
.B(n_28),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_13),
.B(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_15),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_15),
.B(n_71),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_71),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_16),
.B(n_54),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_16),
.B(n_59),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_16),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_16),
.B(n_28),
.Y(n_187)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_17),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_157),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_134),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_56),
.C(n_63),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_22),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.C(n_48),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_23),
.B(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_25),
.B(n_30),
.C(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_27),
.B(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_40),
.A2(n_41),
.B(n_44),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_40),
.B(n_48),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_43),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.C(n_55),
.Y(n_48)
);

FAx1_ASAP7_75t_SL g138 ( 
.A(n_49),
.B(n_53),
.CI(n_55),
.CON(n_138),
.SN(n_138)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_51),
.B(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_56),
.B(n_63),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_61),
.C(n_62),
.Y(n_123)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_59),
.Y(n_220)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_73),
.C(n_75),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_64),
.B(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.C(n_70),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_65),
.B(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_66),
.B(n_220),
.Y(n_219)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_69),
.B(n_70),
.Y(n_256)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_100),
.B2(n_133),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_90),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_85),
.B(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_86),
.A2(n_88),
.B1(n_92),
.B2(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_87),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_92),
.C(n_93),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_92),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_94),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_96),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.CI(n_99),
.CON(n_96),
.SN(n_96)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_122),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_112),
.C(n_118),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_107),
.C(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_108),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_118),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.C(n_116),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_132),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_128),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_153),
.C(n_155),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_135),
.A2(n_136),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_149),
.C(n_151),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_137),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.C(n_145),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_138),
.B(n_249),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_138),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_139),
.A2(n_140),
.B1(n_145),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_145),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.C(n_148),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_146),
.B(n_147),
.CI(n_148),
.CON(n_235),
.SN(n_235)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_149),
.B(n_151),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_153),
.B(n_155),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_269),
.C(n_270),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_259),
.C(n_260),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_242),
.C(n_243),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_229),
.C(n_230),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_191),
.C(n_203),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_176),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_171),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_164),
.B(n_171),
.C(n_176),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_169),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_166),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_172),
.B(n_174),
.C(n_175),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_184),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_177),
.B(n_185),
.C(n_186),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_182),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_178),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_202)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_188),
.B(n_190),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.C(n_202),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_196),
.B1(n_202),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_207)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_225),
.C(n_226),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_212),
.C(n_217),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_210),
.C(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.C(n_221),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_237),
.C(n_241),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_234),
.C(n_235),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_235),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_237),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.CI(n_240),
.CON(n_237),
.SN(n_237)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_251),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_247),
.C(n_251),
.Y(n_259)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_255),
.C(n_257),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_254),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_255),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_268),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_265),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);


endmodule