module real_jpeg_5958_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_1),
.A2(n_83),
.B1(n_86),
.B2(n_89),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_1),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_1),
.A2(n_89),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_1),
.A2(n_89),
.B1(n_206),
.B2(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_1),
.A2(n_89),
.B1(n_269),
.B2(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_2),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_2),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_2),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_114),
.B1(n_116),
.B2(n_119),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_3),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_3),
.A2(n_119),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_5),
.Y(n_157)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_5),
.Y(n_170)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_5),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_5),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_5),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_5),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_6),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_6),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_9),
.A2(n_49),
.B1(n_244),
.B2(n_247),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_9),
.B(n_259),
.C(n_261),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_9),
.B(n_74),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_9),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_9),
.B(n_98),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_9),
.B(n_337),
.Y(n_336)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_10),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_10),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_10),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_11),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_11),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_11),
.A2(n_94),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_11),
.A2(n_94),
.B1(n_255),
.B2(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_12),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_12),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_165),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_13),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_14),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_14),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_14),
.A2(n_168),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_15),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_15),
.A2(n_58),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_15),
.A2(n_58),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_15),
.A2(n_58),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_235),
.B1(n_236),
.B2(n_376),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_18),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_234),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_196),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_20),
.B(n_196),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_135),
.C(n_176),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_21),
.B(n_373),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_62),
.B2(n_134),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_22),
.B(n_63),
.C(n_96),
.Y(n_215)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_46),
.B(n_55),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_24),
.B(n_57),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_32),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_SL g147 ( 
.A(n_28),
.Y(n_147)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_40),
.B2(n_44),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_35),
.Y(n_149)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_39),
.Y(n_182)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_43),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_43),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_49),
.B(n_50),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_49),
.B(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_49),
.A2(n_155),
.B(n_272),
.Y(n_298)
);

OAI21xp33_ASAP7_75t_SL g331 ( 
.A1(n_49),
.A2(n_332),
.B(n_335),
.Y(n_331)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_50),
.A2(n_139),
.A3(n_142),
.B1(n_146),
.B2(n_148),
.Y(n_138)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_61),
.Y(n_195)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_96),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_82),
.B1(n_90),
.B2(n_91),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_64),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_74),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_70),
.Y(n_350)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_70),
.Y(n_357)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_74)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_77),
.Y(n_206)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_77),
.Y(n_257)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_77),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_77),
.Y(n_328)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_79),
.Y(n_246)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_79),
.Y(n_250)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_82),
.A2(n_90),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_85),
.Y(n_334)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_90),
.B(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_91),
.Y(n_232)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_92),
.Y(n_183)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g344 ( 
.A1(n_95),
.A2(n_336),
.A3(n_345),
.B1(n_347),
.B2(n_351),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_113),
.B(n_120),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_97),
.A2(n_113),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_97),
.A2(n_200),
.B1(n_282),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_98),
.B(n_121),
.Y(n_251)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_99),
.A2(n_120),
.B(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_107),
.B2(n_110),
.Y(n_99)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_105),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_105),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_112),
.Y(n_260)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_127),
.B1(n_130),
.B2(n_133),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_125),
.Y(n_200)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_135),
.A2(n_136),
.B1(n_176),
.B2(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_153),
.B2(n_154),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_138),
.B(n_153),
.Y(n_219)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_163),
.B1(n_169),
.B2(n_171),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_155),
.A2(n_265),
.B(n_272),
.Y(n_264)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_156),
.A2(n_164),
.B1(n_186),
.B2(n_190),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_156),
.A2(n_172),
.B1(n_208),
.B2(n_213),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_156),
.B(n_275),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_156),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_162),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_162),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_SL g278 ( 
.A(n_166),
.Y(n_278)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_174),
.Y(n_267)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_176),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_185),
.C(n_194),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_177),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_184),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_184),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_184),
.A2(n_233),
.B(n_331),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_185),
.B(n_194),
.Y(n_367)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_186),
.Y(n_341)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_189),
.Y(n_276)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_193),
.Y(n_297)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_193),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_223),
.B(n_229),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_218),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_197)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_207),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_200),
.A2(n_243),
.B(n_251),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_200),
.A2(n_251),
.B(n_327),
.Y(n_364)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_230),
.B2(n_231),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AOI21x1_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_370),
.B(n_375),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_359),
.B(n_369),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_321),
.B(n_358),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_288),
.B(n_320),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_263),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_241),
.B(n_263),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_252),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_242),
.A2(n_252),
.B1(n_253),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_242),
.Y(n_318)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_250),
.Y(n_346)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_250),
.Y(n_354)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_279),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_264),
.B(n_280),
.C(n_287),
.Y(n_322)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_286),
.B2(n_287),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_311),
.B(n_319),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_299),
.B(n_310),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_298),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_296),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_309),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_309),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_305),
.B(n_308),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_307),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_308),
.A2(n_341),
.B(n_342),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_317),
.Y(n_319)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_323),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_339),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_329),
.B2(n_330),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_329),
.C(n_339),
.Y(n_360)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_344),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_340),
.B(n_344),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_355),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_360),
.B(n_361),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_366),
.B2(n_368),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_364),
.B(n_365),
.C(n_368),
.Y(n_371)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_366),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_371),
.B(n_372),
.Y(n_375)
);


endmodule