module fake_jpeg_14595_n_348 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_38),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_8),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_41),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

HAxp5_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_0),
.CON(n_43),
.SN(n_43)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_26),
.B(n_29),
.C(n_32),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_50),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_20),
.B1(n_27),
.B2(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_66),
.C(n_68),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_22),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_60),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_28),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_28),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_20),
.B1(n_27),
.B2(n_29),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_18),
.B1(n_32),
.B2(n_21),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_42),
.B1(n_21),
.B2(n_18),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_19),
.B1(n_24),
.B2(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_36),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_59),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_86),
.C(n_90),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_34),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_34),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_99),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_53),
.B(n_56),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_47),
.B(n_36),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_63),
.B(n_65),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_58),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_40),
.B(n_19),
.C(n_41),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_70),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_72),
.Y(n_97)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_64),
.B(n_40),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_100),
.A2(n_75),
.B(n_85),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_42),
.B1(n_54),
.B2(n_45),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_101),
.A2(n_111),
.B1(n_115),
.B2(n_117),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_110),
.Y(n_135)
);

BUFx24_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_112),
.B(n_118),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_54),
.B1(n_45),
.B2(n_71),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_63),
.B(n_48),
.C(n_40),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_78),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_124),
.B1(n_97),
.B2(n_89),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_84),
.A2(n_54),
.B1(n_45),
.B2(n_41),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_33),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_126),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_73),
.A2(n_45),
.B1(n_41),
.B2(n_52),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_97),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_37),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_88),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_91),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_73),
.B(n_76),
.Y(n_141)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_78),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_77),
.A2(n_16),
.B1(n_24),
.B2(n_23),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_88),
.B1(n_73),
.B2(n_98),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_33),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_128),
.B(n_130),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_121),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_142),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_90),
.B1(n_86),
.B2(n_79),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_146),
.B(n_147),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_150),
.B1(n_119),
.B2(n_48),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_39),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_94),
.C(n_92),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_153),
.C(n_117),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_127),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_103),
.A2(n_81),
.B(n_79),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_94),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_110),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_103),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_149),
.A2(n_152),
.B(n_156),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_81),
.B1(n_94),
.B2(n_76),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

NOR2x1_ASAP7_75t_R g152 ( 
.A(n_109),
.B(n_76),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_75),
.C(n_39),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_107),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_162),
.C(n_168),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_156),
.A2(n_118),
.B1(n_112),
.B2(n_102),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_184),
.B1(n_131),
.B2(n_155),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_122),
.B1(n_105),
.B2(n_101),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_160),
.A2(n_181),
.B1(n_146),
.B2(n_114),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_179),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_115),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_143),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_140),
.A2(n_141),
.B(n_152),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_167),
.A2(n_143),
.B(n_137),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_39),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_93),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_169),
.B(n_137),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_135),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_170),
.B(n_180),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_108),
.Y(n_173)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_143),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_128),
.A2(n_124),
.B1(n_114),
.B2(n_48),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_148),
.A2(n_139),
.B1(n_145),
.B2(n_134),
.Y(n_184)
);

NOR2x1_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_153),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_185),
.A2(n_194),
.B1(n_203),
.B2(n_211),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_145),
.C(n_130),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_168),
.C(n_163),
.Y(n_225)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_198),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_177),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_209),
.B1(n_212),
.B2(n_0),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_200),
.B(n_33),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_202),
.B(n_205),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_159),
.A2(n_124),
.B1(n_129),
.B2(n_85),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_204),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_165),
.B(n_129),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_151),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_39),
.Y(n_236)
);

AO22x2_ASAP7_75t_L g207 ( 
.A1(n_159),
.A2(n_106),
.B1(n_78),
.B2(n_62),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_208),
.B1(n_39),
.B2(n_25),
.Y(n_237)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_93),
.B(n_74),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_210),
.A2(n_183),
.B(n_172),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_171),
.A2(n_55),
.B1(n_57),
.B2(n_106),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_201),
.A2(n_160),
.B1(n_184),
.B2(n_173),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_197),
.A2(n_185),
.B1(n_191),
.B2(n_210),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_220),
.B(n_224),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_238),
.Y(n_246)
);

OAI22x1_ASAP7_75t_SL g223 ( 
.A1(n_207),
.A2(n_162),
.B1(n_172),
.B2(n_161),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_223),
.A2(n_237),
.B1(n_207),
.B2(n_195),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_166),
.B1(n_167),
.B2(n_179),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_227),
.C(n_229),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_163),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_228),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_106),
.C(n_62),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_46),
.C(n_37),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_46),
.C(n_37),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_233),
.C(n_234),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_194),
.C(n_200),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_46),
.C(n_37),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_37),
.C(n_39),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_239),
.C(n_31),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_30),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_212),
.A2(n_16),
.B1(n_23),
.B2(n_24),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_211),
.B(n_30),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_193),
.Y(n_247)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_247),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_214),
.B1(n_16),
.B2(n_3),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_214),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_251),
.B(n_252),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_216),
.B(n_193),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_207),
.B1(n_188),
.B2(n_203),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_253),
.A2(n_255),
.B1(n_261),
.B2(n_235),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_258),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_233),
.A2(n_25),
.B1(n_31),
.B2(n_24),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_0),
.Y(n_256)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_222),
.B(n_11),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_257),
.B(n_10),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_1),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_0),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_213),
.A2(n_31),
.B1(n_16),
.B2(n_23),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_30),
.C(n_31),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_225),
.C(n_227),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_279),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_271),
.C(n_278),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_248),
.B1(n_250),
.B2(n_244),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_253),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_231),
.C(n_229),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_245),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_221),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_276),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_228),
.C(n_239),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_273),
.B(n_256),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_261),
.B1(n_2),
.B2(n_3),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_9),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_281),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_276),
.B(n_249),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_296),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_290),
.C(n_297),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_4),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_245),
.C(n_262),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_246),
.B1(n_254),
.B2(n_241),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_292),
.A2(n_294),
.B1(n_5),
.B2(n_6),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_9),
.B(n_15),
.Y(n_295)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_7),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_1),
.C(n_2),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_1),
.C(n_3),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_5),
.C(n_6),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_263),
.A2(n_11),
.B(n_14),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_7),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_266),
.B(n_277),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_303),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_282),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_302),
.B(n_308),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_11),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_288),
.A2(n_274),
.B(n_12),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_294),
.B1(n_5),
.B2(n_12),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_10),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_307),
.Y(n_320)
);

XNOR2x1_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_5),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_297),
.B(n_298),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_312),
.B(n_313),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_322),
.Y(n_334)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_318),
.B(n_321),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_283),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_283),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_309),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_325),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_10),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_12),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_13),
.B(n_14),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_316),
.A2(n_310),
.B1(n_314),
.B2(n_306),
.Y(n_327)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_327),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_331),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_307),
.B(n_35),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_35),
.C(n_330),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_320),
.A2(n_35),
.B(n_315),
.C(n_323),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_332),
.A2(n_333),
.B(n_35),
.Y(n_338)
);

O2A1O1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_320),
.A2(n_35),
.B(n_321),
.C(n_316),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_336),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_337),
.A2(n_335),
.B(n_35),
.Y(n_344)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_338),
.A2(n_339),
.B(n_341),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_35),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_344),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_340),
.C(n_342),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_343),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_336),
.Y(n_348)
);


endmodule