module fake_jpeg_12941_n_286 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_83),
.Y(n_105)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_54),
.B(n_58),
.Y(n_102)
);

BUFx12f_ASAP7_75t_SL g55 ( 
.A(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_77),
.Y(n_100)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_3),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx5_ASAP7_75t_SL g116 ( 
.A(n_59),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_60),
.Y(n_90)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_26),
.B(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_63),
.B(n_78),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_23),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_68),
.A2(n_38),
.B1(n_42),
.B2(n_45),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_26),
.B(n_15),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_28),
.B(n_5),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_85),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_17),
.B(n_30),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_40),
.Y(n_117)
);

HAxp5_ASAP7_75t_SL g85 ( 
.A(n_38),
.B(n_6),
.CON(n_85),
.SN(n_85)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_88),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_54),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_111),
.B(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_58),
.B(n_44),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_9),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_44),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_17),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_43),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_43),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_75),
.A2(n_40),
.B1(n_45),
.B2(n_24),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_130),
.B1(n_132),
.B2(n_87),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_59),
.B1(n_7),
.B2(n_8),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_42),
.B1(n_37),
.B2(n_30),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_37),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_24),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_81),
.A2(n_84),
.B1(n_57),
.B2(n_67),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_137),
.B(n_153),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_145),
.Y(n_168)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_47),
.B1(n_46),
.B2(n_60),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_160),
.B1(n_97),
.B2(n_118),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_149),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_150),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_161),
.B1(n_92),
.B2(n_133),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_6),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_151),
.B(n_155),
.Y(n_183)
);

NAND2x1_ASAP7_75t_L g152 ( 
.A(n_93),
.B(n_7),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_156),
.C(n_166),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_15),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_12),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_101),
.A2(n_13),
.B(n_14),
.C(n_126),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_162),
.B(n_91),
.Y(n_190)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_109),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_163),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_14),
.B1(n_103),
.B2(n_121),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_102),
.A2(n_14),
.B1(n_130),
.B2(n_114),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_118),
.A2(n_94),
.B1(n_97),
.B2(n_95),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_92),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_95),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_165),
.Y(n_178)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_100),
.B(n_128),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_159),
.A2(n_123),
.B1(n_121),
.B2(n_96),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_185),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_96),
.B1(n_133),
.B2(n_114),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_190),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_165),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_160),
.A2(n_106),
.B1(n_89),
.B2(n_120),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_89),
.B1(n_120),
.B2(n_98),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_134),
.B1(n_145),
.B2(n_144),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_91),
.B1(n_98),
.B2(n_137),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_191),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_149),
.A2(n_147),
.B1(n_166),
.B2(n_155),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_181),
.B(n_155),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_183),
.C(n_171),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_188),
.A2(n_134),
.B1(n_145),
.B2(n_144),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_200),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_169),
.B(n_187),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_198),
.B(n_203),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_169),
.B(n_138),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_187),
.B(n_140),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_211),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_181),
.A2(n_146),
.B(n_135),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_183),
.B(n_152),
.Y(n_215)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_170),
.B(n_136),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_152),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_227),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_223),
.C(n_228),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_189),
.C(n_168),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_201),
.A2(n_204),
.B1(n_211),
.B2(n_182),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_204),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_175),
.B1(n_177),
.B2(n_185),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_226),
.A2(n_200),
.B1(n_197),
.B2(n_202),
.Y(n_242)
);

AOI221xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_190),
.B1(n_168),
.B2(n_179),
.C(n_174),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_184),
.C(n_179),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_228),
.A2(n_209),
.B(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_213),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_238),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_209),
.C(n_207),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_245),
.C(n_215),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_241),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_244),
.B1(n_224),
.B2(n_217),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_225),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_231),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_249),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_232),
.B(n_237),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_241),
.A2(n_226),
.B1(n_220),
.B2(n_227),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_253),
.A2(n_256),
.B1(n_242),
.B2(n_244),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_230),
.C(n_224),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_239),
.C(n_233),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_243),
.A2(n_221),
.B1(n_196),
.B2(n_195),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_256),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_261),
.C(n_263),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_252),
.C(n_246),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_265),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_233),
.C(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_235),
.C(n_229),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_266),
.C(n_249),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_221),
.B1(n_176),
.B2(n_158),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_270),
.B(n_253),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_248),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_250),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_248),
.B(n_255),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_262),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_274),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_250),
.B(n_268),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_275),
.A2(n_176),
.B1(n_173),
.B2(n_154),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_276),
.B(n_271),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_173),
.C(n_167),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_278),
.C(n_167),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_281),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_282),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_283),
.B(n_141),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_164),
.Y(n_286)
);


endmodule