module fake_jpeg_24772_n_306 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_155;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_0),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_28),
.Y(n_73)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_24),
.B1(n_18),
.B2(n_29),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_53),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_24),
.B1(n_18),
.B2(n_29),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_54),
.A2(n_55),
.B1(n_71),
.B2(n_75),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_18),
.B1(n_29),
.B2(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_63),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_66),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_34),
.B1(n_38),
.B2(n_23),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_72),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_34),
.B1(n_38),
.B2(n_23),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_34),
.B1(n_25),
.B2(n_33),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_25),
.B1(n_33),
.B2(n_35),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_77),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_28),
.B1(n_35),
.B2(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_31),
.Y(n_100)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_79),
.B(n_83),
.Y(n_128)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_84),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_49),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_85),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_88),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_44),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_87),
.B(n_105),
.Y(n_141)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_49),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_2),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_52),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_90),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_93),
.B(n_97),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_37),
.B(n_45),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_94),
.B(n_21),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_32),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_104),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_73),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_31),
.B1(n_22),
.B2(n_30),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_77),
.B1(n_57),
.B2(n_72),
.Y(n_124)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx5_ASAP7_75t_SL g118 ( 
.A(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_37),
.Y(n_104)
);

AND2x6_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_1),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_37),
.C(n_22),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_114),
.C(n_21),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_54),
.A2(n_22),
.B1(n_30),
.B2(n_27),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

BUFx16f_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

BUFx16f_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_62),
.B(n_1),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_37),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_115),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_37),
.C(n_30),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_27),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_50),
.A2(n_27),
.B1(n_21),
.B2(n_4),
.Y(n_116)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_109),
.B1(n_114),
.B2(n_102),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_137),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_60),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_142),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_143),
.Y(n_164)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_112),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_79),
.B(n_60),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_144),
.A2(n_146),
.B(n_147),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_96),
.A2(n_57),
.B1(n_74),
.B2(n_50),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_145),
.A2(n_116),
.B1(n_94),
.B2(n_107),
.Y(n_150)
);

NAND2x1_ASAP7_75t_SL g147 ( 
.A(n_89),
.B(n_50),
.Y(n_147)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_111),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_155),
.B1(n_156),
.B2(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_83),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_153),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_84),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_109),
.B1(n_97),
.B2(n_105),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_157),
.B(n_160),
.Y(n_197)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_120),
.B(n_93),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_173),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_57),
.B1(n_106),
.B2(n_104),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_113),
.CI(n_100),
.CON(n_163),
.SN(n_163)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_95),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_166),
.A2(n_178),
.B(n_121),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_170),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_126),
.A2(n_68),
.B1(n_63),
.B2(n_91),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_169),
.A2(n_126),
.B1(n_140),
.B2(n_145),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_128),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_175),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_122),
.B(n_82),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_122),
.B(n_143),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_82),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_139),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_177),
.A2(n_149),
.B1(n_99),
.B2(n_117),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_136),
.A2(n_3),
.B(n_4),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_SL g226 ( 
.A1(n_181),
.A2(n_188),
.B(n_192),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_176),
.C(n_180),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_172),
.C(n_173),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_146),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_186),
.B(n_190),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_141),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_199),
.B1(n_169),
.B2(n_155),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_148),
.B(n_117),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_198),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_156),
.A2(n_145),
.A3(n_133),
.B1(n_130),
.B2(n_108),
.C1(n_81),
.C2(n_88),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_145),
.B1(n_130),
.B2(n_99),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_207),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_133),
.Y(n_204)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_219),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_166),
.B(n_153),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_210),
.A2(n_229),
.B1(n_6),
.B2(n_7),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_227),
.B1(n_228),
.B2(n_184),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_214),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_218),
.C(n_222),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_162),
.C(n_163),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_159),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_163),
.C(n_152),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_177),
.C(n_160),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_8),
.C(n_10),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_125),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_224),
.B(n_188),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_194),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g237 ( 
.A(n_225),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_158),
.B1(n_125),
.B2(n_127),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_189),
.A2(n_137),
.B1(n_127),
.B2(n_110),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_SL g229 ( 
.A1(n_193),
.A2(n_200),
.B(n_195),
.C(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_110),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_230),
.A2(n_185),
.B(n_190),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_226),
.A2(n_182),
.B1(n_185),
.B2(n_202),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_240),
.B1(n_245),
.B2(n_247),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_243),
.C(n_244),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_212),
.B1(n_224),
.B2(n_222),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_197),
.B1(n_203),
.B2(n_208),
.Y(n_240)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_246),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_188),
.C(n_181),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_184),
.C(n_207),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_214),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_248),
.A2(n_212),
.B1(n_230),
.B2(n_12),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_223),
.C(n_231),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_234),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_251),
.A2(n_253),
.B(n_259),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_248),
.B1(n_216),
.B2(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_239),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_216),
.B(n_217),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_254),
.A2(n_264),
.B(n_265),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_220),
.Y(n_258)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_266),
.C(n_11),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_252),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_231),
.Y(n_264)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_15),
.C(n_17),
.Y(n_266)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_235),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_271),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_233),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_260),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_272)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_276),
.C(n_272),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_12),
.C(n_14),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_258),
.B(n_255),
.CI(n_260),
.CON(n_277),
.SN(n_277)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_277),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_275),
.B(n_253),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_285),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_251),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_262),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_287),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_286),
.A2(n_269),
.B(n_278),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_289),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_271),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_284),
.A2(n_263),
.B1(n_259),
.B2(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_291),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_275),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_257),
.B1(n_263),
.B2(n_268),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_282),
.B1(n_287),
.B2(n_276),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_261),
.C(n_277),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_295),
.A2(n_292),
.B(n_274),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_295),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_301),
.A3(n_292),
.B1(n_296),
.B2(n_267),
.C1(n_270),
.C2(n_254),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_302),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_303),
.C(n_266),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_265),
.Y(n_306)
);


endmodule