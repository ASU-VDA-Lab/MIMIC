module real_jpeg_5879_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_9;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_18),
.C(n_19),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_1),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_1),
.A2(n_45),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_1),
.B(n_31),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_1),
.B(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_3),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_3),
.A2(n_27),
.B1(n_66),
.B2(n_69),
.Y(n_65)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_4),
.Y(n_134)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_5),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_7),
.A2(n_37),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_7),
.A2(n_83),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_109),
.Y(n_8)
);

OAI21xp5_ASAP7_75t_SL g9 ( 
.A1(n_10),
.A2(n_84),
.B(n_108),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_59),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_11),
.B(n_59),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_22),
.B1(n_57),
.B2(n_58),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_17),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_15),
.Y(n_124)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_16),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_16),
.Y(n_135)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_18),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_18),
.A2(n_50),
.B1(n_52),
.B2(n_55),
.Y(n_49)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_22),
.B(n_57),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_31),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_24),
.B(n_48),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_31),
.B(n_122),
.Y(n_121)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_48),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_56),
.A2(n_131),
.B1(n_135),
.B2(n_136),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_73),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_75),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_103),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_100),
.B(n_107),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_94),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_106),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_140),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_113),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_128),
.B1(n_138),
.B2(n_139),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);


endmodule