module fake_aes_5057_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g11 ( .A(n_3), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_3), .B(n_6), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_5), .Y(n_14) );
INVx5_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
NOR2xp33_ASAP7_75t_L g16 ( .A(n_11), .B(n_0), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_15), .B(n_0), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_12), .B(n_1), .Y(n_18) );
OAI21x1_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_13), .B(n_9), .Y(n_19) );
AOI21xp5_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_15), .B(n_14), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_19), .B(n_15), .Y(n_21) );
INVx3_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_22), .B(n_16), .Y(n_24) );
AOI22xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_22), .B1(n_21), .B2(n_15), .Y(n_25) );
O2A1O1Ixp5_ASAP7_75t_L g26 ( .A1(n_23), .A2(n_21), .B(n_22), .C(n_7), .Y(n_26) );
OAI21xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_21), .B(n_22), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_21), .B1(n_4), .B2(n_2), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
NAND4xp75_ASAP7_75t_L g30 ( .A(n_28), .B(n_4), .C(n_21), .D(n_10), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
NAND2xp5_ASAP7_75t_SL g32 ( .A(n_30), .B(n_21), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
AOI22xp33_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_32), .B1(n_30), .B2(n_8), .Y(n_34) );
endmodule