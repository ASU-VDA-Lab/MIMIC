module real_jpeg_12122_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_275, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_275;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_249;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_38),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_0),
.A2(n_38),
.B1(n_56),
.B2(n_57),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_0),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_227)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_5),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_5),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_5),
.A2(n_24),
.B1(n_44),
.B2(n_45),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_5),
.A2(n_24),
.B1(n_56),
.B2(n_57),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_9),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_10),
.A2(n_20),
.B1(n_21),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_10),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_30),
.B(n_41),
.C(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_10),
.A2(n_34),
.B1(n_56),
.B2(n_57),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_10),
.B(n_35),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_10),
.B(n_54),
.C(n_57),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_10),
.B(n_46),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_10),
.B(n_27),
.C(n_31),
.Y(n_173)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_84),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_82),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_69),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_15),
.B(n_69),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_62),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_36),
.C(n_49),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_17),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_17),
.A2(n_71),
.B1(n_123),
.B2(n_125),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_17),
.B(n_123),
.C(n_185),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_17),
.A2(n_71),
.B1(n_93),
.B2(n_94),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_25),
.B1(n_33),
.B2(n_35),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OA21x2_ASAP7_75t_L g76 ( 
.A1(n_19),
.A2(n_29),
.B(n_65),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_21),
.B(n_173),
.Y(n_172)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_25),
.B(n_35),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_29),
.A2(n_64),
.B(n_65),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_31),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_33),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_34),
.A2(n_42),
.B(n_44),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_34),
.B(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_34),
.B(n_60),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_36),
.A2(n_49),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_36),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_46),
.B2(n_47),
.Y(n_36)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_39),
.B(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_39),
.A2(n_46),
.B1(n_81),
.B2(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_41),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_43),
.A2(n_80),
.B(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_43),
.A2(n_68),
.B(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_45),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_45),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_67),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_76),
.C(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_49),
.A2(n_75),
.B1(n_78),
.B2(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_60),
.B(n_61),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_50),
.A2(n_60),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_100),
.Y(n_99)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_51),
.A2(n_55),
.B1(n_98),
.B2(n_100),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_51),
.A2(n_55),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

AO22x1_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_56),
.B(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_97),
.B(n_99),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_60),
.A2(n_99),
.B(n_227),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_61),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.C(n_77),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_70),
.A2(n_76),
.B1(n_175),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_70),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_71),
.B(n_94),
.C(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_76),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_76),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_76),
.A2(n_175),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_76),
.A2(n_175),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_77),
.B(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_78),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_81),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_253),
.B(n_270),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_231),
.B(n_252),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_214),
.B(n_230),
.Y(n_87)
);

OAI321xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_182),
.A3(n_209),
.B1(n_212),
.B2(n_213),
.C(n_275),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_165),
.B(n_181),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_131),
.B(n_164),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_112),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_92),
.B(n_112),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.C(n_101),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_148),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_93),
.A2(n_94),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_94),
.B(n_175),
.C(n_179),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_96),
.B(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_96),
.A2(n_135),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_96),
.A2(n_148),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_100),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_101),
.A2(n_102),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_106),
.A2(n_110),
.B1(n_111),
.B2(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_107),
.B(n_207),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_110),
.A2(n_111),
.B1(n_189),
.B2(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_111),
.A2(n_121),
.B(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_126),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_128),
.C(n_129),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_123),
.B2(n_125),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_116),
.B(n_119),
.C(n_125),
.Y(n_169)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_118),
.B(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_119),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_123),
.A2(n_247),
.B(n_250),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_123),
.B(n_247),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_127),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_130),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_140),
.C(n_142),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_128),
.A2(n_130),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_128),
.B(n_206),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_158),
.B(n_163),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_144),
.B(n_157),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_137),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_142),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_154),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_171),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_149),
.B(n_156),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_188),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_153),
.B(n_155),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_160),
.Y(n_163)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_167),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_170),
.C(n_174),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_196),
.C(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_192),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_192),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_191),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_184),
.B(n_187),
.CI(n_191),
.CON(n_211),
.SN(n_211)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_188),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_208),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_203),
.B2(n_204),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_204),
.C(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_210),
.B(n_211),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g274 ( 
.A(n_211),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_229),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_229),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_218),
.C(n_223),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_224),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_226),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_224),
.A2(n_228),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_228),
.A2(n_237),
.B(n_242),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_233),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_251),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_245),
.B2(n_246),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_245),
.C(n_251),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_250),
.A2(n_257),
.B1(n_258),
.B2(n_262),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_250),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_265),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_264),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_264),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_263),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_262),
.C(n_263),
.Y(n_269)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_265),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_269),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_269),
.Y(n_272)
);


endmodule