module fake_ariane_1131_n_1824 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1824);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1824;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_122),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_36),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_73),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_108),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_63),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_100),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_134),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_60),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_57),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_2),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_81),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_127),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_80),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_15),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_67),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_114),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_135),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_70),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_71),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_110),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_10),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_141),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_3),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_35),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_105),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_27),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_74),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_42),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_62),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_25),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_155),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_96),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_101),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_1),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_24),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_14),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_156),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_40),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_57),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_168),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_167),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_48),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_98),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g218 ( 
.A(n_39),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_28),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_130),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_83),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_86),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_165),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_91),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_24),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_76),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_28),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_51),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_117),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_82),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_103),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_31),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_30),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_148),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_129),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_131),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_162),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_7),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_104),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_26),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_125),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_160),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_159),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_111),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_89),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_85),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_69),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_25),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_92),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_60),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_138),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_90),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_29),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_51),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_48),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_12),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_58),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_16),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_8),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_119),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_11),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_1),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_32),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_27),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_7),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_143),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_120),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_164),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_142),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_12),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_66),
.Y(n_271)
);

BUFx2_ASAP7_75t_SL g272 ( 
.A(n_49),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_112),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_0),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_20),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_64),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_68),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_13),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_30),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_79),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_8),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_62),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_15),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_37),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_26),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_152),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_145),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_95),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_21),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_116),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_33),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_53),
.Y(n_292)
);

CKINVDCx11_ASAP7_75t_R g293 ( 
.A(n_6),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_78),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_65),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_45),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_14),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_34),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_44),
.Y(n_299)
);

BUFx2_ASAP7_75t_SL g300 ( 
.A(n_169),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_55),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_42),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_39),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_50),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_32),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_133),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_16),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_153),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_50),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_20),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_6),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_118),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_99),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_166),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_43),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_55),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_23),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_18),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_59),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_23),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_58),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_61),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_22),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_47),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_43),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_121),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_47),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_136),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_17),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_21),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_102),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_41),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_54),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_77),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_109),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_9),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_158),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_115),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_293),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_218),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_190),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_184),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_305),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_218),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_197),
.B(n_0),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_218),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_192),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_218),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_218),
.B(n_2),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_272),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_237),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_244),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_218),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_294),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_218),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_197),
.B(n_3),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_186),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_218),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_278),
.B(n_4),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_212),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_278),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_326),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_250),
.Y(n_363)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_171),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_254),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_278),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_210),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_253),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_204),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_269),
.B(n_4),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_253),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_208),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_209),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_219),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_212),
.B(n_5),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_225),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_253),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_227),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_232),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_253),
.Y(n_380)
);

XNOR2x1_ASAP7_75t_L g381 ( 
.A(n_171),
.B(n_5),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_259),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_253),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_233),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_258),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_255),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_262),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_289),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_303),
.B(n_210),
.Y(n_389)
);

BUFx6f_ASAP7_75t_SL g390 ( 
.A(n_174),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_258),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_258),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_258),
.Y(n_393)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_191),
.A2(n_231),
.B(n_187),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_256),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_303),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_258),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_292),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_263),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_336),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_336),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_265),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_336),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_301),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_322),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_178),
.Y(n_407)
);

INVxp33_ASAP7_75t_L g408 ( 
.A(n_193),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_325),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_270),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_275),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_183),
.B(n_9),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_214),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_287),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_178),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_279),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_213),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_281),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_179),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_213),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_340),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_361),
.B(n_235),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_394),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_340),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_361),
.B(n_274),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_366),
.B(n_274),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_344),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_348),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_407),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_363),
.A2(n_299),
.B1(n_180),
.B2(n_333),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_366),
.B(n_306),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_348),
.Y(n_437)
);

INVx6_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_353),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_355),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_350),
.B(n_246),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_355),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_342),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_358),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_368),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_368),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_389),
.B(n_200),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_371),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_377),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_377),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_359),
.B(n_203),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_380),
.Y(n_456)
);

CKINVDCx8_ASAP7_75t_R g457 ( 
.A(n_357),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_343),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_383),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_383),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_385),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_385),
.B(n_217),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_391),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_367),
.B(n_302),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_391),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_392),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_392),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_393),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_390),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_408),
.B(n_418),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_369),
.Y(n_471)
);

OA21x2_ASAP7_75t_L g472 ( 
.A1(n_349),
.A2(n_226),
.B(n_220),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_393),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_345),
.B(n_302),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_397),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_397),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_400),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_400),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_401),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_401),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_403),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_403),
.Y(n_482)
);

OR2x6_ASAP7_75t_L g483 ( 
.A(n_356),
.B(n_297),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_406),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_356),
.B(n_418),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_415),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_416),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_416),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_421),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_421),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_412),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_360),
.B(n_396),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_375),
.B(n_297),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_420),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_390),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_370),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_438),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_471),
.B(n_372),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_443),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_425),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_443),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_373),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_443),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_447),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_R g506 ( 
.A(n_445),
.B(n_351),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_450),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_447),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_445),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_447),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_364),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_492),
.B(n_374),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_445),
.Y(n_513)
);

NAND2xp33_ASAP7_75t_L g514 ( 
.A(n_425),
.B(n_376),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_447),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_483),
.A2(n_390),
.B1(n_381),
.B2(n_319),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_450),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_451),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_451),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_483),
.A2(n_494),
.B1(n_438),
.B2(n_497),
.Y(n_520)
);

BUFx4f_ASAP7_75t_L g521 ( 
.A(n_472),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_492),
.B(n_454),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_425),
.B(n_378),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_433),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_433),
.Y(n_525)
);

AO21x2_ASAP7_75t_L g526 ( 
.A1(n_454),
.A2(n_268),
.B(n_239),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g527 ( 
.A(n_422),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_433),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_483),
.A2(n_438),
.B1(n_381),
.B2(n_435),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_483),
.A2(n_240),
.B1(n_309),
.B2(n_315),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_425),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_471),
.B(n_379),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_423),
.B(n_384),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_452),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_423),
.B(n_386),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_433),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_458),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_438),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_433),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_458),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_433),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_471),
.B(n_395),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_496),
.B(n_399),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_456),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_470),
.B(n_402),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_440),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_440),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_456),
.Y(n_549)
);

INVxp33_ASAP7_75t_L g550 ( 
.A(n_435),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_460),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_496),
.B(n_410),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_496),
.B(n_411),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_422),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_460),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_496),
.B(n_417),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_438),
.B(n_419),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_447),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_425),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_422),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_465),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_SL g562 ( 
.A(n_469),
.B(n_339),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_465),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_496),
.B(n_245),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_442),
.B(n_170),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g566 ( 
.A(n_426),
.B(n_199),
.C(n_196),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_465),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_425),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_461),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_465),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_470),
.B(n_319),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_461),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_483),
.A2(n_228),
.B1(n_332),
.B2(n_330),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_463),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_438),
.B(n_413),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_458),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_436),
.B(n_414),
.Y(n_577)
);

OR2x6_ASAP7_75t_L g578 ( 
.A(n_483),
.B(n_300),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_465),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_440),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_434),
.Y(n_581)
);

NOR3xp33_ASAP7_75t_L g582 ( 
.A(n_434),
.B(n_296),
.C(n_216),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_479),
.Y(n_583)
);

OAI21xp33_ASAP7_75t_SL g584 ( 
.A1(n_483),
.A2(n_238),
.B(n_202),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_440),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_422),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_479),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_463),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_487),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_493),
.B(n_179),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_470),
.B(n_248),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_473),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_440),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_473),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_440),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_442),
.B(n_170),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_436),
.B(n_173),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_475),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_494),
.A2(n_307),
.B1(n_299),
.B2(n_317),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_485),
.B(n_257),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_440),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_457),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_475),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_469),
.B(n_173),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_469),
.B(n_175),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_449),
.B(n_341),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_428),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_493),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_493),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_494),
.A2(n_485),
.B1(n_474),
.B2(n_307),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_425),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_479),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_477),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_428),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_477),
.Y(n_615)
);

AO21x2_ASAP7_75t_L g616 ( 
.A1(n_426),
.A2(n_295),
.B(n_290),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_469),
.B(n_175),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_485),
.B(n_261),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_494),
.A2(n_304),
.B1(n_321),
.B2(n_264),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_449),
.B(n_347),
.Y(n_620)
);

AND2x6_ASAP7_75t_L g621 ( 
.A(n_424),
.B(n_191),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_480),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_469),
.B(n_176),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_424),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_424),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_424),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_485),
.B(n_176),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_485),
.B(n_246),
.Y(n_628)
);

INVxp33_ASAP7_75t_SL g629 ( 
.A(n_495),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_424),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_487),
.B(n_177),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_428),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_L g633 ( 
.A(n_432),
.B(n_310),
.C(n_285),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_474),
.B(n_177),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_428),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_428),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_495),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_479),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_480),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_474),
.B(n_352),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_479),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_474),
.B(n_181),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_482),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_474),
.B(n_354),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_424),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_494),
.B(n_181),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_422),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_457),
.B(n_182),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_428),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_507),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_507),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_504),
.Y(n_652)
);

NOR2xp67_ASAP7_75t_L g653 ( 
.A(n_513),
.B(n_491),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_578),
.B(n_600),
.Y(n_654)
);

NAND2x1_ASAP7_75t_L g655 ( 
.A(n_501),
.B(n_424),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_522),
.B(n_431),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_581),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_624),
.B(n_424),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_557),
.B(n_431),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_606),
.A2(n_432),
.B1(n_439),
.B2(n_441),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_517),
.Y(n_661)
);

NOR2x1p5_ASAP7_75t_L g662 ( 
.A(n_590),
.B(n_457),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_624),
.B(n_431),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_554),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_624),
.B(n_431),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_578),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_577),
.B(n_362),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_504),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_511),
.B(n_431),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_624),
.B(n_444),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_520),
.B(n_444),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_504),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_503),
.B(n_444),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_629),
.B(n_365),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_500),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_L g676 ( 
.A(n_501),
.B(n_444),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_512),
.B(n_444),
.Y(n_677)
);

NOR2xp67_ASAP7_75t_L g678 ( 
.A(n_576),
.B(n_491),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_517),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_500),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_620),
.B(n_533),
.Y(n_681)
);

NAND2x1_ASAP7_75t_L g682 ( 
.A(n_501),
.B(n_437),
.Y(n_682)
);

BUFx6f_ASAP7_75t_SL g683 ( 
.A(n_637),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_578),
.B(n_464),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_535),
.B(n_382),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_597),
.B(n_437),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_501),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_498),
.B(n_439),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_581),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_589),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_518),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_498),
.B(n_441),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_538),
.B(n_446),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_608),
.B(n_464),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_578),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_518),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_624),
.B(n_446),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_550),
.A2(n_472),
.B1(n_464),
.B2(n_429),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_578),
.A2(n_472),
.B1(n_464),
.B2(n_313),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_538),
.A2(n_472),
.B1(n_464),
.B2(n_313),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_519),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_519),
.Y(n_702)
);

AO22x2_ASAP7_75t_L g703 ( 
.A1(n_529),
.A2(n_427),
.B1(n_429),
.B2(n_324),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_625),
.B(n_626),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_502),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_565),
.B(n_596),
.Y(n_706)
);

NOR3xp33_ASAP7_75t_L g707 ( 
.A(n_541),
.B(n_316),
.C(n_201),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_628),
.A2(n_320),
.B1(n_201),
.B2(n_311),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_608),
.B(n_472),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_527),
.B(n_427),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_589),
.B(n_427),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_628),
.A2(n_182),
.B1(n_185),
.B2(n_198),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_502),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_509),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_505),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_534),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_534),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_609),
.B(n_387),
.Y(n_718)
);

BUFx5_ASAP7_75t_L g719 ( 
.A(n_621),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_505),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_637),
.B(n_427),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_575),
.B(n_388),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_560),
.B(n_427),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_586),
.B(n_544),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_545),
.Y(n_725)
);

AOI22x1_ASAP7_75t_R g726 ( 
.A1(n_509),
.A2(n_405),
.B1(n_409),
.B2(n_404),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_625),
.B(n_428),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_552),
.B(n_429),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_545),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_553),
.B(n_429),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_625),
.B(n_428),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_625),
.B(n_430),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_546),
.B(n_429),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_628),
.A2(n_318),
.B1(n_311),
.B2(n_317),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_549),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_508),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_625),
.B(n_430),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_508),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_549),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_556),
.B(n_430),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_571),
.B(n_430),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_510),
.Y(n_742)
);

AND2x6_ASAP7_75t_SL g743 ( 
.A(n_640),
.B(n_398),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_551),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_571),
.B(n_430),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_626),
.B(n_430),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_551),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_546),
.B(n_430),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_499),
.B(n_180),
.Y(n_749)
);

AOI221xp5_ASAP7_75t_L g750 ( 
.A1(n_599),
.A2(n_323),
.B1(n_329),
.B2(n_327),
.C(n_320),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_554),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_555),
.Y(n_752)
);

NOR3xp33_ASAP7_75t_L g753 ( 
.A(n_537),
.B(n_323),
.C(n_318),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_510),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_627),
.B(n_430),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_555),
.Y(n_756)
);

O2A1O1Ixp5_ASAP7_75t_L g757 ( 
.A1(n_525),
.A2(n_536),
.B(n_540),
.C(n_528),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_569),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_626),
.B(n_630),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_569),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_515),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_610),
.B(n_490),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_515),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_610),
.B(n_490),
.Y(n_764)
);

NOR2xp67_ASAP7_75t_L g765 ( 
.A(n_602),
.B(n_462),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_558),
.Y(n_766)
);

NOR2x1p5_ASAP7_75t_L g767 ( 
.A(n_590),
.B(n_327),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_558),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_554),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_572),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_572),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_626),
.B(n_490),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_574),
.Y(n_773)
);

AOI221xp5_ASAP7_75t_L g774 ( 
.A1(n_599),
.A2(n_329),
.B1(n_333),
.B2(n_284),
.C(n_291),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_564),
.B(n_490),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_647),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_626),
.B(n_490),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_584),
.A2(n_462),
.B(n_486),
.C(n_489),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_574),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_628),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_588),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_600),
.B(n_490),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_630),
.B(n_490),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_618),
.B(n_490),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_588),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_630),
.B(n_185),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_618),
.B(n_486),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_537),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_L g789 ( 
.A(n_501),
.B(n_172),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_526),
.B(n_486),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_526),
.B(n_486),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_561),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_630),
.B(n_188),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_592),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_561),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_563),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_592),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_526),
.B(n_486),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_630),
.B(n_188),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_L g800 ( 
.A(n_531),
.B(n_172),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_628),
.B(n_482),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_584),
.A2(n_189),
.B1(n_198),
.B2(n_195),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_506),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_573),
.B(n_484),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_645),
.B(n_531),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_532),
.B(n_282),
.Y(n_806)
);

BUFx8_ASAP7_75t_L g807 ( 
.A(n_591),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_594),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_591),
.B(n_484),
.Y(n_809)
);

AND2x2_ASAP7_75t_SL g810 ( 
.A(n_529),
.B(n_516),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_594),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_543),
.B(n_283),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_598),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_647),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_647),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_563),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_567),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_644),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_567),
.B(n_488),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_570),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_657),
.B(n_602),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_659),
.A2(n_645),
.B(n_559),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_689),
.B(n_530),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_662),
.B(n_648),
.Y(n_824)
);

AOI21x1_ASAP7_75t_L g825 ( 
.A1(n_655),
.A2(n_603),
.B(n_598),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_681),
.B(n_530),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_658),
.A2(n_645),
.B(n_559),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_658),
.A2(n_645),
.B(n_559),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_748),
.A2(n_646),
.B(n_634),
.C(n_642),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_740),
.A2(n_645),
.B(n_559),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_780),
.B(n_531),
.Y(n_831)
);

O2A1O1Ixp5_ASAP7_75t_L g832 ( 
.A1(n_786),
.A2(n_603),
.B(n_643),
.C(n_613),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_690),
.B(n_582),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_656),
.A2(n_559),
.B(n_531),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_751),
.Y(n_835)
);

NOR2x1_ASAP7_75t_R g836 ( 
.A(n_654),
.B(n_631),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_818),
.B(n_524),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_687),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_669),
.B(n_619),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_727),
.A2(n_611),
.B(n_531),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_727),
.A2(n_611),
.B(n_568),
.Y(n_841)
);

AND2x2_ASAP7_75t_SL g842 ( 
.A(n_810),
.B(n_521),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_780),
.B(n_611),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_722),
.B(n_667),
.Y(n_844)
);

AOI33xp33_ASAP7_75t_L g845 ( 
.A1(n_750),
.A2(n_622),
.A3(n_643),
.B1(n_613),
.B2(n_639),
.B3(n_615),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_706),
.B(n_524),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_809),
.B(n_611),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_809),
.B(n_615),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_652),
.Y(n_849)
);

AOI21x1_ASAP7_75t_L g850 ( 
.A1(n_805),
.A2(n_639),
.B(n_622),
.Y(n_850)
);

INVx11_ASAP7_75t_L g851 ( 
.A(n_807),
.Y(n_851)
);

BUFx12f_ASAP7_75t_L g852 ( 
.A(n_807),
.Y(n_852)
);

OAI21xp33_ASAP7_75t_L g853 ( 
.A1(n_774),
.A2(n_298),
.B(n_514),
.Y(n_853)
);

AOI21x1_ASAP7_75t_L g854 ( 
.A1(n_805),
.A2(n_759),
.B(n_704),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_652),
.Y(n_855)
);

OAI21xp33_ASAP7_75t_L g856 ( 
.A1(n_749),
.A2(n_523),
.B(n_617),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_714),
.B(n_566),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_721),
.B(n_694),
.Y(n_858)
);

O2A1O1Ixp5_ASAP7_75t_L g859 ( 
.A1(n_786),
.A2(n_521),
.B(n_542),
.C(n_525),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_685),
.B(n_524),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_731),
.A2(n_568),
.B(n_521),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_721),
.B(n_570),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_668),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_732),
.A2(n_568),
.B(n_737),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_788),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_674),
.B(n_566),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_654),
.B(n_524),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_732),
.A2(n_568),
.B(n_528),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_694),
.B(n_765),
.Y(n_869)
);

BUFx4f_ASAP7_75t_L g870 ( 
.A(n_654),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_810),
.A2(n_562),
.B1(n_604),
.B2(n_605),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_737),
.A2(n_568),
.B(n_528),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_733),
.B(n_579),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_802),
.A2(n_579),
.B(n_641),
.C(n_638),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_650),
.A2(n_633),
.B(n_641),
.C(n_638),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_718),
.B(n_633),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_803),
.B(n_711),
.Y(n_877)
);

NAND3xp33_ASAP7_75t_SL g878 ( 
.A(n_806),
.B(n_623),
.C(n_194),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_651),
.A2(n_587),
.B1(n_583),
.B2(n_612),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_686),
.B(n_539),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_807),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_746),
.A2(n_536),
.B(n_525),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_746),
.A2(n_540),
.B(n_536),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_733),
.B(n_583),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_704),
.A2(n_542),
.B(n_540),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_703),
.A2(n_616),
.B1(n_621),
.B2(n_489),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_684),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_751),
.Y(n_888)
);

NOR2xp67_ASAP7_75t_L g889 ( 
.A(n_653),
.B(n_587),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_759),
.A2(n_593),
.B(n_542),
.Y(n_890)
);

OAI21xp33_ASAP7_75t_L g891 ( 
.A1(n_812),
.A2(n_612),
.B(n_539),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_676),
.A2(n_547),
.B(n_593),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_678),
.A2(n_621),
.B1(n_616),
.B2(n_539),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_661),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_679),
.A2(n_585),
.B1(n_580),
.B2(n_539),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_676),
.A2(n_547),
.B(n_593),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_663),
.A2(n_547),
.B(n_595),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_663),
.A2(n_595),
.B(n_649),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_660),
.B(n_616),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_691),
.B(n_621),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_665),
.A2(n_595),
.B(n_649),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_696),
.B(n_621),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_665),
.A2(n_649),
.B(n_607),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_670),
.A2(n_635),
.B(n_614),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_670),
.A2(n_635),
.B(n_614),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_769),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_673),
.A2(n_635),
.B(n_614),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_701),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_702),
.A2(n_585),
.B1(n_548),
.B2(n_580),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_683),
.B(n_548),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_668),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_677),
.A2(n_724),
.B(n_697),
.Y(n_912)
);

OAI321xp33_ASAP7_75t_L g913 ( 
.A1(n_708),
.A2(n_488),
.A3(n_338),
.B1(n_337),
.B2(n_312),
.C(n_459),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_726),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_684),
.B(n_666),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_672),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_683),
.B(n_548),
.Y(n_917)
);

OAI321xp33_ASAP7_75t_L g918 ( 
.A1(n_734),
.A2(n_459),
.A3(n_467),
.B1(n_476),
.B2(n_468),
.C(n_478),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_684),
.Y(n_919)
);

BUFx12f_ASAP7_75t_L g920 ( 
.A(n_743),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_716),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_675),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_717),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_697),
.A2(n_607),
.B(n_548),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_SL g925 ( 
.A(n_683),
.B(n_174),
.Y(n_925)
);

AOI21xp33_ASAP7_75t_L g926 ( 
.A1(n_671),
.A2(n_607),
.B(n_601),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_725),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_729),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_787),
.A2(n_601),
.B(n_585),
.C(n_580),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_735),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_753),
.B(n_174),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_739),
.B(n_621),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_687),
.B(n_719),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_772),
.A2(n_601),
.B(n_585),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_744),
.B(n_621),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_710),
.A2(n_601),
.B(n_580),
.C(n_636),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_703),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_767),
.B(n_288),
.Y(n_938)
);

AOI21x1_ASAP7_75t_L g939 ( 
.A1(n_772),
.A2(n_467),
.B(n_448),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_723),
.A2(n_784),
.B(n_782),
.C(n_760),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_747),
.B(n_636),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_707),
.B(n_288),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_752),
.B(n_636),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_666),
.B(n_632),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_687),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_L g946 ( 
.A(n_728),
.B(n_636),
.C(n_632),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_756),
.B(n_632),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_758),
.B(n_632),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_703),
.Y(n_949)
);

NOR3xp33_ASAP7_75t_L g950 ( 
.A(n_730),
.B(n_331),
.C(n_335),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_770),
.B(n_195),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_801),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_771),
.B(n_308),
.Y(n_953)
);

NOR2x1_ASAP7_75t_L g954 ( 
.A(n_769),
.B(n_224),
.Y(n_954)
);

BUFx12f_ASAP7_75t_L g955 ( 
.A(n_695),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_777),
.A2(n_308),
.B(n_314),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_773),
.B(n_314),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_779),
.B(n_328),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_687),
.Y(n_959)
);

AOI21x1_ASAP7_75t_L g960 ( 
.A1(n_783),
.A2(n_478),
.B(n_476),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_719),
.B(n_664),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_781),
.A2(n_448),
.B(n_478),
.C(n_476),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_783),
.A2(n_328),
.B(n_331),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_695),
.B(n_448),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_755),
.A2(n_334),
.B(n_335),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_776),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_785),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_794),
.A2(n_459),
.B(n_467),
.C(n_468),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_719),
.B(n_334),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_688),
.A2(n_247),
.B(n_221),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_692),
.A2(n_249),
.B(n_222),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_797),
.B(n_468),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_719),
.B(n_466),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_693),
.A2(n_251),
.B(n_205),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_675),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_808),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_811),
.Y(n_977)
);

NOR2x2_ASAP7_75t_L g978 ( 
.A(n_712),
.B(n_715),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_813),
.B(n_288),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_775),
.A2(n_243),
.B(n_223),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_664),
.B(n_10),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_741),
.A2(n_231),
.B(n_224),
.C(n_17),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_715),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_664),
.B(n_11),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_745),
.B(n_206),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_776),
.B(n_13),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_720),
.A2(n_260),
.B(n_230),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_719),
.B(n_466),
.Y(n_988)
);

AO21x1_ASAP7_75t_L g989 ( 
.A1(n_790),
.A2(n_172),
.B(n_455),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_736),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_719),
.B(n_466),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_814),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_699),
.A2(n_266),
.B1(n_211),
.B2(n_229),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_738),
.A2(n_820),
.B(n_763),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_814),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_757),
.A2(n_267),
.B(n_215),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_820),
.A2(n_18),
.B(n_19),
.C(n_22),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_719),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_698),
.B(n_234),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_SL g1000 ( 
.A1(n_709),
.A2(n_207),
.B(n_273),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_815),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_738),
.A2(n_271),
.B(n_242),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_742),
.A2(n_19),
.B(n_29),
.C(n_31),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_804),
.Y(n_1004)
);

AOI21xp33_ASAP7_75t_L g1005 ( 
.A1(n_762),
.A2(n_277),
.B(n_236),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_815),
.B(n_241),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_742),
.A2(n_280),
.B(n_252),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_870),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_844),
.B(n_754),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_842),
.B(n_764),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_852),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_826),
.A2(n_799),
.B1(n_793),
.B2(n_700),
.Y(n_1012)
);

OAI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_848),
.A2(n_791),
.B1(n_798),
.B2(n_816),
.Y(n_1013)
);

NAND2xp33_ASAP7_75t_L g1014 ( 
.A(n_847),
.B(n_754),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_822),
.A2(n_789),
.B(n_800),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_922),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_834),
.A2(n_789),
.B(n_800),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_SL g1018 ( 
.A(n_821),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_830),
.A2(n_793),
.B(n_799),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_860),
.A2(n_778),
.B(n_817),
.C(n_816),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_894),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_827),
.A2(n_682),
.B(n_819),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_828),
.A2(n_817),
.B(n_796),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_865),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_840),
.A2(n_796),
.B(n_795),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_846),
.A2(n_795),
.B(n_792),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_908),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_876),
.B(n_761),
.Y(n_1028)
);

INVxp67_ASAP7_75t_SL g1029 ( 
.A(n_887),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_846),
.A2(n_768),
.B(n_766),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_866),
.B(n_763),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_858),
.A2(n_761),
.B(n_713),
.C(n_705),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1004),
.B(n_713),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_975),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_849),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_841),
.A2(n_705),
.B(n_680),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_823),
.B(n_33),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_952),
.B(n_34),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_865),
.B(n_453),
.Y(n_1039)
);

BUFx2_ASAP7_75t_SL g1040 ( 
.A(n_881),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_870),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_966),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_952),
.B(n_35),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_920),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_912),
.A2(n_286),
.B(n_276),
.Y(n_1045)
);

NOR2x1_ASAP7_75t_SL g1046 ( 
.A(n_838),
.B(n_455),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_855),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_861),
.A2(n_207),
.B(n_466),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_921),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_880),
.A2(n_207),
.B(n_466),
.Y(n_1050)
);

AO32x1_ASAP7_75t_L g1051 ( 
.A1(n_949),
.A2(n_895),
.A3(n_909),
.B1(n_879),
.B2(n_989),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_880),
.A2(n_940),
.B(n_907),
.Y(n_1052)
);

BUFx8_ASAP7_75t_L g1053 ( 
.A(n_833),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_842),
.B(n_481),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_868),
.A2(n_207),
.B(n_466),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_838),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_966),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_872),
.A2(n_207),
.B(n_466),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_857),
.B(n_455),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_864),
.A2(n_481),
.B(n_466),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_860),
.A2(n_871),
.B1(n_837),
.B2(n_928),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_877),
.A2(n_455),
.B1(n_453),
.B2(n_481),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_961),
.A2(n_481),
.B(n_455),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_863),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_838),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_R g1066 ( 
.A(n_925),
.B(n_94),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_836),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_838),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_R g1069 ( 
.A(n_914),
.B(n_878),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_837),
.A2(n_455),
.B1(n_453),
.B2(n_481),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_911),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_873),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_877),
.B(n_38),
.Y(n_1073)
);

NOR2x1_ASAP7_75t_L g1074 ( 
.A(n_835),
.B(n_455),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_923),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_927),
.A2(n_453),
.B1(n_481),
.B2(n_44),
.Y(n_1076)
);

BUFx2_ASAP7_75t_SL g1077 ( 
.A(n_824),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_945),
.B(n_481),
.Y(n_1078)
);

NAND2x1_ASAP7_75t_SL g1079 ( 
.A(n_824),
.B(n_938),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_937),
.A2(n_453),
.B1(n_481),
.B2(n_172),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_930),
.A2(n_453),
.B1(n_41),
.B2(n_45),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_919),
.B(n_40),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_851),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_961),
.A2(n_453),
.B(n_107),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_884),
.A2(n_46),
.B(n_49),
.C(n_52),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_967),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_955),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_916),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_976),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_885),
.A2(n_113),
.B(n_163),
.Y(n_1090)
);

O2A1O1Ixp5_ASAP7_75t_SL g1091 ( 
.A1(n_969),
.A2(n_172),
.B(n_52),
.C(n_53),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_977),
.A2(n_46),
.B1(n_54),
.B2(n_56),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_887),
.B(n_56),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_931),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_890),
.A2(n_126),
.B(n_161),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_875),
.A2(n_59),
.B(n_61),
.C(n_172),
.Y(n_1096)
);

AOI21x1_ASAP7_75t_L g1097 ( 
.A1(n_825),
.A2(n_172),
.B(n_75),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_839),
.B(n_172),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_SL g1099 ( 
.A1(n_874),
.A2(n_72),
.B(n_84),
.C(n_87),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_869),
.B(n_88),
.Y(n_1100)
);

OAI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_845),
.A2(n_950),
.B(n_853),
.Y(n_1101)
);

AO32x1_ASAP7_75t_L g1102 ( 
.A1(n_983),
.A2(n_93),
.A3(n_97),
.B1(n_106),
.B2(n_123),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_945),
.B(n_128),
.Y(n_1103)
);

BUFx12f_ASAP7_75t_L g1104 ( 
.A(n_966),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_942),
.B(n_915),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_915),
.B(n_132),
.Y(n_1106)
);

INVxp67_ASAP7_75t_SL g1107 ( 
.A(n_945),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_856),
.A2(n_139),
.B(n_144),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_829),
.A2(n_899),
.B(n_913),
.C(n_986),
.Y(n_1109)
);

NOR2x1_ASAP7_75t_SL g1110 ( 
.A(n_945),
.B(n_157),
.Y(n_1110)
);

INVx5_ASAP7_75t_L g1111 ( 
.A(n_959),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_986),
.A2(n_146),
.B(n_147),
.C(n_149),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_867),
.B(n_151),
.Y(n_1113)
);

BUFx12f_ASAP7_75t_L g1114 ( 
.A(n_966),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_867),
.B(n_1001),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_1001),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_990),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_979),
.B(n_951),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_959),
.B(n_995),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_953),
.A2(n_958),
.B1(n_957),
.B2(n_862),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_832),
.A2(n_984),
.B(n_981),
.C(n_889),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_959),
.B(n_995),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_950),
.B(n_981),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_978),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_999),
.A2(n_886),
.B1(n_1005),
.B2(n_993),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_972),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_835),
.B(n_888),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_888),
.A2(n_906),
.B1(n_992),
.B2(n_984),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_906),
.A2(n_992),
.B1(n_995),
.B2(n_941),
.Y(n_1129)
);

AND2x6_ASAP7_75t_L g1130 ( 
.A(n_959),
.B(n_995),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_962),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_892),
.A2(n_896),
.B(n_883),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_954),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_944),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_910),
.B(n_917),
.Y(n_1135)
);

OAI22x1_ASAP7_75t_L g1136 ( 
.A1(n_893),
.A2(n_917),
.B1(n_910),
.B2(n_964),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_944),
.B(n_886),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_850),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_964),
.B(n_1006),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_998),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_943),
.A2(n_947),
.B1(n_948),
.B2(n_935),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_946),
.A2(n_985),
.B1(n_926),
.B2(n_891),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_882),
.A2(n_905),
.B(n_904),
.Y(n_1143)
);

AO21x2_ASAP7_75t_L g1144 ( 
.A1(n_996),
.A2(n_946),
.B(n_900),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_854),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_831),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_968),
.Y(n_1147)
);

O2A1O1Ixp5_ASAP7_75t_L g1148 ( 
.A1(n_859),
.A2(n_969),
.B(n_832),
.C(n_932),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_903),
.A2(n_901),
.B(n_898),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_875),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_902),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_939),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_994),
.B(n_831),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_998),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_997),
.A2(n_1003),
.B(n_982),
.C(n_936),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_843),
.B(n_963),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_843),
.B(n_956),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_897),
.A2(n_924),
.B(n_934),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_933),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_960),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_859),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_965),
.B(n_970),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1052),
.A2(n_991),
.B(n_988),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1031),
.B(n_929),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_SL g1165 ( 
.A1(n_1123),
.A2(n_991),
.B(n_973),
.C(n_988),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1021),
.Y(n_1166)
);

BUFx12f_ASAP7_75t_L g1167 ( 
.A(n_1083),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1061),
.A2(n_971),
.B(n_974),
.C(n_1002),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1037),
.A2(n_973),
.B1(n_987),
.B2(n_1007),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1132),
.A2(n_1000),
.B(n_980),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1121),
.A2(n_918),
.B(n_1143),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1149),
.A2(n_1158),
.B(n_1020),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1141),
.A2(n_1015),
.B(n_1017),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1025),
.A2(n_1023),
.B(n_1036),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_SL g1175 ( 
.A(n_1037),
.B(n_1066),
.C(n_1069),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1073),
.A2(n_1120),
.B(n_1096),
.C(n_1101),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1048),
.A2(n_1097),
.B(n_1019),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_1024),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1018),
.B(n_1053),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1124),
.B(n_1105),
.Y(n_1180)
);

INVx4_ASAP7_75t_SL g1181 ( 
.A(n_1130),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1162),
.A2(n_1022),
.B(n_1050),
.Y(n_1182)
);

OA21x2_ASAP7_75t_L g1183 ( 
.A1(n_1148),
.A2(n_1161),
.B(n_1142),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1096),
.A2(n_1118),
.B(n_1109),
.C(n_1116),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_SL g1185 ( 
.A1(n_1066),
.A2(n_1137),
.B1(n_1094),
.B2(n_1053),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1012),
.A2(n_1148),
.B(n_1026),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1116),
.A2(n_1085),
.B(n_1072),
.C(n_1092),
.Y(n_1187)
);

OR2x6_ASAP7_75t_L g1188 ( 
.A(n_1077),
.B(n_1008),
.Y(n_1188)
);

CKINVDCx11_ASAP7_75t_R g1189 ( 
.A(n_1044),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1030),
.A2(n_1013),
.B(n_1108),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1028),
.B(n_1126),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1009),
.B(n_1079),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1160),
.A2(n_1153),
.B(n_1058),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1013),
.A2(n_1128),
.B(n_1113),
.Y(n_1194)
);

AOI221xp5_ASAP7_75t_L g1195 ( 
.A1(n_1072),
.A2(n_1085),
.B1(n_1125),
.B2(n_1081),
.C(n_1089),
.Y(n_1195)
);

BUFx2_ASAP7_75t_R g1196 ( 
.A(n_1011),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1027),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1160),
.A2(n_1055),
.B(n_1152),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1029),
.B(n_1135),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1049),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1138),
.A2(n_1136),
.A3(n_1098),
.B(n_1150),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1075),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_1156),
.A2(n_1157),
.A3(n_1100),
.B(n_1117),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1029),
.B(n_1115),
.Y(n_1204)
);

INVxp67_ASAP7_75t_SL g1205 ( 
.A(n_1033),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1067),
.B(n_1039),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1113),
.A2(n_1142),
.B(n_1014),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1093),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1140),
.A2(n_1078),
.B(n_1100),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1086),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1041),
.A2(n_1134),
.B1(n_1040),
.B2(n_1125),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1134),
.B(n_1010),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1104),
.Y(n_1213)
);

AOI221xp5_ASAP7_75t_L g1214 ( 
.A1(n_1155),
.A2(n_1043),
.B1(n_1038),
.B2(n_1069),
.C(n_1076),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1131),
.A2(n_1147),
.B1(n_1062),
.B2(n_1082),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1016),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1010),
.B(n_1127),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1140),
.A2(n_1078),
.B(n_1099),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_1114),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1041),
.B(n_1008),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1060),
.A2(n_1090),
.B(n_1095),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1155),
.A2(n_1032),
.B(n_1139),
.C(n_1045),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1034),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1087),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1035),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1059),
.A2(n_1112),
.B1(n_1054),
.B2(n_1080),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1032),
.A2(n_1084),
.B(n_1063),
.Y(n_1227)
);

AO22x2_ASAP7_75t_L g1228 ( 
.A1(n_1054),
.A2(n_1064),
.B1(n_1047),
.B2(n_1071),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1088),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1111),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1099),
.A2(n_1129),
.B(n_1146),
.C(n_1103),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1146),
.A2(n_1103),
.B(n_1070),
.C(n_1133),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1151),
.A2(n_1080),
.B1(n_1106),
.B2(n_1159),
.Y(n_1233)
);

OAI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1159),
.A2(n_1042),
.B1(n_1057),
.B2(n_1111),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1051),
.A2(n_1110),
.A3(n_1046),
.B(n_1144),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1042),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1130),
.B(n_1107),
.Y(n_1237)
);

INVx3_ASAP7_75t_SL g1238 ( 
.A(n_1111),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1159),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1119),
.B(n_1122),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1130),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1091),
.A2(n_1074),
.B(n_1122),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1051),
.A2(n_1144),
.A3(n_1145),
.B(n_1102),
.Y(n_1243)
);

INVx4_ASAP7_75t_L g1244 ( 
.A(n_1130),
.Y(n_1244)
);

OAI22x1_ASAP7_75t_L g1245 ( 
.A1(n_1119),
.A2(n_1102),
.B1(n_1051),
.B2(n_1159),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1102),
.A2(n_1154),
.B(n_1145),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1145),
.A2(n_1056),
.B(n_1065),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1145),
.A2(n_1056),
.B(n_1065),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1065),
.A2(n_1132),
.B(n_1143),
.Y(n_1249)
);

AO21x2_ASAP7_75t_L g1250 ( 
.A1(n_1068),
.A2(n_1013),
.B(n_989),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1068),
.A2(n_531),
.B(n_501),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1068),
.A2(n_1132),
.B(n_1143),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1052),
.A2(n_531),
.B(n_501),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1052),
.A2(n_531),
.B(n_501),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_1083),
.Y(n_1255)
);

OR2x6_ASAP7_75t_L g1256 ( 
.A(n_1077),
.B(n_1008),
.Y(n_1256)
);

AOI221x1_ASAP7_75t_L g1257 ( 
.A1(n_1101),
.A2(n_1109),
.B1(n_1061),
.B2(n_1123),
.C(n_826),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1021),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1132),
.A2(n_1143),
.B(n_1149),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1052),
.A2(n_531),
.B(n_501),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1021),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1037),
.A2(n_826),
.B1(n_848),
.B2(n_1061),
.Y(n_1262)
);

AOI221x1_ASAP7_75t_L g1263 ( 
.A1(n_1101),
.A2(n_1109),
.B1(n_1061),
.B2(n_1123),
.C(n_826),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1021),
.Y(n_1264)
);

AO21x2_ASAP7_75t_L g1265 ( 
.A1(n_1013),
.A2(n_989),
.B(n_1138),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1052),
.A2(n_531),
.B(n_501),
.Y(n_1266)
);

AO21x1_ASAP7_75t_L g1267 ( 
.A1(n_1123),
.A2(n_1061),
.B(n_1096),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1021),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1031),
.B(n_1028),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_1053),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1052),
.A2(n_531),
.B(n_501),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1031),
.B(n_1028),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1132),
.A2(n_1143),
.B(n_1149),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1052),
.A2(n_531),
.B(n_501),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1061),
.A2(n_1020),
.B(n_1012),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1083),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_SL g1277 ( 
.A1(n_1123),
.A2(n_1121),
.B(n_1061),
.C(n_847),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1037),
.B(n_844),
.Y(n_1278)
);

NOR2xp67_ASAP7_75t_L g1279 ( 
.A(n_1083),
.B(n_852),
.Y(n_1279)
);

AOI221xp5_ASAP7_75t_SL g1280 ( 
.A1(n_1072),
.A2(n_1085),
.B1(n_1101),
.B2(n_1061),
.C(n_1096),
.Y(n_1280)
);

INVx8_ASAP7_75t_L g1281 ( 
.A(n_1104),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1037),
.A2(n_844),
.B1(n_674),
.B2(n_667),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1008),
.Y(n_1283)
);

AOI221xp5_ASAP7_75t_SL g1284 ( 
.A1(n_1072),
.A2(n_1085),
.B1(n_1101),
.B2(n_1061),
.C(n_1096),
.Y(n_1284)
);

INVx2_ASAP7_75t_SL g1285 ( 
.A(n_1083),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1024),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1052),
.A2(n_531),
.B(n_501),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1061),
.A2(n_1020),
.B(n_1012),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1024),
.Y(n_1289)
);

AOI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1052),
.A2(n_1132),
.B(n_1143),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1132),
.A2(n_1143),
.B(n_1149),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1037),
.A2(n_844),
.B1(n_674),
.B2(n_667),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1037),
.B(n_844),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1117),
.Y(n_1294)
);

O2A1O1Ixp5_ASAP7_75t_L g1295 ( 
.A1(n_1052),
.A2(n_844),
.B(n_1123),
.C(n_681),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1031),
.B(n_1028),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1123),
.A2(n_681),
.B(n_826),
.C(n_844),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1037),
.B(n_844),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1031),
.B(n_1028),
.Y(n_1299)
);

AOI221x1_ASAP7_75t_L g1300 ( 
.A1(n_1101),
.A2(n_1109),
.B1(n_1061),
.B2(n_1123),
.C(n_826),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1008),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1135),
.B(n_844),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1132),
.A2(n_1143),
.B(n_1149),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1052),
.A2(n_531),
.B(n_501),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1052),
.A2(n_531),
.B(n_501),
.Y(n_1305)
);

O2A1O1Ixp5_ASAP7_75t_L g1306 ( 
.A1(n_1052),
.A2(n_844),
.B(n_1123),
.C(n_681),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1037),
.A2(n_844),
.B1(n_674),
.B2(n_667),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1052),
.A2(n_531),
.B(n_501),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1278),
.B(n_1293),
.Y(n_1309)
);

CKINVDCx6p67_ASAP7_75t_R g1310 ( 
.A(n_1189),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1244),
.B(n_1241),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1166),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1206),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1197),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1282),
.A2(n_1307),
.B1(n_1292),
.B2(n_1262),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1262),
.A2(n_1175),
.B1(n_1267),
.B2(n_1298),
.Y(n_1316)
);

INVx6_ASAP7_75t_L g1317 ( 
.A(n_1281),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1200),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1202),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1257),
.A2(n_1300),
.B1(n_1263),
.B2(n_1275),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1195),
.A2(n_1275),
.B1(n_1288),
.B2(n_1214),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1210),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1288),
.A2(n_1302),
.B1(n_1185),
.B2(n_1207),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1258),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1238),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1208),
.A2(n_1194),
.B1(n_1215),
.B2(n_1272),
.Y(n_1326)
);

INVxp67_ASAP7_75t_SL g1327 ( 
.A(n_1183),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1261),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1215),
.A2(n_1226),
.B1(n_1284),
.B2(n_1280),
.Y(n_1329)
);

INVx3_ASAP7_75t_SL g1330 ( 
.A(n_1281),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1230),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1269),
.A2(n_1272),
.B1(n_1296),
.B2(n_1299),
.Y(n_1332)
);

INVx6_ASAP7_75t_L g1333 ( 
.A(n_1181),
.Y(n_1333)
);

BUFx2_ASAP7_75t_SL g1334 ( 
.A(n_1279),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1264),
.Y(n_1335)
);

INVx6_ASAP7_75t_L g1336 ( 
.A(n_1181),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1268),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1167),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_1255),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1196),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1181),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1289),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1226),
.A2(n_1284),
.B1(n_1280),
.B2(n_1205),
.Y(n_1343)
);

BUFx4_ASAP7_75t_R g1344 ( 
.A(n_1224),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1199),
.B(n_1204),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1176),
.A2(n_1199),
.B1(n_1184),
.B2(n_1187),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_SL g1347 ( 
.A1(n_1270),
.A2(n_1211),
.B(n_1179),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1192),
.A2(n_1216),
.B1(n_1294),
.B2(n_1299),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1213),
.Y(n_1349)
);

CKINVDCx11_ASAP7_75t_R g1350 ( 
.A(n_1178),
.Y(n_1350)
);

BUFx12f_ASAP7_75t_L g1351 ( 
.A(n_1285),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1269),
.A2(n_1296),
.B1(n_1229),
.B2(n_1223),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1225),
.A2(n_1180),
.B1(n_1191),
.B2(n_1233),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1178),
.A2(n_1204),
.B1(n_1217),
.B2(n_1222),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1217),
.A2(n_1169),
.B1(n_1286),
.B2(n_1164),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1188),
.A2(n_1256),
.B1(n_1219),
.B2(n_1220),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1228),
.A2(n_1212),
.B1(n_1164),
.B2(n_1256),
.Y(n_1357)
);

BUFx8_ASAP7_75t_L g1358 ( 
.A(n_1196),
.Y(n_1358)
);

BUFx8_ASAP7_75t_L g1359 ( 
.A(n_1301),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1219),
.B(n_1283),
.Y(n_1360)
);

INVx8_ASAP7_75t_L g1361 ( 
.A(n_1188),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1212),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1228),
.A2(n_1239),
.B1(n_1245),
.B2(n_1186),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1186),
.A2(n_1183),
.B1(n_1171),
.B2(n_1265),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1265),
.A2(n_1190),
.B1(n_1250),
.B2(n_1283),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1237),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1242),
.A2(n_1236),
.B1(n_1240),
.B2(n_1250),
.Y(n_1367)
);

CKINVDCx6p67_ASAP7_75t_R g1368 ( 
.A(n_1237),
.Y(n_1368)
);

CKINVDCx11_ASAP7_75t_R g1369 ( 
.A(n_1277),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1209),
.A2(n_1173),
.B1(n_1168),
.B2(n_1231),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1248),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1234),
.Y(n_1372)
);

INVx6_ASAP7_75t_L g1373 ( 
.A(n_1248),
.Y(n_1373)
);

CKINVDCx11_ASAP7_75t_R g1374 ( 
.A(n_1295),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1247),
.Y(n_1375)
);

BUFx4f_ASAP7_75t_SL g1376 ( 
.A(n_1232),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1242),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1246),
.A2(n_1218),
.B1(n_1163),
.B2(n_1198),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1306),
.A2(n_1172),
.B1(n_1227),
.B2(n_1203),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_SL g1380 ( 
.A1(n_1221),
.A2(n_1170),
.B1(n_1243),
.B2(n_1182),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1249),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1251),
.A2(n_1260),
.B(n_1305),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1243),
.A2(n_1235),
.B1(n_1249),
.B2(n_1201),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1243),
.A2(n_1235),
.B1(n_1201),
.B2(n_1177),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1253),
.A2(n_1271),
.B1(n_1304),
.B2(n_1287),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1254),
.Y(n_1386)
);

BUFx12f_ASAP7_75t_L g1387 ( 
.A(n_1165),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1235),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1266),
.A2(n_1308),
.B1(n_1274),
.B2(n_1290),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1193),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1252),
.B(n_1259),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1273),
.A2(n_1291),
.B1(n_1303),
.B2(n_1174),
.Y(n_1392)
);

OAI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1282),
.A2(n_1292),
.B1(n_1307),
.B2(n_826),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1282),
.A2(n_1307),
.B1(n_1292),
.B2(n_844),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1289),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1206),
.Y(n_1396)
);

CKINVDCx11_ASAP7_75t_R g1397 ( 
.A(n_1189),
.Y(n_1397)
);

INVx6_ASAP7_75t_L g1398 ( 
.A(n_1281),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1282),
.A2(n_1307),
.B1(n_1292),
.B2(n_844),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1278),
.B(n_1293),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1282),
.A2(n_810),
.B1(n_667),
.B2(n_844),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1282),
.A2(n_810),
.B1(n_1307),
.B2(n_1292),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1166),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1282),
.A2(n_810),
.B1(n_1307),
.B2(n_1292),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1282),
.A2(n_810),
.B1(n_1307),
.B2(n_1292),
.Y(n_1405)
);

INVx6_ASAP7_75t_L g1406 ( 
.A(n_1281),
.Y(n_1406)
);

INVxp67_ASAP7_75t_SL g1407 ( 
.A(n_1183),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1282),
.A2(n_1292),
.B1(n_1307),
.B2(n_1297),
.Y(n_1408)
);

CKINVDCx11_ASAP7_75t_R g1409 ( 
.A(n_1189),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1262),
.A2(n_810),
.B1(n_1037),
.B2(n_1124),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1276),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_SL g1412 ( 
.A1(n_1262),
.A2(n_810),
.B1(n_1037),
.B2(n_1124),
.Y(n_1412)
);

BUFx8_ASAP7_75t_SL g1413 ( 
.A(n_1167),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1282),
.A2(n_810),
.B1(n_667),
.B2(n_844),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1282),
.A2(n_810),
.B1(n_667),
.B2(n_844),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1289),
.Y(n_1416)
);

OAI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1282),
.A2(n_1292),
.B1(n_1307),
.B2(n_826),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1282),
.A2(n_810),
.B1(n_1307),
.B2(n_1292),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1282),
.A2(n_1292),
.B1(n_1307),
.B2(n_1297),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1289),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1278),
.B(n_1293),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1282),
.A2(n_810),
.B1(n_667),
.B2(n_844),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1362),
.B(n_1400),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1375),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_1421),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1375),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1382),
.A2(n_1389),
.B(n_1385),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1391),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1313),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1312),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1314),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1318),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1319),
.B(n_1322),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1345),
.B(n_1366),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1396),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1324),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1328),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1335),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1364),
.A2(n_1365),
.B(n_1327),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1337),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1355),
.B(n_1354),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1387),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1370),
.A2(n_1365),
.B(n_1378),
.Y(n_1443)
);

AO31x2_ASAP7_75t_L g1444 ( 
.A1(n_1346),
.A2(n_1377),
.A3(n_1390),
.B(n_1419),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1373),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1332),
.B(n_1326),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1381),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1364),
.A2(n_1363),
.B(n_1367),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1403),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1327),
.A2(n_1407),
.B(n_1311),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1407),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1329),
.B(n_1343),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1368),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1386),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1373),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1329),
.B(n_1343),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1309),
.B(n_1326),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1371),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1383),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1321),
.B(n_1384),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1383),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1321),
.A2(n_1408),
.B(n_1393),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1388),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1384),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1379),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1374),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1379),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1320),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1357),
.B(n_1316),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1372),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1320),
.A2(n_1393),
.B(n_1417),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1360),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1352),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1410),
.B(n_1412),
.Y(n_1474)
);

AO21x2_ASAP7_75t_L g1475 ( 
.A1(n_1417),
.A2(n_1394),
.B(n_1399),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1401),
.A2(n_1422),
.B1(n_1414),
.B2(n_1415),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1315),
.B(n_1323),
.Y(n_1477)
);

OR2x6_ASAP7_75t_L g1478 ( 
.A(n_1333),
.B(n_1341),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1392),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1372),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1372),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1392),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1380),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1413),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1323),
.B(n_1418),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1376),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1331),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1331),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1348),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1402),
.B(n_1418),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1402),
.B(n_1405),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1325),
.Y(n_1492)
);

INVx4_ASAP7_75t_L g1493 ( 
.A(n_1336),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1404),
.B(n_1405),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1325),
.B(n_1404),
.Y(n_1495)
);

NAND4xp25_ASAP7_75t_L g1496 ( 
.A(n_1347),
.B(n_1420),
.C(n_1416),
.D(n_1342),
.Y(n_1496)
);

INVx4_ASAP7_75t_L g1497 ( 
.A(n_1341),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1353),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1359),
.Y(n_1499)
);

AO21x1_ASAP7_75t_L g1500 ( 
.A1(n_1441),
.A2(n_1356),
.B(n_1344),
.Y(n_1500)
);

O2A1O1Ixp5_ASAP7_75t_L g1501 ( 
.A1(n_1462),
.A2(n_1369),
.B(n_1350),
.C(n_1358),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1474),
.A2(n_1361),
.B(n_1340),
.C(n_1334),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1457),
.B(n_1349),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1434),
.B(n_1395),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1430),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1457),
.B(n_1339),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1484),
.Y(n_1507)
);

AOI211xp5_ASAP7_75t_L g1508 ( 
.A1(n_1471),
.A2(n_1330),
.B(n_1411),
.C(n_1338),
.Y(n_1508)
);

AOI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1474),
.A2(n_1351),
.B1(n_1358),
.B2(n_1317),
.Y(n_1509)
);

NAND2xp33_ASAP7_75t_L g1510 ( 
.A(n_1442),
.B(n_1330),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1486),
.B(n_1406),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1434),
.B(n_1310),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1483),
.B(n_1423),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1430),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1429),
.B(n_1409),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1486),
.B(n_1454),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1428),
.B(n_1398),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1454),
.Y(n_1518)
);

NOR2x1_ASAP7_75t_SL g1519 ( 
.A(n_1478),
.B(n_1397),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1455),
.B(n_1428),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1453),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1477),
.A2(n_1476),
.B1(n_1452),
.B2(n_1456),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1428),
.B(n_1479),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1472),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1447),
.B(n_1435),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1475),
.A2(n_1494),
.B(n_1446),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1499),
.Y(n_1527)
);

AO32x2_ASAP7_75t_L g1528 ( 
.A1(n_1445),
.A2(n_1492),
.A3(n_1460),
.B1(n_1493),
.B2(n_1497),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1458),
.B(n_1433),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1496),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1486),
.B(n_1475),
.Y(n_1531)
);

A2O1A1Ixp33_ASAP7_75t_SL g1532 ( 
.A1(n_1482),
.A2(n_1424),
.B(n_1426),
.C(n_1468),
.Y(n_1532)
);

AOI221x1_ASAP7_75t_SL g1533 ( 
.A1(n_1431),
.A2(n_1449),
.B1(n_1440),
.B2(n_1438),
.C(n_1437),
.Y(n_1533)
);

AO32x2_ASAP7_75t_L g1534 ( 
.A1(n_1492),
.A2(n_1460),
.A3(n_1497),
.B1(n_1493),
.B2(n_1499),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1433),
.B(n_1465),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1465),
.B(n_1467),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1456),
.A2(n_1485),
.B(n_1495),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1485),
.A2(n_1443),
.B(n_1490),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1444),
.Y(n_1539)
);

OA21x2_ASAP7_75t_L g1540 ( 
.A1(n_1427),
.A2(n_1443),
.B(n_1448),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1448),
.A2(n_1467),
.B(n_1450),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1432),
.Y(n_1542)
);

A2O1A1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1490),
.A2(n_1491),
.B(n_1469),
.C(n_1464),
.Y(n_1543)
);

AO32x2_ASAP7_75t_L g1544 ( 
.A1(n_1493),
.A2(n_1497),
.A3(n_1461),
.B1(n_1459),
.B2(n_1444),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1425),
.B(n_1463),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1436),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1498),
.A2(n_1469),
.B1(n_1491),
.B2(n_1489),
.Y(n_1547)
);

NAND3xp33_ASAP7_75t_SL g1548 ( 
.A(n_1466),
.B(n_1453),
.C(n_1464),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1436),
.B(n_1437),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1505),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1523),
.B(n_1439),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1531),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1529),
.B(n_1444),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1514),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1542),
.Y(n_1555)
);

NAND3xp33_ASAP7_75t_L g1556 ( 
.A(n_1526),
.B(n_1487),
.C(n_1488),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1523),
.B(n_1439),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1546),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1520),
.B(n_1439),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1522),
.A2(n_1498),
.B1(n_1489),
.B2(n_1459),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1540),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1531),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1533),
.B(n_1444),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1538),
.A2(n_1461),
.B1(n_1473),
.B2(n_1439),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1508),
.B(n_1442),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1549),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1527),
.B(n_1442),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1549),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1520),
.B(n_1540),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1543),
.A2(n_1470),
.B1(n_1480),
.B2(n_1481),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1534),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1540),
.B(n_1444),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1541),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1535),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1535),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1513),
.B(n_1528),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1524),
.B(n_1444),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1528),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1513),
.B(n_1451),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1541),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1528),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1518),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1544),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1544),
.B(n_1451),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1576),
.B(n_1525),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1550),
.Y(n_1586)
);

BUFx2_ASAP7_75t_SL g1587 ( 
.A(n_1565),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1577),
.B(n_1506),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1554),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1576),
.B(n_1571),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1567),
.B(n_1530),
.Y(n_1591)
);

AO21x2_ASAP7_75t_L g1592 ( 
.A1(n_1573),
.A2(n_1532),
.B(n_1539),
.Y(n_1592)
);

AOI221xp5_ASAP7_75t_L g1593 ( 
.A1(n_1563),
.A2(n_1543),
.B1(n_1537),
.B2(n_1548),
.C(n_1536),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1554),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1577),
.B(n_1553),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1553),
.B(n_1503),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1576),
.B(n_1518),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1571),
.Y(n_1598)
);

NOR3xp33_ASAP7_75t_L g1599 ( 
.A(n_1563),
.B(n_1501),
.C(n_1521),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1584),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1559),
.B(n_1519),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1574),
.B(n_1545),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1579),
.B(n_1504),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1555),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1574),
.B(n_1517),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1555),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1564),
.A2(n_1500),
.B1(n_1536),
.B2(n_1547),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1575),
.B(n_1517),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1558),
.Y(n_1609)
);

INVx4_ASAP7_75t_L g1610 ( 
.A(n_1582),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1558),
.Y(n_1611)
);

NOR3xp33_ASAP7_75t_SL g1612 ( 
.A(n_1556),
.B(n_1527),
.C(n_1516),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1551),
.B(n_1532),
.Y(n_1613)
);

OAI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1564),
.A2(n_1570),
.B1(n_1560),
.B2(n_1556),
.C(n_1502),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1566),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1561),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1590),
.B(n_1569),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1592),
.Y(n_1618)
);

NAND2xp33_ASAP7_75t_L g1619 ( 
.A(n_1612),
.B(n_1442),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1598),
.B(n_1578),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1590),
.B(n_1569),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1598),
.B(n_1578),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1586),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1600),
.B(n_1569),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1588),
.B(n_1581),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1597),
.B(n_1551),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1586),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1613),
.B(n_1583),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1589),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1613),
.B(n_1557),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1601),
.B(n_1559),
.Y(n_1631)
);

NOR2x1_ASAP7_75t_SL g1632 ( 
.A(n_1587),
.B(n_1582),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1585),
.B(n_1559),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1585),
.B(n_1599),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1601),
.B(n_1587),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1594),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1594),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1601),
.B(n_1605),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1604),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1606),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1605),
.B(n_1568),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1595),
.B(n_1583),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1606),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1608),
.B(n_1584),
.Y(n_1644)
);

INVx3_ASAP7_75t_L g1645 ( 
.A(n_1616),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1592),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1637),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1618),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1630),
.B(n_1593),
.Y(n_1649)
);

NAND3xp33_ASAP7_75t_L g1650 ( 
.A(n_1628),
.B(n_1614),
.C(n_1561),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1637),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1623),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1632),
.B(n_1610),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1632),
.B(n_1610),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1618),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1638),
.B(n_1610),
.Y(n_1656)
);

NAND2x1p5_ASAP7_75t_L g1657 ( 
.A(n_1635),
.B(n_1610),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1630),
.B(n_1609),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1638),
.B(n_1608),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1623),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1638),
.B(n_1602),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1627),
.Y(n_1662)
);

NAND3x1_ASAP7_75t_L g1663 ( 
.A(n_1634),
.B(n_1509),
.C(n_1591),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1627),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1630),
.B(n_1609),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1618),
.Y(n_1666)
);

OAI33xp33_ASAP7_75t_L g1667 ( 
.A1(n_1628),
.A2(n_1595),
.A3(n_1552),
.B1(n_1562),
.B2(n_1611),
.B3(n_1596),
.Y(n_1667)
);

INVxp67_ASAP7_75t_SL g1668 ( 
.A(n_1628),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1629),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1642),
.B(n_1603),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1641),
.B(n_1634),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1634),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1635),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1641),
.B(n_1625),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1629),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1619),
.A2(n_1614),
.B1(n_1607),
.B2(n_1572),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1636),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1636),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1635),
.B(n_1602),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1618),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1641),
.B(n_1611),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1642),
.B(n_1603),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1617),
.B(n_1615),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1625),
.B(n_1596),
.Y(n_1684)
);

NOR2x1_ASAP7_75t_L g1685 ( 
.A(n_1619),
.B(n_1515),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1639),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1639),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1652),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1668),
.B(n_1640),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1661),
.B(n_1659),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1671),
.B(n_1620),
.Y(n_1691)
);

NOR3xp33_ASAP7_75t_L g1692 ( 
.A(n_1650),
.B(n_1646),
.C(n_1645),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1649),
.B(n_1640),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1652),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1648),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1661),
.B(n_1617),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1670),
.B(n_1620),
.Y(n_1697)
);

NOR2x1_ASAP7_75t_L g1698 ( 
.A(n_1685),
.B(n_1647),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1676),
.A2(n_1583),
.B1(n_1572),
.B2(n_1646),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_1673),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1672),
.B(n_1647),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1659),
.B(n_1617),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1660),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1679),
.B(n_1621),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1651),
.B(n_1643),
.Y(n_1705)
);

INVxp67_ASAP7_75t_SL g1706 ( 
.A(n_1663),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1670),
.B(n_1620),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1679),
.B(n_1621),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1653),
.B(n_1631),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1653),
.B(n_1654),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1651),
.B(n_1643),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1660),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1656),
.B(n_1621),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1669),
.B(n_1644),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1656),
.B(n_1626),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1658),
.B(n_1665),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1662),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1682),
.B(n_1644),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1662),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1657),
.B(n_1626),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1664),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1682),
.B(n_1644),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1657),
.B(n_1626),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_1701),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1693),
.B(n_1674),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1700),
.Y(n_1726)
);

OAI22xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1706),
.A2(n_1663),
.B1(n_1642),
.B2(n_1622),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1700),
.B(n_1683),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1699),
.A2(n_1667),
.B1(n_1572),
.B2(n_1646),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1693),
.B(n_1507),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1717),
.Y(n_1731)
);

AOI222xp33_ASAP7_75t_L g1732 ( 
.A1(n_1698),
.A2(n_1646),
.B1(n_1655),
.B2(n_1648),
.C1(n_1666),
.C2(n_1680),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1718),
.B(n_1684),
.Y(n_1733)
);

OAI31xp33_ASAP7_75t_L g1734 ( 
.A1(n_1692),
.A2(n_1622),
.A3(n_1657),
.B(n_1502),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1690),
.B(n_1683),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1688),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1690),
.B(n_1681),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1698),
.A2(n_1718),
.B1(n_1722),
.B2(n_1709),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1710),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1722),
.A2(n_1631),
.B1(n_1624),
.B2(n_1654),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1697),
.B(n_1622),
.Y(n_1741)
);

OAI32xp33_ASAP7_75t_L g1742 ( 
.A1(n_1691),
.A2(n_1645),
.A3(n_1624),
.B1(n_1686),
.B2(n_1675),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1688),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1701),
.B(n_1633),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1694),
.Y(n_1745)
);

NOR4xp25_ASAP7_75t_SL g1746 ( 
.A(n_1694),
.B(n_1687),
.C(n_1664),
.D(n_1686),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1703),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1695),
.A2(n_1584),
.B1(n_1592),
.B2(n_1580),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1703),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1745),
.Y(n_1750)
);

NAND2xp33_ASAP7_75t_SL g1751 ( 
.A(n_1746),
.B(n_1697),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1745),
.Y(n_1752)
);

NAND2xp33_ASAP7_75t_SL g1753 ( 
.A(n_1728),
.B(n_1707),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1726),
.B(n_1507),
.Y(n_1754)
);

A2O1A1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1729),
.A2(n_1707),
.B(n_1691),
.C(n_1689),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1730),
.B(n_1710),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1739),
.Y(n_1757)
);

NAND3xp33_ASAP7_75t_L g1758 ( 
.A(n_1732),
.B(n_1689),
.C(n_1712),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1724),
.B(n_1696),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1736),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1743),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1724),
.B(n_1696),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1747),
.Y(n_1763)
);

AO22x1_ASAP7_75t_L g1764 ( 
.A1(n_1730),
.A2(n_1710),
.B1(n_1709),
.B2(n_1720),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1749),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1735),
.A2(n_1709),
.B1(n_1708),
.B2(n_1704),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1727),
.A2(n_1734),
.B1(n_1748),
.B2(n_1738),
.C(n_1741),
.Y(n_1767)
);

O2A1O1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1742),
.A2(n_1721),
.B(n_1712),
.C(n_1719),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1725),
.B(n_1702),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1731),
.B(n_1702),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1750),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1757),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1756),
.B(n_1754),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1757),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1769),
.B(n_1733),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1751),
.A2(n_1740),
.B(n_1744),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1759),
.B(n_1737),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1755),
.A2(n_1695),
.B1(n_1714),
.B2(n_1716),
.C(n_1719),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1754),
.B(n_1710),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1758),
.B(n_1709),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1764),
.B(n_1704),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1752),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1772),
.Y(n_1783)
);

NAND3xp33_ASAP7_75t_L g1784 ( 
.A(n_1774),
.B(n_1753),
.C(n_1767),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1773),
.B(n_1762),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1780),
.A2(n_1695),
.B1(n_1763),
.B2(n_1765),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1775),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1773),
.B(n_1770),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1779),
.B(n_1766),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1771),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1781),
.B(n_1760),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1781),
.B(n_1768),
.Y(n_1792)
);

INVxp67_ASAP7_75t_L g1793 ( 
.A(n_1789),
.Y(n_1793)
);

OAI211xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1792),
.A2(n_1776),
.B(n_1780),
.C(n_1778),
.Y(n_1794)
);

AOI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1784),
.A2(n_1755),
.B1(n_1771),
.B2(n_1782),
.Y(n_1795)
);

NOR2x1_ASAP7_75t_L g1796 ( 
.A(n_1787),
.B(n_1782),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1788),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1797),
.B(n_1785),
.Y(n_1798)
);

AOI211xp5_ASAP7_75t_L g1799 ( 
.A1(n_1794),
.A2(n_1791),
.B(n_1783),
.C(n_1790),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1796),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1795),
.A2(n_1786),
.B1(n_1777),
.B2(n_1761),
.Y(n_1801)
);

AOI211xp5_ASAP7_75t_SL g1802 ( 
.A1(n_1793),
.A2(n_1786),
.B(n_1723),
.C(n_1720),
.Y(n_1802)
);

AOI211xp5_ASAP7_75t_L g1803 ( 
.A1(n_1794),
.A2(n_1721),
.B(n_1723),
.C(n_1705),
.Y(n_1803)
);

NAND2x1p5_ASAP7_75t_L g1804 ( 
.A(n_1800),
.B(n_1512),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1798),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1801),
.Y(n_1806)
);

INVxp67_ASAP7_75t_L g1807 ( 
.A(n_1802),
.Y(n_1807)
);

INVxp67_ASAP7_75t_SL g1808 ( 
.A(n_1799),
.Y(n_1808)
);

NAND4xp75_ASAP7_75t_L g1809 ( 
.A(n_1806),
.B(n_1803),
.C(n_1708),
.D(n_1705),
.Y(n_1809)
);

NOR2x1p5_ASAP7_75t_L g1810 ( 
.A(n_1805),
.B(n_1711),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_SL g1811 ( 
.A1(n_1807),
.A2(n_1716),
.B(n_1711),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1809),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1812),
.A2(n_1808),
.B1(n_1804),
.B2(n_1810),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1812),
.B1(n_1811),
.B2(n_1804),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1813),
.B(n_1675),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1814),
.A2(n_1815),
.B1(n_1714),
.B2(n_1713),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1815),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1817),
.A2(n_1666),
.B(n_1655),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1816),
.A2(n_1680),
.B1(n_1713),
.B2(n_1715),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1818),
.A2(n_1678),
.B(n_1677),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1820),
.B(n_1819),
.Y(n_1821)
);

XNOR2xp5_ASAP7_75t_L g1822 ( 
.A(n_1821),
.B(n_1715),
.Y(n_1822)
);

AOI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1822),
.A2(n_1687),
.B1(n_1678),
.B2(n_1677),
.Y(n_1823)
);

AOI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1823),
.A2(n_1510),
.B(n_1516),
.C(n_1511),
.Y(n_1824)
);


endmodule