module fake_netlist_6_2642_n_78 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_78);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_78;

wire n_52;
wire n_46;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_50;
wire n_49;
wire n_77;
wire n_42;
wire n_54;
wire n_32;
wire n_66;
wire n_47;
wire n_62;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_38;
wire n_61;
wire n_59;
wire n_76;
wire n_36;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_40;
wire n_41;
wire n_71;
wire n_74;
wire n_72;
wire n_60;
wire n_35;
wire n_69;
wire n_43;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_27),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_10),
.B(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_8),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_21),
.B(n_3),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_13),
.B(n_23),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

AND2x4_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_0),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

AND2x4_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_42),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_48),
.B1(n_39),
.B2(n_46),
.Y(n_59)
);

OAI21x1_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_47),
.B(n_37),
.Y(n_60)
);

AOI221xp5_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_36),
.B1(n_35),
.B2(n_32),
.C(n_45),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_9),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

AO21x2_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_50),
.B(n_55),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

AND2x4_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_61),
.B1(n_59),
.B2(n_69),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_58),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_69),
.B(n_66),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_65),
.B1(n_57),
.B2(n_68),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_56),
.C(n_0),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_74),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

AOI322xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_2),
.A3(n_4),
.B1(n_7),
.B2(n_16),
.C1(n_26),
.C2(n_28),
.Y(n_78)
);


endmodule