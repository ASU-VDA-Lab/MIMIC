module fake_jpeg_17898_n_353 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_12),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

AND2x4_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_47),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_51),
.Y(n_68)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_30),
.B1(n_23),
.B2(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_52),
.A2(n_65),
.B1(n_71),
.B2(n_26),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_54),
.B(n_55),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_23),
.B1(n_30),
.B2(n_31),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_34),
.B1(n_22),
.B2(n_29),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_70),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_35),
.B1(n_31),
.B2(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_32),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_49),
.B1(n_45),
.B2(n_48),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_18),
.B(n_17),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_18),
.B1(n_36),
.B2(n_17),
.Y(n_111)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_34),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_64),
.Y(n_84)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_50),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_74),
.B(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_79),
.B(n_83),
.Y(n_144)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_22),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_94),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_50),
.B1(n_44),
.B2(n_40),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_86),
.A2(n_36),
.B1(n_1),
.B2(n_2),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_89),
.B1(n_99),
.B2(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_96),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_26),
.B1(n_28),
.B2(n_34),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_90),
.B(n_92),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_29),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_20),
.Y(n_93)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_20),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_97),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_32),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_108),
.Y(n_122)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_17),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_73),
.A2(n_21),
.B1(n_16),
.B2(n_36),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_76),
.B1(n_69),
.B2(n_67),
.Y(n_136)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_59),
.A2(n_36),
.B1(n_14),
.B2(n_13),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_59),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_115),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_17),
.C(n_51),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_138),
.C(n_111),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_77),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_76),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_88),
.Y(n_134)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_141),
.B1(n_106),
.B2(n_104),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_85),
.B(n_18),
.C(n_27),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_69),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_86),
.Y(n_150)
);

AO22x1_ASAP7_75t_SL g145 ( 
.A1(n_107),
.A2(n_17),
.B1(n_27),
.B2(n_2),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_114),
.B1(n_105),
.B2(n_102),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_146),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_152),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_148),
.B(n_144),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_168),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_87),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_151),
.A2(n_165),
.B(n_170),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_146),
.Y(n_152)
);

AND2x4_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_90),
.Y(n_153)
);

AOI21x1_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_121),
.B(n_122),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_135),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_154),
.A2(n_133),
.B1(n_104),
.B2(n_118),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_158),
.Y(n_200)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_122),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_162),
.B1(n_129),
.B2(n_125),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_103),
.C(n_93),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_129),
.C(n_126),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_142),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_166),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_97),
.B1(n_100),
.B2(n_99),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_163),
.A2(n_179),
.B1(n_131),
.B2(n_119),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_91),
.Y(n_164)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_108),
.B(n_110),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_81),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_103),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_135),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_177),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_95),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_172),
.Y(n_180)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_83),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_144),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_120),
.B(n_80),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_176),
.A2(n_118),
.B1(n_80),
.B2(n_124),
.Y(n_195)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_127),
.A2(n_106),
.B1(n_113),
.B2(n_82),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_182),
.A2(n_186),
.B1(n_204),
.B2(n_206),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_183),
.A2(n_192),
.B(n_211),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_189),
.C(n_196),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_150),
.A2(n_141),
.B1(n_121),
.B2(n_145),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_188),
.A2(n_175),
.B1(n_163),
.B2(n_176),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_81),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_125),
.B(n_145),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_201),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_136),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_202),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_149),
.B(n_116),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_207),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_151),
.A2(n_124),
.B1(n_101),
.B2(n_133),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_151),
.A2(n_98),
.B1(n_123),
.B2(n_109),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_149),
.B(n_0),
.Y(n_209)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_153),
.A2(n_27),
.B(n_14),
.C(n_10),
.D(n_3),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_98),
.C(n_10),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_0),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_176),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_231),
.Y(n_253)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_197),
.B(n_168),
.CI(n_160),
.CON(n_215),
.SN(n_215)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_215),
.B(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_217),
.Y(n_261)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_177),
.Y(n_223)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_170),
.B1(n_152),
.B2(n_147),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_227),
.A2(n_239),
.B1(n_204),
.B2(n_180),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_195),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_182),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_161),
.B1(n_172),
.B2(n_174),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_194),
.B1(n_208),
.B2(n_209),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_191),
.B(n_193),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_170),
.B(n_156),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_186),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_189),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_236),
.C(n_187),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g235 ( 
.A1(n_203),
.A2(n_156),
.B(n_154),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_213),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_169),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_190),
.Y(n_238)
);

NAND3xp33_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_240),
.C(n_200),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_197),
.A2(n_167),
.B1(n_157),
.B2(n_171),
.Y(n_239)
);

NOR2x1_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_1),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_262),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_196),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_249),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_198),
.C(n_188),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_256),
.C(n_267),
.Y(n_268)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_225),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_255),
.B(n_266),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_219),
.Y(n_256)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_221),
.A2(n_202),
.B1(n_181),
.B2(n_210),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_264),
.A2(n_265),
.B1(n_240),
.B2(n_214),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_181),
.B1(n_210),
.B2(n_3),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_226),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_220),
.B(n_1),
.C(n_2),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_220),
.C(n_215),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_276),
.C(n_283),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_244),
.B(n_218),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_267),
.B(n_246),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_218),
.B1(n_214),
.B2(n_217),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_273),
.A2(n_278),
.B1(n_282),
.B2(n_4),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_257),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_285),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_215),
.C(n_227),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_214),
.B1(n_231),
.B2(n_235),
.Y(n_278)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_233),
.B1(n_232),
.B2(n_3),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_1),
.C(n_2),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_3),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_247),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_4),
.Y(n_302)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_243),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_284),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_283),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_248),
.C(n_263),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_295),
.C(n_303),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_251),
.B1(n_264),
.B2(n_254),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_305),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_259),
.C(n_258),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_297),
.B(n_300),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_273),
.A2(n_265),
.B(n_260),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_297),
.A2(n_300),
.B(n_306),
.Y(n_314)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_4),
.B(n_5),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_282),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_5),
.C(n_6),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_304)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_274),
.A2(n_271),
.B1(n_270),
.B2(n_279),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_277),
.A2(n_6),
.B(n_7),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_302),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_309),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_284),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_321),
.C(n_290),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_313),
.A2(n_292),
.B(n_296),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_318),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_291),
.B(n_286),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_316),
.B(n_320),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_8),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_295),
.B(n_288),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_290),
.B(n_288),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_327),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_328),
.C(n_332),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_303),
.Y(n_325)
);

OAI211xp5_ASAP7_75t_L g340 ( 
.A1(n_325),
.A2(n_326),
.B(n_314),
.C(n_308),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_305),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_310),
.A2(n_9),
.B1(n_294),
.B2(n_319),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_9),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_329),
.B(n_309),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_9),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_334),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_312),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_338),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_312),
.Y(n_338)
);

AOI21x1_ASAP7_75t_L g339 ( 
.A1(n_324),
.A2(n_317),
.B(n_314),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_339),
.A2(n_340),
.B1(n_324),
.B2(n_317),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_331),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_342),
.B(n_344),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_322),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_340),
.C(n_334),
.Y(n_348)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_345),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_346),
.Y(n_349)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_349),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_344),
.Y(n_351)
);

OAI211xp5_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_347),
.B(n_348),
.C(n_341),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_343),
.Y(n_353)
);


endmodule