module fake_jpeg_22638_n_225 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_15),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_37),
.Y(n_73)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_42),
.B(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_0),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_20),
.C(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_50),
.B(n_55),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_19),
.B1(n_33),
.B2(n_20),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_63),
.B1(n_21),
.B2(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_74),
.Y(n_82)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_65),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_16),
.B1(n_34),
.B2(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_36),
.A2(n_19),
.B1(n_16),
.B2(n_34),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_17),
.B1(n_20),
.B2(n_33),
.Y(n_88)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_44),
.B1(n_38),
.B2(n_19),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_23),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_30),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_98),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_64),
.B1(n_71),
.B2(n_29),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_85),
.A2(n_86),
.B1(n_96),
.B2(n_104),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_33),
.B1(n_20),
.B2(n_43),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_89),
.B1(n_26),
.B2(n_2),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_23),
.B1(n_28),
.B2(n_30),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_30),
.B1(n_28),
.B2(n_40),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_37),
.B(n_35),
.C(n_3),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_71),
.B(n_35),
.C(n_29),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_79),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_105),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_70),
.B1(n_68),
.B2(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_26),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_35),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_26),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_66),
.C(n_73),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_126),
.C(n_93),
.Y(n_147)
);

AO22x1_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_59),
.B1(n_60),
.B2(n_54),
.Y(n_111)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_122),
.B(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_113),
.Y(n_153)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_1),
.Y(n_114)
);

XOR2x1_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_116),
.Y(n_160)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_118),
.Y(n_158)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

AO22x2_ASAP7_75t_L g121 ( 
.A1(n_81),
.A2(n_60),
.B1(n_62),
.B2(n_67),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_111),
.B1(n_130),
.B2(n_108),
.Y(n_150)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_96),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_87),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_123),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_130),
.B1(n_131),
.B2(n_99),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_64),
.C(n_29),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_29),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_95),
.Y(n_144)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_129),
.B(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_94),
.A2(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_102),
.B(n_106),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_122),
.A2(n_129),
.B1(n_121),
.B2(n_116),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_146),
.B1(n_155),
.B2(n_121),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_135),
.B1(n_117),
.B2(n_3),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_141),
.B(n_115),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_114),
.B(n_95),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_120),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_108),
.B1(n_102),
.B2(n_92),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_152),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_95),
.B(n_93),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_156),
.B(n_121),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_154),
.B1(n_157),
.B2(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_114),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_91),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_84),
.B(n_1),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_84),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_151),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_166),
.B1(n_170),
.B2(n_172),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_143),
.Y(n_178)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_171),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_115),
.A3(n_127),
.B1(n_1),
.B2(n_4),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_6),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_113),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_173),
.A2(n_155),
.B1(n_154),
.B2(n_138),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_142),
.C(n_149),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_6),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_145),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_185),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_162),
.B(n_140),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_189),
.C(n_167),
.Y(n_190)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_184),
.Y(n_196)
);

OAI322xp33_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_159),
.A3(n_152),
.B1(n_148),
.B2(n_147),
.C1(n_138),
.C2(n_156),
.Y(n_183)
);

OA21x2_ASAP7_75t_SL g191 ( 
.A1(n_183),
.A2(n_167),
.B(n_169),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_150),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_187),
.A2(n_172),
.B1(n_170),
.B2(n_175),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_193),
.C(n_198),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_191),
.B(n_178),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_197),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_174),
.C(n_165),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_182),
.A2(n_173),
.B1(n_142),
.B2(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_161),
.C(n_12),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_10),
.C(n_13),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_201),
.Y(n_204)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_190),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_196),
.A2(n_187),
.B(n_180),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_207),
.B(n_200),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_196),
.A2(n_177),
.B(n_186),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_10),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_208),
.B(n_13),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_203),
.A2(n_194),
.B1(n_193),
.B2(n_199),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_211),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_198),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_206),
.C(n_13),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_207),
.B(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_213),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_217),
.C(n_216),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_15),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_218),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_220),
.B(n_15),
.Y(n_224)
);


endmodule