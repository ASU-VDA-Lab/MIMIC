module real_jpeg_1291_n_7 (n_5, n_4, n_0, n_1, n_2, n_6, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_57;
wire n_43;
wire n_37;
wire n_21;
wire n_54;
wire n_65;
wire n_33;
wire n_35;
wire n_50;
wire n_38;
wire n_29;
wire n_55;
wire n_58;
wire n_10;
wire n_31;
wire n_9;
wire n_49;
wire n_52;
wire n_67;
wire n_63;
wire n_12;
wire n_24;
wire n_66;
wire n_34;
wire n_28;
wire n_60;
wire n_44;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_51;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_56;
wire n_30;
wire n_48;
wire n_16;
wire n_15;
wire n_13;

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_2),
.B(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_2),
.A2(n_12),
.B1(n_22),
.B2(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_2),
.B(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_2),
.A2(n_26),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_2),
.B(n_12),
.C(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_2),
.B(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_3),
.A2(n_12),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_3),
.A2(n_21),
.B1(n_40),
.B2(n_41),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_51),
.Y(n_7)
);

OAI21xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_34),
.B(n_50),
.Y(n_8)
);

AOI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_27),
.B(n_33),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_17),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_15),
.Y(n_11)
);

INVx3_ASAP7_75t_SL g22 ( 
.A(n_12),
.Y(n_22)
);

AO22x1_ASAP7_75t_SL g29 ( 
.A1(n_12),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_22),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_16),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

OA21x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B(n_23),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_32),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_31),
.B1(n_40),
.B2(n_41),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_32),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_39),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_65)
);

AOI22x1_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_41),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_67),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);


endmodule