module fake_netlist_6_791_n_2305 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2305);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2305;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_343;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_2292;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_1093;
wire n_418;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_1098;
wire n_391;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_SL g219 ( 
.A(n_27),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_191),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_36),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_207),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_205),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_68),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_61),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_159),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_201),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_120),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_78),
.Y(n_231)
);

BUFx2_ASAP7_75t_SL g232 ( 
.A(n_122),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_47),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_22),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_151),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_187),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_92),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_138),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_165),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_184),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_50),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_166),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_128),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_127),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_82),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_19),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_88),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_124),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_176),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_107),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_170),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_143),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_188),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_9),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_135),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_83),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_32),
.Y(n_258)
);

BUFx2_ASAP7_75t_SL g259 ( 
.A(n_137),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_3),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_103),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_68),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_95),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_18),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_161),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_82),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_139),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_160),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_164),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_28),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_76),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_131),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_55),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_35),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_154),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_60),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_198),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_216),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_60),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_40),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_209),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_42),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_47),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_152),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_63),
.Y(n_285)
);

BUFx2_ASAP7_75t_SL g286 ( 
.A(n_93),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_113),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_54),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_5),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_142),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_133),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_145),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_3),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_130),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_157),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_202),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_25),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_185),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_55),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_97),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_98),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_79),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_109),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_48),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_200),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_210),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_50),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_29),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_45),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_146),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_79),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_203),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_57),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_11),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_118),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_192),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_66),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_168),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_92),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_58),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_17),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_12),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_132),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_95),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_80),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_116),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_62),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_18),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_104),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_171),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_134),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_28),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_1),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_156),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_24),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_175),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_93),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_36),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_101),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_172),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_52),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_27),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_33),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_52),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_25),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_10),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_86),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_70),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_162),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_62),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_64),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_67),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_206),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_80),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_29),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_181),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_105),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_106),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_14),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_63),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_33),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_37),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_111),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_19),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_196),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_147),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_99),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_11),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_149),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_101),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_40),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_148),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_123),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_114),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_66),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_88),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_70),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_194),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_17),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_208),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_98),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_197),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_10),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_41),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_144),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_61),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_14),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_57),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_4),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_77),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_12),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_38),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_71),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_0),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_7),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_110),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_32),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_38),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_94),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_126),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_15),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_15),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_179),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_215),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_72),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_212),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_87),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_180),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_35),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_87),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_43),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_51),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_31),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_59),
.Y(n_415)
);

BUFx10_ASAP7_75t_L g416 ( 
.A(n_217),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_136),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_81),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_96),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_218),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_65),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_1),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_39),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_96),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_64),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_99),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_5),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_0),
.Y(n_428)
);

INVxp33_ASAP7_75t_L g429 ( 
.A(n_42),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_155),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_233),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_220),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_222),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_251),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_223),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_233),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_233),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_233),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_233),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_231),
.B(n_2),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_233),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_227),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_229),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_256),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_256),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_253),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_246),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_246),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_246),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_246),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_246),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_246),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_230),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_236),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_241),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_238),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_413),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_413),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_413),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_319),
.B(n_2),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_413),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_358),
.B(n_4),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_267),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_239),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_358),
.B(n_6),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_240),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_281),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_383),
.B(n_6),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_242),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_383),
.B(n_7),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_413),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_366),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_373),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_243),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_413),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_342),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_273),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_249),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_250),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_342),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_420),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_252),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_255),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_256),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_342),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_330),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_269),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_419),
.Y(n_488)
);

NOR2xp67_ASAP7_75t_L g489 ( 
.A(n_319),
.B(n_8),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_299),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_419),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_419),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_282),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_282),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_299),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_241),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_330),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_268),
.Y(n_498)
);

BUFx2_ASAP7_75t_SL g499 ( 
.A(n_354),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_282),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_399),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_399),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_399),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_231),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_272),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_247),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_277),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_247),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_260),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_354),
.B(n_8),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_260),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_284),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_274),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_248),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_274),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_287),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_280),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_280),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_319),
.B(n_9),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_289),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_289),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_291),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_294),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_300),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_308),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_300),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_248),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_295),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_304),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_309),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_309),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_299),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_318),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_318),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_329),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_329),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_324),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_340),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_331),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_335),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_322),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_322),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_340),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_225),
.B(n_228),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_444),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_487),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_487),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_432),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_460),
.B(n_308),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_450),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_487),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_489),
.B(n_328),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_484),
.B(n_306),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_450),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_496),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_490),
.B(n_219),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_433),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_450),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_431),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_435),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_431),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_434),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_446),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_519),
.B(n_219),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_436),
.B(n_306),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_436),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_487),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_495),
.B(n_219),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_542),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_532),
.B(n_293),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_442),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_486),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_463),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_487),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_437),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_514),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_437),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_438),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_438),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_443),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_453),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_514),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_444),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_454),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_499),
.B(n_429),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_439),
.B(n_306),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_439),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_441),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_445),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g590 ( 
.A(n_476),
.B(n_319),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_456),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_464),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_441),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_447),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_447),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_466),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_469),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_474),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_497),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_499),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_525),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_544),
.B(n_293),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_448),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_448),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_L g605 ( 
.A(n_440),
.B(n_293),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_478),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_449),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_510),
.B(n_493),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_449),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_451),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_451),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_527),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_479),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_452),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_482),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_527),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_445),
.B(n_314),
.Y(n_617)
);

BUFx8_ASAP7_75t_L g618 ( 
.A(n_440),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_452),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_483),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_493),
.B(n_430),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_457),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_467),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_494),
.B(n_341),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_472),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_498),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_455),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_457),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_458),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_507),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_494),
.B(n_350),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_458),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_459),
.B(n_248),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_473),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_600),
.B(n_500),
.Y(n_635)
);

INVxp67_ASAP7_75t_SL g636 ( 
.A(n_589),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_569),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_553),
.B(n_512),
.Y(n_638)
);

INVxp33_ASAP7_75t_L g639 ( 
.A(n_627),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_569),
.B(n_541),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_575),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_600),
.B(n_516),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_585),
.B(n_522),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_553),
.B(n_500),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_575),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_605),
.A2(n_477),
.B1(n_465),
.B2(n_468),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_559),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_559),
.Y(n_648)
);

NOR2x1p5_ASAP7_75t_L g649 ( 
.A(n_548),
.B(n_344),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_561),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_583),
.B(n_523),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_561),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_617),
.B(n_501),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_553),
.B(n_501),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_575),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_566),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_565),
.B(n_225),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_608),
.B(n_539),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_545),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_608),
.B(n_459),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_566),
.Y(n_661)
);

CKINVDCx16_ASAP7_75t_R g662 ( 
.A(n_601),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_577),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_583),
.B(n_505),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_577),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_587),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_565),
.B(n_586),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_578),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_545),
.B(n_528),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_545),
.B(n_529),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_587),
.Y(n_671)
);

BUFx4f_ASAP7_75t_L g672 ( 
.A(n_633),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_549),
.B(n_537),
.Y(n_673)
);

NAND3x1_ASAP7_75t_L g674 ( 
.A(n_585),
.B(n_470),
.C(n_462),
.Y(n_674)
);

NAND2x1p5_ASAP7_75t_L g675 ( 
.A(n_633),
.B(n_275),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_565),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_578),
.Y(n_677)
);

CKINVDCx8_ASAP7_75t_R g678 ( 
.A(n_601),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_578),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_594),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_594),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_589),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_602),
.B(n_502),
.Y(n_683)
);

OAI221xp5_ASAP7_75t_L g684 ( 
.A1(n_602),
.A2(n_314),
.B1(n_349),
.B2(n_320),
.C(n_345),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_604),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_551),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_621),
.B(n_624),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_582),
.Y(n_688)
);

INVxp67_ASAP7_75t_SL g689 ( 
.A(n_546),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_557),
.B(n_540),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_549),
.B(n_502),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_552),
.A2(n_328),
.B1(n_410),
.B2(n_376),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_556),
.B(n_503),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_551),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_582),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_551),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_551),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_605),
.A2(n_410),
.B1(n_263),
.B2(n_283),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_624),
.B(n_631),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_560),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_564),
.A2(n_349),
.B1(n_320),
.B2(n_344),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_604),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_SL g703 ( 
.A(n_571),
.B(n_481),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_582),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_552),
.B(n_503),
.Y(n_705)
);

BUFx6f_ASAP7_75t_SL g706 ( 
.A(n_565),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_546),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_580),
.B(n_235),
.Y(n_708)
);

AND2x6_ASAP7_75t_L g709 ( 
.A(n_633),
.B(n_265),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_565),
.B(n_228),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_581),
.B(n_275),
.Y(n_711)
);

BUFx4f_ASAP7_75t_L g712 ( 
.A(n_633),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_551),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_584),
.B(n_296),
.Y(n_714)
);

OAI21xp33_ASAP7_75t_SL g715 ( 
.A1(n_556),
.A2(n_362),
.B(n_355),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_591),
.B(n_235),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_579),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_631),
.B(n_461),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_607),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_627),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_586),
.B(n_471),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_592),
.B(n_296),
.Y(n_722)
);

NAND3x1_ASAP7_75t_L g723 ( 
.A(n_568),
.B(n_362),
.C(n_355),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_596),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_607),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_579),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_586),
.B(n_261),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_611),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_579),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_568),
.B(n_476),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_551),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_588),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_551),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_586),
.B(n_261),
.Y(n_734)
);

INVx6_ASAP7_75t_L g735 ( 
.A(n_586),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_546),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_588),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_617),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_582),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_546),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_R g741 ( 
.A(n_597),
.B(n_598),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_570),
.B(n_480),
.Y(n_742)
);

XNOR2xp5_ASAP7_75t_L g743 ( 
.A(n_634),
.B(n_226),
.Y(n_743)
);

OR2x6_ASAP7_75t_L g744 ( 
.A(n_570),
.B(n_232),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_606),
.B(n_235),
.Y(n_745)
);

AND2x6_ASAP7_75t_L g746 ( 
.A(n_633),
.B(n_265),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_588),
.Y(n_747)
);

INVx5_ASAP7_75t_L g748 ( 
.A(n_582),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_617),
.B(n_480),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_582),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_550),
.B(n_471),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_546),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_611),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_593),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_564),
.A2(n_377),
.B1(n_380),
.B2(n_365),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_590),
.B(n_290),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_618),
.A2(n_377),
.B1(n_380),
.B2(n_365),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_593),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_614),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_555),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_614),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_547),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_593),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_582),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_618),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_555),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_613),
.B(n_235),
.Y(n_767)
);

AND2x2_ASAP7_75t_SL g768 ( 
.A(n_626),
.B(n_265),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_615),
.B(n_221),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_622),
.B(n_485),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_620),
.B(n_244),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_599),
.B(n_369),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_595),
.Y(n_773)
);

BUFx10_ASAP7_75t_L g774 ( 
.A(n_550),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_562),
.Y(n_775)
);

INVx5_ASAP7_75t_L g776 ( 
.A(n_612),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_626),
.B(n_232),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_595),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_595),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_603),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_618),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_603),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_630),
.B(n_244),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_603),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_622),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_609),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_609),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_687),
.B(n_699),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_647),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_642),
.B(n_630),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_768),
.B(n_618),
.Y(n_791)
);

INVx8_ASAP7_75t_L g792 ( 
.A(n_706),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_676),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_768),
.B(n_658),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_711),
.B(n_618),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_768),
.B(n_357),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_691),
.A2(n_292),
.B(n_337),
.C(n_297),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_660),
.B(n_616),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_738),
.B(n_364),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_637),
.Y(n_800)
);

OR2x6_ASAP7_75t_L g801 ( 
.A(n_781),
.B(n_259),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_683),
.B(n_616),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_738),
.B(n_367),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_714),
.B(n_599),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_637),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_635),
.B(n_370),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_683),
.B(n_616),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_676),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_SL g809 ( 
.A(n_765),
.B(n_244),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_647),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_705),
.B(n_337),
.C(n_292),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_635),
.B(n_375),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_718),
.B(n_616),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_730),
.B(n_629),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_L g815 ( 
.A1(n_698),
.A2(n_744),
.B1(n_638),
.B2(n_777),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_674),
.A2(n_644),
.B1(n_654),
.B2(n_723),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_730),
.B(n_629),
.Y(n_817)
);

NOR2xp67_ASAP7_75t_L g818 ( 
.A(n_659),
.B(n_667),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_648),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_676),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_657),
.A2(n_292),
.B(n_337),
.C(n_297),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_674),
.A2(n_325),
.B1(n_346),
.B2(n_302),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_742),
.B(n_632),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_722),
.B(n_639),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_SL g825 ( 
.A(n_700),
.B(n_623),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_651),
.B(n_623),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_648),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_643),
.B(n_572),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_742),
.B(n_632),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_739),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_657),
.A2(n_307),
.B1(n_311),
.B2(n_290),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_659),
.B(n_307),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_769),
.B(n_562),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_657),
.A2(n_313),
.B1(n_317),
.B2(n_311),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_693),
.B(n_554),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_650),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_682),
.B(n_386),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_682),
.B(n_397),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_640),
.B(n_563),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_693),
.B(n_554),
.Y(n_840)
);

BUFx8_ASAP7_75t_L g841 ( 
.A(n_765),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_650),
.Y(n_842)
);

OAI22xp33_ASAP7_75t_L g843 ( 
.A1(n_698),
.A2(n_313),
.B1(n_327),
.B2(n_317),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_644),
.B(n_558),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_654),
.B(n_558),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_640),
.B(n_563),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_657),
.A2(n_332),
.B1(n_374),
.B2(n_327),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_652),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_667),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_636),
.B(n_573),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_652),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_675),
.B(n_619),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_772),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_675),
.B(n_619),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_720),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_646),
.B(n_401),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_673),
.B(n_404),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_675),
.B(n_656),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_723),
.A2(n_384),
.B1(n_388),
.B2(n_372),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_656),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_661),
.B(n_663),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_661),
.B(n_619),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_757),
.A2(n_332),
.B1(n_379),
.B2(n_374),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_663),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_L g865 ( 
.A(n_710),
.B(n_381),
.C(n_379),
.Y(n_865)
);

NAND2x1_ASAP7_75t_L g866 ( 
.A(n_735),
.B(n_619),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_760),
.B(n_573),
.Y(n_867)
);

NOR2x2_ASAP7_75t_L g868 ( 
.A(n_777),
.B(n_408),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_672),
.A2(n_574),
.B(n_567),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_665),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_664),
.B(n_405),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_772),
.B(n_369),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_766),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_665),
.Y(n_874)
);

INVxp67_ASAP7_75t_SL g875 ( 
.A(n_739),
.Y(n_875)
);

INVx8_ASAP7_75t_L g876 ( 
.A(n_706),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_666),
.B(n_619),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_666),
.B(n_628),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_667),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_671),
.B(n_628),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_667),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_781),
.B(n_407),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_671),
.B(n_628),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_680),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_735),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_775),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_692),
.B(n_409),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_653),
.B(n_244),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_680),
.B(n_628),
.Y(n_889)
);

OR2x6_ASAP7_75t_L g890 ( 
.A(n_777),
.B(n_259),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_681),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_681),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_653),
.B(n_278),
.Y(n_893)
);

O2A1O1Ixp5_ASAP7_75t_L g894 ( 
.A1(n_710),
.A2(n_628),
.B(n_574),
.C(n_417),
.Y(n_894)
);

AND2x6_ASAP7_75t_SL g895 ( 
.A(n_777),
.B(n_385),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_749),
.B(n_504),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_669),
.B(n_278),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_783),
.B(n_625),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_685),
.B(n_547),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_672),
.A2(n_574),
.B(n_590),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_670),
.B(n_625),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_685),
.B(n_547),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_702),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_702),
.B(n_547),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_710),
.A2(n_417),
.B1(n_381),
.B2(n_286),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_SL g906 ( 
.A(n_777),
.B(n_278),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_708),
.B(n_634),
.Y(n_907)
);

NAND2x1_ASAP7_75t_L g908 ( 
.A(n_735),
.B(n_547),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_749),
.Y(n_909)
);

AOI221xp5_ASAP7_75t_L g910 ( 
.A1(n_684),
.A2(n_400),
.B1(n_376),
.B2(n_411),
.C(n_414),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_741),
.B(n_278),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_735),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_719),
.B(n_567),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_715),
.A2(n_286),
.B1(n_270),
.B2(n_411),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_715),
.A2(n_270),
.B(n_414),
.C(n_475),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_774),
.B(n_416),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_743),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_710),
.A2(n_269),
.B1(n_316),
.B2(n_359),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_719),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_716),
.B(n_745),
.Y(n_920)
);

NAND2xp33_ASAP7_75t_L g921 ( 
.A(n_709),
.B(n_269),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_725),
.B(n_567),
.Y(n_922)
);

NOR2xp67_ASAP7_75t_L g923 ( 
.A(n_721),
.B(n_475),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_725),
.B(n_567),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_767),
.B(n_400),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_727),
.A2(n_269),
.B1(n_316),
.B2(n_359),
.Y(n_926)
);

NOR2xp67_ASAP7_75t_L g927 ( 
.A(n_751),
.B(n_567),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_771),
.B(n_224),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_727),
.A2(n_269),
.B1(n_316),
.B2(n_359),
.Y(n_929)
);

NOR3xp33_ASAP7_75t_L g930 ( 
.A(n_662),
.B(n_237),
.C(n_234),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_728),
.Y(n_931)
);

AND3x1_ASAP7_75t_L g932 ( 
.A(n_701),
.B(n_387),
.C(n_385),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_727),
.A2(n_279),
.B1(n_315),
.B2(n_312),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_SL g934 ( 
.A1(n_764),
.A2(n_576),
.B(n_610),
.C(n_609),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_728),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_744),
.B(n_504),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_744),
.B(n_506),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_672),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_753),
.B(n_612),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_774),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_774),
.B(n_416),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_774),
.B(n_416),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_727),
.A2(n_269),
.B1(n_316),
.B2(n_359),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_744),
.A2(n_387),
.B(n_424),
.C(n_415),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_753),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_736),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_759),
.B(n_612),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_734),
.A2(n_316),
.B1(n_359),
.B2(n_610),
.Y(n_948)
);

BUFx8_ASAP7_75t_L g949 ( 
.A(n_706),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_759),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_761),
.B(n_612),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_761),
.B(n_612),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_712),
.B(n_700),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_734),
.A2(n_316),
.B1(n_359),
.B2(n_610),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_785),
.B(n_612),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_785),
.B(n_612),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_712),
.B(n_416),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_734),
.B(n_576),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_789),
.Y(n_959)
);

NAND2x1p5_ASAP7_75t_L g960 ( 
.A(n_938),
.B(n_712),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_789),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_792),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_900),
.A2(n_707),
.B(n_689),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_788),
.A2(n_734),
.B1(n_649),
.B2(n_744),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_810),
.Y(n_965)
);

OR2x6_ASAP7_75t_L g966 ( 
.A(n_792),
.B(n_690),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_824),
.B(n_700),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_SL g968 ( 
.A(n_843),
.B(n_662),
.C(n_743),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_792),
.B(n_649),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_909),
.B(n_842),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_792),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_885),
.B(n_736),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_949),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_810),
.Y(n_974)
);

INVxp67_ASAP7_75t_SL g975 ( 
.A(n_946),
.Y(n_975)
);

AO22x1_ASAP7_75t_L g976 ( 
.A1(n_795),
.A2(n_746),
.B1(n_709),
.B2(n_756),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_909),
.B(n_770),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_819),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_SL g979 ( 
.A(n_839),
.B(n_254),
.C(n_245),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_819),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_827),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_827),
.Y(n_982)
);

INVx5_ASAP7_75t_L g983 ( 
.A(n_881),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_881),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_842),
.B(n_770),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_805),
.Y(n_986)
);

NOR3xp33_ASAP7_75t_SL g987 ( 
.A(n_846),
.B(n_258),
.C(n_257),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_805),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_800),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_896),
.B(n_700),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_SL g991 ( 
.A(n_867),
.B(n_264),
.C(n_262),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_836),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_851),
.B(n_736),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_836),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_802),
.A2(n_746),
.B(n_709),
.Y(n_995)
);

BUFx4_ASAP7_75t_SL g996 ( 
.A(n_895),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_848),
.Y(n_997)
);

AND2x6_ASAP7_75t_L g998 ( 
.A(n_881),
.B(n_756),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_876),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_848),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_R g1001 ( 
.A(n_825),
.B(n_703),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_864),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_864),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_851),
.B(n_740),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_881),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_870),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_860),
.B(n_740),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_870),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_860),
.B(n_740),
.Y(n_1009)
);

NOR3xp33_ASAP7_75t_SL g1010 ( 
.A(n_850),
.B(n_271),
.C(n_266),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_884),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_874),
.B(n_752),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_874),
.B(n_752),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_855),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_881),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_855),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_896),
.B(n_724),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_853),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_891),
.B(n_752),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_884),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_885),
.B(n_762),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_790),
.B(n_724),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_892),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_892),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_849),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_894),
.A2(n_764),
.B(n_733),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_931),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_931),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_SL g1029 ( 
.A(n_886),
.B(n_724),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_935),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_938),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_872),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_935),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_804),
.B(n_678),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_873),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_936),
.B(n_724),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_SL g1037 ( 
.A(n_925),
.B(n_285),
.C(n_276),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_945),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_849),
.Y(n_1039)
);

NOR2x1_ASAP7_75t_L g1040 ( 
.A(n_940),
.B(n_762),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_891),
.B(n_762),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_936),
.B(n_678),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_794),
.A2(n_709),
.B1(n_746),
.B2(n_756),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_938),
.B(n_756),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_849),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_937),
.B(n_755),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_903),
.B(n_709),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_937),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_872),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_879),
.Y(n_1050)
);

NAND2xp33_ASAP7_75t_SL g1051 ( 
.A(n_791),
.B(n_938),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_SL g1052 ( 
.A(n_938),
.B(n_694),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_949),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_879),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_945),
.Y(n_1055)
);

NOR2x1_ASAP7_75t_L g1056 ( 
.A(n_940),
.B(n_686),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_950),
.Y(n_1057)
);

NAND2xp33_ASAP7_75t_SL g1058 ( 
.A(n_953),
.B(n_694),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_879),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_832),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_815),
.A2(n_746),
.B1(n_709),
.B2(n_645),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_793),
.B(n_709),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_903),
.B(n_746),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_793),
.B(n_746),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_832),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_832),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_876),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_950),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_808),
.B(n_746),
.Y(n_1069)
);

BUFx4f_ASAP7_75t_L g1070 ( 
.A(n_876),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_826),
.B(n_920),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_917),
.B(n_506),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_828),
.B(n_288),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_808),
.B(n_764),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_919),
.B(n_686),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_SL g1076 ( 
.A(n_898),
.B(n_301),
.C(n_298),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_919),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_R g1078 ( 
.A(n_876),
.B(n_906),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_833),
.B(n_303),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_R g1080 ( 
.A(n_906),
.B(n_686),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_835),
.B(n_645),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_814),
.B(n_686),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_820),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_820),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_958),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_840),
.B(n_655),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_912),
.B(n_764),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_946),
.Y(n_1088)
);

INVx4_ASAP7_75t_L g1089 ( 
.A(n_912),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_949),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_946),
.Y(n_1091)
);

CKINVDCx6p67_ASAP7_75t_R g1092 ( 
.A(n_890),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_871),
.B(n_305),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_858),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_912),
.B(n_733),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_868),
.Y(n_1096)
);

INVxp67_ASAP7_75t_SL g1097 ( 
.A(n_818),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_SL g1098 ( 
.A(n_910),
.B(n_321),
.C(n_310),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_862),
.Y(n_1099)
);

AO22x1_ASAP7_75t_L g1100 ( 
.A1(n_863),
.A2(n_396),
.B1(n_415),
.B2(n_424),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_796),
.A2(n_747),
.B(n_668),
.C(n_677),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_901),
.B(n_323),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_877),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_R g1104 ( 
.A(n_809),
.B(n_733),
.Y(n_1104)
);

NAND2xp33_ASAP7_75t_R g1105 ( 
.A(n_907),
.B(n_326),
.Y(n_1105)
);

INVx5_ASAP7_75t_L g1106 ( 
.A(n_890),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_816),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_841),
.Y(n_1108)
);

OAI21xp33_ASAP7_75t_SL g1109 ( 
.A1(n_816),
.A2(n_861),
.B(n_823),
.Y(n_1109)
);

NOR3xp33_ASAP7_75t_SL g1110 ( 
.A(n_888),
.B(n_334),
.C(n_333),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_878),
.Y(n_1111)
);

BUFx8_ASAP7_75t_L g1112 ( 
.A(n_841),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_880),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_890),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_866),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_883),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_889),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_939),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_817),
.B(n_733),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_829),
.B(n_655),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_807),
.A2(n_729),
.B1(n_668),
.B2(n_677),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_947),
.Y(n_1122)
);

OR2x6_ASAP7_75t_L g1123 ( 
.A(n_890),
.B(n_508),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_899),
.Y(n_1124)
);

BUFx12f_ASAP7_75t_L g1125 ( 
.A(n_841),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_SL g1126 ( 
.A(n_809),
.B(n_421),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_856),
.A2(n_747),
.B1(n_679),
.B2(n_726),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_844),
.B(n_679),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_845),
.B(n_726),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_902),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_933),
.B(n_729),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_908),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_908),
.Y(n_1133)
);

NOR3xp33_ASAP7_75t_SL g1134 ( 
.A(n_893),
.B(n_338),
.C(n_336),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_904),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_818),
.B(n_754),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_913),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_866),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_951),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_952),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_933),
.B(n_928),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_955),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_956),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_868),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_852),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_922),
.Y(n_1146)
);

NOR3xp33_ASAP7_75t_SL g1147 ( 
.A(n_837),
.B(n_343),
.C(n_339),
.Y(n_1147)
);

NOR3xp33_ASAP7_75t_SL g1148 ( 
.A(n_838),
.B(n_348),
.C(n_347),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_806),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_895),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_798),
.B(n_754),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_963),
.A2(n_921),
.B(n_854),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1071),
.B(n_812),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1073),
.B(n_857),
.Y(n_1154)
);

BUFx8_ASAP7_75t_L g1155 ( 
.A(n_1125),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1026),
.A2(n_869),
.B(n_924),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1094),
.B(n_813),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_SL g1158 ( 
.A1(n_1094),
.A2(n_944),
.B(n_915),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_1107),
.A2(n_797),
.A3(n_821),
.B(n_717),
.Y(n_1159)
);

OAI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1126),
.A2(n_822),
.B1(n_859),
.B2(n_801),
.Y(n_1160)
);

OAI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_1079),
.A2(n_822),
.B(n_859),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_959),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_965),
.Y(n_1163)
);

INVxp67_ASAP7_75t_L g1164 ( 
.A(n_1014),
.Y(n_1164)
);

AOI21xp33_ASAP7_75t_L g1165 ( 
.A1(n_1102),
.A2(n_887),
.B(n_897),
.Y(n_1165)
);

OA22x2_ASAP7_75t_L g1166 ( 
.A1(n_1107),
.A2(n_914),
.B1(n_801),
.B2(n_941),
.Y(n_1166)
);

NOR2x1_ASAP7_75t_R g1167 ( 
.A(n_1125),
.B(n_911),
.Y(n_1167)
);

AOI31xp67_ASAP7_75t_L g1168 ( 
.A1(n_959),
.A2(n_961),
.A3(n_978),
.B(n_974),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_977),
.B(n_970),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_990),
.B(n_905),
.Y(n_1170)
);

BUFx4f_ASAP7_75t_L g1171 ( 
.A(n_1067),
.Y(n_1171)
);

AND3x2_ASAP7_75t_L g1172 ( 
.A(n_1034),
.B(n_930),
.C(n_428),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_990),
.B(n_831),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1017),
.B(n_834),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1026),
.A2(n_960),
.B(n_1101),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1017),
.B(n_916),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_960),
.A2(n_875),
.B(n_830),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_SL g1178 ( 
.A1(n_1145),
.A2(n_914),
.B(n_847),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_960),
.A2(n_811),
.B(n_957),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1075),
.A2(n_811),
.B(n_865),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_SL g1181 ( 
.A(n_1029),
.B(n_801),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1141),
.A2(n_942),
.B1(n_882),
.B2(n_803),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1001),
.B(n_799),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_983),
.B(n_1031),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1089),
.Y(n_1185)
);

AOI221x1_ASAP7_75t_L g1186 ( 
.A1(n_1051),
.A2(n_865),
.B1(n_758),
.B2(n_779),
.C(n_773),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_961),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_993),
.A2(n_927),
.B(n_923),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_983),
.B(n_688),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1046),
.B(n_932),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1081),
.B(n_948),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1109),
.A2(n_964),
.B(n_1093),
.C(n_1085),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1004),
.A2(n_927),
.B(n_923),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1014),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1081),
.B(n_954),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1007),
.A2(n_926),
.B(n_918),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1085),
.A2(n_921),
.B(n_929),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_974),
.Y(n_1198)
);

NOR2xp67_ASAP7_75t_L g1199 ( 
.A(n_1032),
.B(n_108),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1060),
.A2(n_801),
.B1(n_943),
.B2(n_932),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_978),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_989),
.B(n_351),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1009),
.A2(n_717),
.B(n_641),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_1112),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_995),
.A2(n_695),
.B(n_688),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1082),
.A2(n_934),
.B(n_773),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1151),
.A2(n_695),
.B(n_688),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1012),
.A2(n_717),
.B(n_641),
.Y(n_1208)
);

AOI21xp33_ASAP7_75t_L g1209 ( 
.A1(n_1105),
.A2(n_353),
.B(n_352),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_965),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1031),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_980),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1086),
.B(n_758),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1016),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_980),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1044),
.A2(n_695),
.B(n_688),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1136),
.A2(n_779),
.B(n_778),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1013),
.A2(n_732),
.B(n_641),
.Y(n_1218)
);

AOI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1128),
.A2(n_778),
.B(n_737),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1019),
.A2(n_1041),
.B(n_1056),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1086),
.B(n_732),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1097),
.A2(n_704),
.B(n_695),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1046),
.B(n_732),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_983),
.A2(n_704),
.B(n_696),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_986),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1131),
.A2(n_428),
.B(n_396),
.C(n_356),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1131),
.A2(n_1065),
.B(n_1060),
.C(n_1098),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1036),
.B(n_694),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_983),
.A2(n_704),
.B(n_696),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1047),
.A2(n_763),
.B(n_737),
.Y(n_1230)
);

INVxp67_ASAP7_75t_L g1231 ( 
.A(n_1049),
.Y(n_1231)
);

CKINVDCx14_ASAP7_75t_R g1232 ( 
.A(n_973),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_992),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1065),
.A2(n_704),
.B1(n_750),
.B2(n_739),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1048),
.B(n_737),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1031),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_983),
.A2(n_696),
.B(n_694),
.Y(n_1237)
);

OA21x2_ASAP7_75t_L g1238 ( 
.A1(n_1118),
.A2(n_780),
.B(n_763),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1063),
.A2(n_780),
.B(n_763),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1099),
.B(n_780),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_SL g1241 ( 
.A(n_973),
.B(n_421),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1119),
.A2(n_784),
.B(n_782),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1036),
.B(n_782),
.Y(n_1243)
);

AO21x2_ASAP7_75t_L g1244 ( 
.A1(n_1080),
.A2(n_784),
.B(n_782),
.Y(n_1244)
);

BUFx12f_ASAP7_75t_L g1245 ( 
.A(n_1112),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1099),
.B(n_1103),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_975),
.A2(n_696),
.B(n_694),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1042),
.B(n_986),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1145),
.A2(n_1120),
.B(n_1129),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_SL g1250 ( 
.A1(n_1083),
.A2(n_786),
.B(n_784),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1066),
.B(n_786),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1091),
.A2(n_786),
.B(n_787),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1091),
.A2(n_787),
.B(n_488),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1067),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1018),
.B(n_360),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_981),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1042),
.B(n_787),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1031),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1091),
.A2(n_488),
.B(n_485),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_985),
.A2(n_1077),
.B1(n_1054),
.B2(n_1059),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_984),
.B(n_696),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_981),
.A2(n_492),
.B(n_491),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1103),
.B(n_739),
.Y(n_1263)
);

AOI21xp33_ASAP7_75t_L g1264 ( 
.A1(n_1149),
.A2(n_363),
.B(n_361),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1111),
.B(n_1113),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1054),
.A2(n_750),
.B1(n_739),
.B2(n_713),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1089),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1111),
.A2(n_576),
.B(n_748),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1113),
.B(n_508),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_992),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1116),
.A2(n_576),
.B(n_748),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1116),
.B(n_750),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1117),
.B(n_750),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_994),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1117),
.B(n_509),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_976),
.A2(n_731),
.B(n_713),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1043),
.A2(n_576),
.B(n_748),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_982),
.A2(n_1008),
.B(n_1003),
.Y(n_1278)
);

NAND2xp33_ASAP7_75t_L g1279 ( 
.A(n_984),
.B(n_750),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_962),
.B(n_491),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_994),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_984),
.B(n_697),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1124),
.A2(n_776),
.B(n_748),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_982),
.A2(n_492),
.B(n_530),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1003),
.B(n_509),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1008),
.A2(n_531),
.B(n_513),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_997),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1020),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1118),
.B(n_697),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_976),
.A2(n_731),
.B(n_713),
.Y(n_1290)
);

INVx5_ASAP7_75t_L g1291 ( 
.A(n_1031),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1020),
.A2(n_531),
.B(n_513),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1052),
.A2(n_1051),
.B(n_1122),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1023),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_SL g1295 ( 
.A1(n_984),
.A2(n_697),
.B(n_731),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1052),
.A2(n_731),
.B(n_713),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_967),
.A2(n_697),
.B1(n_713),
.B2(n_731),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1072),
.B(n_511),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1089),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1023),
.B(n_511),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1024),
.A2(n_1028),
.B(n_1027),
.Y(n_1301)
);

O2A1O1Ixp5_ASAP7_75t_L g1302 ( 
.A1(n_1058),
.A2(n_515),
.B(n_517),
.C(n_543),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1024),
.A2(n_533),
.B(n_517),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1027),
.A2(n_533),
.B(n_518),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1028),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_984),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1122),
.B(n_697),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_SL g1308 ( 
.A(n_1053),
.B(n_421),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1139),
.B(n_368),
.Y(n_1309)
);

AOI31xp67_ASAP7_75t_L g1310 ( 
.A1(n_1030),
.A2(n_530),
.A3(n_515),
.B(n_543),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1015),
.A2(n_129),
.B(n_112),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1067),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1072),
.B(n_518),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1139),
.B(n_371),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1140),
.A2(n_1143),
.B(n_1142),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_997),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1030),
.A2(n_534),
.B(n_521),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1057),
.A2(n_534),
.B(n_521),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1162),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1192),
.A2(n_1061),
.B(n_1130),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1212),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_SL g1322 ( 
.A1(n_1293),
.A2(n_1083),
.B(n_1057),
.Y(n_1322)
);

CKINVDCx11_ASAP7_75t_R g1323 ( 
.A(n_1245),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1190),
.B(n_1000),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1162),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_SL g1326 ( 
.A1(n_1315),
.A2(n_1084),
.B(n_1002),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1246),
.A2(n_1070),
.B1(n_1106),
.B2(n_1022),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1175),
.A2(n_1127),
.B(n_1002),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1212),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1194),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1161),
.A2(n_1096),
.B1(n_1144),
.B2(n_968),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1160),
.A2(n_1114),
.B1(n_1123),
.B2(n_966),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1154),
.A2(n_1165),
.B(n_1182),
.C(n_1227),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1175),
.A2(n_1006),
.B(n_1000),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1190),
.A2(n_1173),
.B1(n_1174),
.B2(n_1170),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1215),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1186),
.A2(n_1011),
.B(n_1006),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1215),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1230),
.A2(n_1038),
.B(n_1011),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1187),
.Y(n_1340)
);

AOI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1219),
.A2(n_1055),
.B(n_1038),
.Y(n_1341)
);

AO21x2_ASAP7_75t_L g1342 ( 
.A1(n_1152),
.A2(n_1104),
.B(n_1055),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1230),
.A2(n_1121),
.B(n_1142),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1239),
.A2(n_1143),
.B(n_1068),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1281),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1281),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1153),
.A2(n_1137),
.B(n_1135),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1239),
.A2(n_1033),
.B(n_1146),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1203),
.A2(n_1146),
.B(n_1088),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1169),
.B(n_988),
.Y(n_1350)
);

INVxp33_ASAP7_75t_SL g1351 ( 
.A(n_1167),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1203),
.A2(n_1088),
.B(n_1084),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1265),
.B(n_1035),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1287),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1214),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1225),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1248),
.A2(n_1181),
.B1(n_1183),
.B2(n_1257),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1166),
.A2(n_1209),
.B1(n_1264),
.B2(n_1114),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1298),
.B(n_1313),
.Y(n_1359)
);

CKINVDCx11_ASAP7_75t_R g1360 ( 
.A(n_1245),
.Y(n_1360)
);

BUFx10_ASAP7_75t_L g1361 ( 
.A(n_1202),
.Y(n_1361)
);

BUFx8_ASAP7_75t_L g1362 ( 
.A(n_1225),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1226),
.B(n_1010),
.C(n_1037),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1164),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_SL g1365 ( 
.A1(n_1241),
.A2(n_1078),
.B1(n_1150),
.B2(n_1112),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1188),
.A2(n_1148),
.B(n_1147),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1287),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1208),
.A2(n_1040),
.B(n_1039),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1257),
.B(n_1269),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1208),
.A2(n_1039),
.B(n_1025),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1218),
.A2(n_1253),
.B(n_1278),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1186),
.A2(n_524),
.B(n_520),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1187),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1218),
.A2(n_1039),
.B(n_1025),
.Y(n_1374)
);

AO21x2_ASAP7_75t_L g1375 ( 
.A1(n_1188),
.A2(n_1076),
.B(n_1110),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1253),
.A2(n_1045),
.B(n_1025),
.Y(n_1376)
);

O2A1O1Ixp33_ASAP7_75t_SL g1377 ( 
.A1(n_1176),
.A2(n_1045),
.B(n_1050),
.C(n_1005),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1198),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1254),
.B(n_1005),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1198),
.Y(n_1380)
);

NAND2x1p5_ASAP7_75t_L g1381 ( 
.A(n_1185),
.B(n_1106),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1171),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1278),
.A2(n_1050),
.B(n_1045),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1269),
.B(n_1035),
.Y(n_1384)
);

NAND2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1185),
.B(n_1106),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1201),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1301),
.A2(n_1050),
.B(n_1115),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1249),
.A2(n_1074),
.B(n_1058),
.Y(n_1388)
);

CKINVDCx8_ASAP7_75t_R g1389 ( 
.A(n_1291),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_1155),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1201),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1301),
.A2(n_1115),
.B(n_1005),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1252),
.A2(n_524),
.B(n_520),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1298),
.B(n_1123),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1313),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1260),
.A2(n_538),
.A3(n_536),
.B(n_535),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1252),
.A2(n_535),
.B(n_526),
.Y(n_1397)
);

AOI22x1_ASAP7_75t_L g1398 ( 
.A1(n_1158),
.A2(n_1074),
.B1(n_1015),
.B2(n_1087),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1193),
.A2(n_1292),
.B(n_1286),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1223),
.B(n_1074),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1256),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1223),
.B(n_1243),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1191),
.A2(n_1021),
.B(n_972),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1309),
.B(n_1123),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1275),
.B(n_1134),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1156),
.A2(n_536),
.B(n_526),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1195),
.A2(n_1021),
.B(n_972),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1256),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1314),
.B(n_1123),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1288),
.Y(n_1410)
);

NOR2x1_ASAP7_75t_SL g1411 ( 
.A(n_1291),
.B(n_1106),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1288),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1166),
.A2(n_966),
.B1(n_1092),
.B2(n_1106),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1166),
.A2(n_966),
.B1(n_1092),
.B2(n_1062),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1294),
.Y(n_1415)
);

AOI31xp67_ASAP7_75t_L g1416 ( 
.A1(n_1310),
.A2(n_1228),
.A3(n_1305),
.B(n_1294),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1157),
.A2(n_1070),
.B1(n_1015),
.B2(n_1059),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1243),
.B(n_972),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1197),
.A2(n_1021),
.B(n_1087),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1156),
.A2(n_538),
.B(n_998),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1305),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_SL g1422 ( 
.A1(n_1261),
.A2(n_979),
.B(n_987),
.C(n_991),
.Y(n_1422)
);

INVxp67_ASAP7_75t_SL g1423 ( 
.A(n_1279),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1231),
.B(n_1150),
.Y(n_1424)
);

OAI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1308),
.A2(n_966),
.B1(n_969),
.B2(n_1090),
.C(n_1108),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1168),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1168),
.Y(n_1427)
);

INVxp33_ASAP7_75t_SL g1428 ( 
.A(n_1255),
.Y(n_1428)
);

OAI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1199),
.A2(n_1053),
.B1(n_1108),
.B2(n_969),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1217),
.A2(n_998),
.B(n_1059),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1286),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1292),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1163),
.B(n_969),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1217),
.A2(n_998),
.B(n_1059),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1303),
.Y(n_1435)
);

BUFx8_ASAP7_75t_L g1436 ( 
.A(n_1254),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1275),
.B(n_1285),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1259),
.A2(n_998),
.B(n_1059),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1303),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1259),
.A2(n_998),
.B(n_1070),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1285),
.B(n_1100),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1304),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1219),
.A2(n_1193),
.B(n_1220),
.Y(n_1443)
);

OAI222xp33_ASAP7_75t_L g1444 ( 
.A1(n_1200),
.A2(n_969),
.B1(n_392),
.B2(n_423),
.C1(n_427),
.C2(n_391),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1171),
.A2(n_1015),
.B1(n_999),
.B2(n_971),
.Y(n_1445)
);

AO21x2_ASAP7_75t_L g1446 ( 
.A1(n_1283),
.A2(n_1087),
.B(n_1095),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1304),
.Y(n_1447)
);

AO31x2_ASAP7_75t_L g1448 ( 
.A1(n_1310),
.A2(n_1100),
.A3(n_998),
.B(n_1015),
.Y(n_1448)
);

AOI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1220),
.A2(n_1095),
.B(n_1062),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1172),
.B(n_1090),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1306),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1295),
.A2(n_1064),
.B(n_1062),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1284),
.A2(n_1067),
.B(n_1138),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1312),
.B(n_1132),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1213),
.A2(n_1095),
.B(n_1069),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1284),
.A2(n_1067),
.B(n_1138),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1291),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1235),
.B(n_1132),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1221),
.A2(n_1069),
.B(n_1064),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1317),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1300),
.B(n_1133),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1317),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_SL g1463 ( 
.A1(n_1282),
.A2(n_1263),
.B(n_1272),
.C(n_1273),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1318),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1262),
.A2(n_1133),
.B(n_971),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1318),
.Y(n_1466)
);

AO31x2_ASAP7_75t_L g1467 ( 
.A1(n_1205),
.A2(n_13),
.A3(n_16),
.B(n_20),
.Y(n_1467)
);

AOI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1178),
.A2(n_406),
.B1(n_382),
.B2(n_389),
.C(n_390),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1280),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1312),
.B(n_962),
.Y(n_1470)
);

INVx5_ASAP7_75t_SL g1471 ( 
.A(n_1211),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1300),
.B(n_999),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1180),
.A2(n_1064),
.B(n_1069),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1210),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1233),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1235),
.B(n_421),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1262),
.A2(n_776),
.B(n_748),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1185),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1171),
.A2(n_412),
.B1(n_393),
.B2(n_394),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1270),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1274),
.Y(n_1481)
);

OA21x2_ASAP7_75t_L g1482 ( 
.A1(n_1206),
.A2(n_418),
.B(n_395),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1316),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1306),
.B(n_115),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1276),
.A2(n_776),
.B(n_748),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1240),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1180),
.A2(n_403),
.B(n_426),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1291),
.A2(n_425),
.B1(n_422),
.B2(n_402),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_SL g1489 ( 
.A1(n_1158),
.A2(n_213),
.B(n_204),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1280),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1267),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1290),
.A2(n_1179),
.B(n_1177),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1179),
.A2(n_776),
.B(n_199),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1178),
.A2(n_398),
.B1(n_378),
.B2(n_996),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1250),
.Y(n_1495)
);

INVx4_ASAP7_75t_SL g1496 ( 
.A(n_1211),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_SL g1497 ( 
.A(n_1333),
.B(n_1204),
.C(n_1302),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1359),
.B(n_1251),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1359),
.B(n_1251),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1362),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1428),
.A2(n_1280),
.B1(n_1204),
.B2(n_1155),
.Y(n_1501)
);

AOI221xp5_ASAP7_75t_L g1502 ( 
.A1(n_1444),
.A2(n_1311),
.B1(n_1232),
.B2(n_1268),
.C(n_1271),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1395),
.B(n_1306),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1384),
.B(n_1289),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1428),
.A2(n_1155),
.B1(n_1244),
.B2(n_1232),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1451),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1323),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1350),
.B(n_1307),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1382),
.B(n_1211),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1357),
.A2(n_1291),
.B1(n_1299),
.B2(n_1267),
.Y(n_1510)
);

A2O1A1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1320),
.A2(n_1279),
.B(n_1196),
.C(n_1299),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1382),
.B(n_1211),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_R g1513 ( 
.A(n_1360),
.B(n_1390),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1476),
.B(n_1159),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1389),
.Y(n_1515)
);

AOI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1468),
.A2(n_1311),
.B1(n_1250),
.B2(n_1242),
.C(n_1277),
.Y(n_1516)
);

NAND3xp33_ASAP7_75t_SL g1517 ( 
.A(n_1358),
.B(n_1297),
.C(n_1184),
.Y(n_1517)
);

NAND2xp33_ASAP7_75t_R g1518 ( 
.A(n_1482),
.B(n_1267),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1474),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1423),
.A2(n_1295),
.B(n_1299),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1319),
.Y(n_1521)
);

INVxp33_ASAP7_75t_L g1522 ( 
.A(n_1330),
.Y(n_1522)
);

NOR2x1p5_ASAP7_75t_L g1523 ( 
.A(n_1405),
.B(n_1236),
.Y(n_1523)
);

OAI211xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1331),
.A2(n_1247),
.B(n_1296),
.C(n_1207),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1361),
.A2(n_1258),
.B1(n_1236),
.B2(n_1184),
.Y(n_1525)
);

NAND2xp33_ASAP7_75t_R g1526 ( 
.A(n_1482),
.B(n_1238),
.Y(n_1526)
);

AND2x2_ASAP7_75t_SL g1527 ( 
.A(n_1413),
.B(n_1236),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1361),
.A2(n_1258),
.B1(n_1236),
.B2(n_1184),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1363),
.A2(n_1244),
.B1(n_1196),
.B2(n_1238),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1452),
.A2(n_1388),
.B(n_1398),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1389),
.Y(n_1531)
);

OR2x6_ASAP7_75t_L g1532 ( 
.A(n_1381),
.B(n_1177),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1451),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_1362),
.Y(n_1534)
);

OAI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1437),
.A2(n_1258),
.B1(n_1236),
.B2(n_1238),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1476),
.B(n_1159),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1457),
.B(n_1258),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1335),
.A2(n_1216),
.B(n_1222),
.Y(n_1538)
);

NAND2xp33_ASAP7_75t_SL g1539 ( 
.A(n_1353),
.B(n_1258),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1361),
.A2(n_1244),
.B1(n_1234),
.B2(n_1266),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1335),
.A2(n_1189),
.B1(n_16),
.B2(n_20),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1324),
.A2(n_1189),
.B1(n_21),
.B2(n_22),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1474),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1470),
.B(n_1159),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1362),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1357),
.A2(n_1189),
.B1(n_21),
.B2(n_23),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1324),
.A2(n_1369),
.B1(n_1394),
.B2(n_1347),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_1356),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1331),
.A2(n_1237),
.B1(n_1229),
.B2(n_1224),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1332),
.A2(n_1409),
.B1(n_1404),
.B2(n_1425),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1475),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1356),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1364),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1404),
.A2(n_1409),
.B1(n_1394),
.B2(n_1414),
.Y(n_1554)
);

AOI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1494),
.A2(n_13),
.B1(n_23),
.B2(n_24),
.C(n_26),
.Y(n_1555)
);

OAI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1441),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1418),
.B(n_1159),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1355),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1457),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1398),
.A2(n_1159),
.B1(n_34),
.B2(n_37),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1325),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1402),
.B(n_30),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1436),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1402),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1433),
.A2(n_776),
.B1(n_44),
.B2(n_45),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1418),
.B(n_43),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1446),
.A2(n_776),
.B(n_193),
.Y(n_1567)
);

INVx4_ASAP7_75t_L g1568 ( 
.A(n_1457),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1475),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1400),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_1570)
);

OR2x6_ASAP7_75t_L g1571 ( 
.A(n_1381),
.B(n_190),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1458),
.B(n_46),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1446),
.A2(n_189),
.B(n_186),
.Y(n_1573)
);

A2O1A1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1419),
.A2(n_49),
.B(n_51),
.C(n_53),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1454),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1446),
.A2(n_183),
.B(n_182),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_SL g1577 ( 
.A1(n_1351),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_1577)
);

NOR2xp67_ASAP7_75t_L g1578 ( 
.A(n_1355),
.B(n_178),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1400),
.B(n_56),
.Y(n_1579)
);

CKINVDCx16_ASAP7_75t_R g1580 ( 
.A(n_1424),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1450),
.A2(n_1351),
.B1(n_1490),
.B2(n_1429),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1469),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_1582)
);

INVx6_ASAP7_75t_L g1583 ( 
.A(n_1436),
.Y(n_1583)
);

OA21x2_ASAP7_75t_L g1584 ( 
.A1(n_1443),
.A2(n_65),
.B(n_67),
.Y(n_1584)
);

OAI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1371),
.A2(n_174),
.B(n_173),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1365),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1458),
.B(n_1486),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1489),
.A2(n_69),
.B1(n_73),
.B2(n_74),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1327),
.B(n_73),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1371),
.A2(n_169),
.B(n_167),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1334),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1492),
.A2(n_163),
.B(n_158),
.Y(n_1592)
);

NAND2x1_ASAP7_75t_L g1593 ( 
.A(n_1326),
.B(n_153),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1489),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_1594)
);

BUFx4f_ASAP7_75t_L g1595 ( 
.A(n_1457),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1483),
.B(n_75),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1436),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1470),
.B(n_150),
.Y(n_1598)
);

AOI21xp33_ASAP7_75t_L g1599 ( 
.A1(n_1461),
.A2(n_77),
.B(n_78),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1480),
.Y(n_1600)
);

INVx4_ASAP7_75t_SL g1601 ( 
.A(n_1457),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1463),
.A2(n_141),
.B(n_140),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1433),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_1603)
);

INVxp33_ASAP7_75t_L g1604 ( 
.A(n_1472),
.Y(n_1604)
);

INVx4_ASAP7_75t_L g1605 ( 
.A(n_1496),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1483),
.B(n_84),
.Y(n_1606)
);

AOI222xp33_ASAP7_75t_L g1607 ( 
.A1(n_1479),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.C1(n_90),
.C2(n_91),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1486),
.A2(n_85),
.B1(n_89),
.B2(n_90),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_SL g1609 ( 
.A1(n_1366),
.A2(n_91),
.B1(n_94),
.B2(n_100),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1480),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1482),
.A2(n_100),
.B1(n_102),
.B2(n_117),
.Y(n_1611)
);

OAI21x1_ASAP7_75t_L g1612 ( 
.A1(n_1492),
.A2(n_119),
.B(n_121),
.Y(n_1612)
);

OAI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1403),
.A2(n_102),
.B1(n_125),
.B2(n_1407),
.C(n_1422),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1390),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1366),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1481),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1482),
.A2(n_1366),
.B1(n_1481),
.B2(n_1375),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_1470),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1342),
.A2(n_1417),
.B(n_1459),
.Y(n_1619)
);

INVx4_ASAP7_75t_L g1620 ( 
.A(n_1496),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1342),
.A2(n_1455),
.B(n_1411),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1420),
.A2(n_1449),
.B(n_1443),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1321),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1454),
.B(n_1321),
.Y(n_1624)
);

INVx4_ASAP7_75t_L g1625 ( 
.A(n_1496),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1375),
.A2(n_1367),
.B1(n_1354),
.B2(n_1338),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1329),
.Y(n_1627)
);

CKINVDCx11_ASAP7_75t_R g1628 ( 
.A(n_1470),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1375),
.A2(n_1484),
.B1(n_1445),
.B2(n_1411),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1334),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1454),
.B(n_1329),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1336),
.Y(n_1632)
);

NAND2xp33_ASAP7_75t_SL g1633 ( 
.A(n_1454),
.B(n_1484),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1336),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1379),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1338),
.A2(n_1345),
.B1(n_1367),
.B2(n_1354),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1379),
.B(n_1484),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1473),
.A2(n_1344),
.B(n_1377),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1345),
.B(n_1346),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1344),
.A2(n_1343),
.B(n_1328),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1346),
.A2(n_1326),
.B1(n_1380),
.B2(n_1378),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1381),
.A2(n_1385),
.B1(n_1471),
.B2(n_1488),
.Y(n_1642)
);

CKINVDCx11_ASAP7_75t_R g1643 ( 
.A(n_1496),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1396),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1342),
.A2(n_1430),
.B(n_1434),
.Y(n_1645)
);

AOI21xp33_ASAP7_75t_L g1646 ( 
.A1(n_1322),
.A2(n_1495),
.B(n_1487),
.Y(n_1646)
);

AND2x6_ASAP7_75t_L g1647 ( 
.A(n_1471),
.B(n_1478),
.Y(n_1647)
);

A2O1A1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1484),
.A2(n_1343),
.B(n_1440),
.C(n_1495),
.Y(n_1648)
);

AOI222xp33_ASAP7_75t_L g1649 ( 
.A1(n_1408),
.A2(n_1415),
.B1(n_1421),
.B2(n_1386),
.C1(n_1401),
.C2(n_1391),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1408),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1325),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1379),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1415),
.Y(n_1653)
);

AOI322xp5_ASAP7_75t_L g1654 ( 
.A1(n_1421),
.A2(n_1412),
.A3(n_1386),
.B1(n_1391),
.B2(n_1373),
.C1(n_1340),
.C2(n_1410),
.Y(n_1654)
);

AND2x6_ASAP7_75t_L g1655 ( 
.A(n_1471),
.B(n_1491),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1373),
.B(n_1412),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1401),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1410),
.A2(n_1322),
.B1(n_1487),
.B2(n_1372),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1393),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1385),
.Y(n_1660)
);

OR2x6_ASAP7_75t_L g1661 ( 
.A(n_1385),
.B(n_1438),
.Y(n_1661)
);

BUFx12f_ASAP7_75t_L g1662 ( 
.A(n_1471),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1487),
.A2(n_1372),
.B1(n_1337),
.B2(n_1432),
.Y(n_1663)
);

INVx4_ASAP7_75t_L g1664 ( 
.A(n_1478),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1487),
.A2(n_1372),
.B1(n_1337),
.B2(n_1462),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1372),
.A2(n_1337),
.B1(n_1432),
.B2(n_1462),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1439),
.A2(n_1460),
.B1(n_1435),
.B2(n_1442),
.C(n_1447),
.Y(n_1667)
);

OR2x6_ASAP7_75t_SL g1668 ( 
.A(n_1431),
.B(n_1447),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1491),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1416),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1467),
.B(n_1396),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1491),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1467),
.B(n_1396),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1467),
.B(n_1396),
.Y(n_1674)
);

CKINVDCx11_ASAP7_75t_R g1675 ( 
.A(n_1431),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1467),
.B(n_1396),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1393),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1337),
.A2(n_1460),
.B1(n_1439),
.B2(n_1466),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1607),
.A2(n_1466),
.B1(n_1464),
.B2(n_1339),
.Y(n_1679)
);

AOI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1556),
.A2(n_1426),
.B1(n_1427),
.B2(n_1467),
.C(n_1416),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1541),
.A2(n_1341),
.B1(n_1399),
.B2(n_1440),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1541),
.A2(n_1341),
.B1(n_1399),
.B2(n_1434),
.Y(n_1682)
);

OAI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1586),
.A2(n_1399),
.B1(n_1493),
.B2(n_1465),
.C(n_1406),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1604),
.B(n_1397),
.Y(n_1684)
);

OAI222xp33_ASAP7_75t_L g1685 ( 
.A1(n_1586),
.A2(n_1448),
.B1(n_1397),
.B2(n_1493),
.C1(n_1339),
.C2(n_1383),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1566),
.B(n_1448),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1555),
.A2(n_1348),
.B1(n_1328),
.B2(n_1352),
.Y(n_1687)
);

BUFx12f_ASAP7_75t_L g1688 ( 
.A(n_1507),
.Y(n_1688)
);

OAI21xp33_ASAP7_75t_L g1689 ( 
.A1(n_1574),
.A2(n_1352),
.B(n_1348),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1577),
.A2(n_1349),
.B1(n_1368),
.B2(n_1370),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1579),
.B(n_1448),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1587),
.B(n_1448),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1509),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1580),
.A2(n_1430),
.B1(n_1438),
.B2(n_1465),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1570),
.A2(n_1349),
.B1(n_1368),
.B2(n_1370),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1572),
.B(n_1448),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1643),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1570),
.A2(n_1374),
.B1(n_1383),
.B2(n_1387),
.Y(n_1698)
);

BUFx6f_ASAP7_75t_L g1699 ( 
.A(n_1628),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1546),
.A2(n_1374),
.B1(n_1387),
.B2(n_1392),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1506),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1544),
.B(n_1575),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1556),
.A2(n_1392),
.B1(n_1453),
.B2(n_1456),
.C(n_1376),
.Y(n_1703)
);

OAI221xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1582),
.A2(n_1453),
.B1(n_1456),
.B2(n_1376),
.C(n_1477),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1506),
.Y(n_1705)
);

NAND3xp33_ASAP7_75t_L g1706 ( 
.A(n_1574),
.B(n_1477),
.C(n_1485),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1623),
.Y(n_1707)
);

AO21x2_ASAP7_75t_L g1708 ( 
.A1(n_1646),
.A2(n_1485),
.B(n_1538),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1572),
.B(n_1637),
.Y(n_1709)
);

CKINVDCx6p67_ASAP7_75t_R g1710 ( 
.A(n_1614),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1501),
.A2(n_1505),
.B1(n_1523),
.B2(n_1547),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1543),
.Y(n_1712)
);

AOI322xp5_ASAP7_75t_L g1713 ( 
.A1(n_1564),
.A2(n_1582),
.A3(n_1546),
.B1(n_1542),
.B2(n_1609),
.C1(n_1611),
.C2(n_1599),
.Y(n_1713)
);

BUFx12f_ASAP7_75t_L g1714 ( 
.A(n_1597),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1550),
.A2(n_1497),
.B1(n_1554),
.B2(n_1501),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1564),
.A2(n_1542),
.B1(n_1589),
.B2(n_1603),
.Y(n_1716)
);

OAI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1589),
.A2(n_1530),
.B(n_1602),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1611),
.A2(n_1608),
.B1(n_1588),
.B2(n_1594),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1596),
.B(n_1606),
.Y(n_1719)
);

INVx4_ASAP7_75t_SL g1720 ( 
.A(n_1583),
.Y(n_1720)
);

A2O1A1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1502),
.A2(n_1633),
.B(n_1619),
.C(n_1576),
.Y(n_1721)
);

A2O1A1Ixp33_ASAP7_75t_L g1722 ( 
.A1(n_1573),
.A2(n_1516),
.B(n_1539),
.C(n_1567),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1551),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1560),
.A2(n_1565),
.B1(n_1562),
.B2(n_1536),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1498),
.B(n_1499),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1544),
.B(n_1575),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1514),
.A2(n_1547),
.B1(n_1615),
.B2(n_1522),
.Y(n_1727)
);

AOI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1522),
.A2(n_1553),
.B1(n_1626),
.B2(n_1548),
.C(n_1617),
.Y(n_1728)
);

OAI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1549),
.A2(n_1524),
.B(n_1508),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1557),
.B(n_1635),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1552),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1527),
.A2(n_1583),
.B1(n_1563),
.B2(n_1531),
.Y(n_1732)
);

AOI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1626),
.A2(n_1617),
.B1(n_1676),
.B2(n_1674),
.C(n_1558),
.Y(n_1733)
);

OR2x6_ASAP7_75t_L g1734 ( 
.A(n_1621),
.B(n_1532),
.Y(n_1734)
);

AOI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1517),
.A2(n_1505),
.B1(n_1503),
.B2(n_1510),
.C(n_1535),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1624),
.B(n_1631),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1504),
.A2(n_1527),
.B1(n_1629),
.B2(n_1583),
.Y(n_1737)
);

OAI221xp5_ASAP7_75t_SL g1738 ( 
.A1(n_1571),
.A2(n_1540),
.B1(n_1673),
.B2(n_1671),
.C(n_1545),
.Y(n_1738)
);

OAI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1578),
.A2(n_1540),
.B1(n_1593),
.B2(n_1571),
.C(n_1500),
.Y(n_1739)
);

A2O1A1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1520),
.A2(n_1598),
.B(n_1511),
.C(n_1531),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1675),
.A2(n_1571),
.B1(n_1500),
.B2(n_1563),
.Y(n_1741)
);

AOI33xp33_ASAP7_75t_L g1742 ( 
.A1(n_1636),
.A2(n_1569),
.A3(n_1600),
.B1(n_1610),
.B2(n_1616),
.B3(n_1641),
.Y(n_1742)
);

OAI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1534),
.A2(n_1515),
.B1(n_1618),
.B2(n_1652),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1627),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1660),
.B(n_1652),
.Y(n_1745)
);

CKINVDCx14_ASAP7_75t_R g1746 ( 
.A(n_1513),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1632),
.Y(n_1747)
);

A2O1A1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1511),
.A2(n_1515),
.B(n_1595),
.C(n_1638),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1525),
.A2(n_1528),
.B1(n_1636),
.B2(n_1595),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1584),
.A2(n_1650),
.B1(n_1653),
.B2(n_1533),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1641),
.A2(n_1668),
.B1(n_1620),
.B2(n_1625),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1535),
.A2(n_1645),
.B(n_1532),
.Y(n_1752)
);

INVx5_ASAP7_75t_L g1753 ( 
.A(n_1647),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1662),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1509),
.Y(n_1755)
);

OAI211xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1649),
.A2(n_1654),
.B(n_1648),
.C(n_1529),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1529),
.A2(n_1648),
.B(n_1642),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1584),
.A2(n_1634),
.B1(n_1644),
.B2(n_1657),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1532),
.A2(n_1640),
.B(n_1661),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1584),
.A2(n_1644),
.B1(n_1651),
.B2(n_1521),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1512),
.B(n_1672),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1639),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1561),
.A2(n_1512),
.B1(n_1660),
.B2(n_1656),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1591),
.Y(n_1764)
);

OR2x6_ASAP7_75t_L g1765 ( 
.A(n_1661),
.B(n_1625),
.Y(n_1765)
);

OAI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1518),
.A2(n_1605),
.B1(n_1620),
.B2(n_1664),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1667),
.Y(n_1767)
);

OAI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1518),
.A2(n_1605),
.B1(n_1664),
.B2(n_1568),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1647),
.A2(n_1655),
.B1(n_1669),
.B2(n_1658),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1669),
.B(n_1559),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1559),
.B(n_1568),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_1647),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_1601),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1601),
.B(n_1537),
.Y(n_1774)
);

OAI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1658),
.A2(n_1665),
.B1(n_1663),
.B2(n_1526),
.C(n_1677),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1647),
.B(n_1655),
.Y(n_1776)
);

BUFx4f_ASAP7_75t_SL g1777 ( 
.A(n_1647),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_SL g1778 ( 
.A1(n_1655),
.A2(n_1585),
.B1(n_1590),
.B2(n_1612),
.Y(n_1778)
);

AOI221xp5_ASAP7_75t_L g1779 ( 
.A1(n_1663),
.A2(n_1665),
.B1(n_1678),
.B2(n_1666),
.C(n_1659),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_SL g1780 ( 
.A1(n_1655),
.A2(n_1592),
.B1(n_1537),
.B2(n_1661),
.Y(n_1780)
);

A2O1A1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1622),
.A2(n_1630),
.B(n_1678),
.C(n_1666),
.Y(n_1781)
);

OAI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1526),
.A2(n_1670),
.B1(n_1601),
.B2(n_1655),
.Y(n_1782)
);

AOI221xp5_ASAP7_75t_L g1783 ( 
.A1(n_1670),
.A2(n_1161),
.B1(n_1073),
.B2(n_1079),
.C(n_1160),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1607),
.A2(n_1161),
.B1(n_1141),
.B2(n_1073),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1607),
.A2(n_1161),
.B1(n_1141),
.B2(n_1073),
.Y(n_1785)
);

OAI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1586),
.A2(n_1161),
.B1(n_790),
.B2(n_1079),
.C(n_1073),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1566),
.B(n_1579),
.Y(n_1787)
);

OAI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1586),
.A2(n_1161),
.B1(n_790),
.B2(n_1079),
.C(n_1073),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1581),
.A2(n_1034),
.B1(n_1428),
.B2(n_790),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1566),
.B(n_1579),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1607),
.A2(n_1161),
.B1(n_1141),
.B2(n_1073),
.Y(n_1791)
);

BUFx4f_ASAP7_75t_SL g1792 ( 
.A(n_1534),
.Y(n_1792)
);

OAI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1586),
.A2(n_1161),
.B1(n_790),
.B2(n_1079),
.C(n_1073),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_L g1794 ( 
.A(n_1643),
.Y(n_1794)
);

AOI21xp33_ASAP7_75t_L g1795 ( 
.A1(n_1613),
.A2(n_1073),
.B(n_1102),
.Y(n_1795)
);

OAI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1613),
.A2(n_1126),
.B1(n_809),
.B2(n_906),
.Y(n_1796)
);

AOI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1550),
.A2(n_1161),
.B1(n_1428),
.B2(n_1034),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1557),
.B(n_1498),
.Y(n_1798)
);

OA21x2_ASAP7_75t_L g1799 ( 
.A1(n_1640),
.A2(n_1443),
.B(n_1646),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1607),
.A2(n_1161),
.B1(n_1141),
.B2(n_1073),
.Y(n_1800)
);

AO221x2_ASAP7_75t_L g1801 ( 
.A1(n_1546),
.A2(n_1160),
.B1(n_1556),
.B2(n_1444),
.C(n_843),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1607),
.A2(n_1161),
.B1(n_1141),
.B2(n_1073),
.Y(n_1802)
);

OAI221xp5_ASAP7_75t_L g1803 ( 
.A1(n_1586),
.A2(n_1161),
.B1(n_790),
.B2(n_1079),
.C(n_1073),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1607),
.A2(n_1161),
.B1(n_1141),
.B2(n_1073),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1581),
.A2(n_1034),
.B1(n_1428),
.B2(n_790),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1555),
.B(n_790),
.C(n_1079),
.Y(n_1806)
);

OAI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1586),
.A2(n_1161),
.B1(n_790),
.B2(n_1079),
.C(n_1073),
.Y(n_1807)
);

AOI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1550),
.A2(n_1161),
.B1(n_1428),
.B2(n_1034),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1546),
.B(n_1333),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1519),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1607),
.A2(n_1161),
.B1(n_1141),
.B2(n_1073),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1581),
.A2(n_1034),
.B1(n_1428),
.B2(n_790),
.Y(n_1812)
);

OAI21xp5_ASAP7_75t_SL g1813 ( 
.A1(n_1586),
.A2(n_1161),
.B(n_790),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1607),
.A2(n_1161),
.B1(n_1141),
.B2(n_1073),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_1507),
.Y(n_1815)
);

AO21x2_ASAP7_75t_L g1816 ( 
.A1(n_1646),
.A2(n_1538),
.B(n_1530),
.Y(n_1816)
);

AOI21xp33_ASAP7_75t_L g1817 ( 
.A1(n_1613),
.A2(n_1073),
.B(n_1102),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1607),
.A2(n_1161),
.B1(n_1141),
.B2(n_1073),
.Y(n_1818)
);

A2O1A1Ixp33_ASAP7_75t_L g1819 ( 
.A1(n_1613),
.A2(n_1161),
.B(n_795),
.C(n_790),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1566),
.B(n_1579),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1607),
.A2(n_1161),
.B1(n_1141),
.B2(n_1073),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1566),
.B(n_1579),
.Y(n_1822)
);

OAI211xp5_ASAP7_75t_L g1823 ( 
.A1(n_1586),
.A2(n_1161),
.B(n_1073),
.C(n_1607),
.Y(n_1823)
);

AO21x2_ASAP7_75t_L g1824 ( 
.A1(n_1646),
.A2(n_1538),
.B(n_1530),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1604),
.B(n_1161),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1566),
.B(n_1579),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1607),
.A2(n_1161),
.B1(n_1141),
.B2(n_1073),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1587),
.B(n_1498),
.Y(n_1828)
);

AO21x2_ASAP7_75t_L g1829 ( 
.A1(n_1646),
.A2(n_1538),
.B(n_1530),
.Y(n_1829)
);

AOI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1556),
.A2(n_1161),
.B1(n_1073),
.B2(n_1079),
.C(n_1160),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1506),
.Y(n_1831)
);

OAI211xp5_ASAP7_75t_L g1832 ( 
.A1(n_1586),
.A2(n_1161),
.B(n_1073),
.C(n_1607),
.Y(n_1832)
);

OAI211xp5_ASAP7_75t_SL g1833 ( 
.A1(n_1607),
.A2(n_1161),
.B(n_1331),
.C(n_646),
.Y(n_1833)
);

AOI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1556),
.A2(n_1161),
.B1(n_1073),
.B2(n_1079),
.C(n_1160),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1707),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1686),
.B(n_1691),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1707),
.Y(n_1837)
);

INVx3_ASAP7_75t_SL g1838 ( 
.A(n_1753),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1747),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1764),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1764),
.B(n_1696),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1744),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1816),
.B(n_1824),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1734),
.B(n_1816),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1824),
.B(n_1829),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1829),
.B(n_1779),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1712),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1723),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1734),
.B(n_1692),
.Y(n_1849)
);

BUFx2_ASAP7_75t_L g1850 ( 
.A(n_1757),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1781),
.B(n_1760),
.Y(n_1851)
);

BUFx2_ASAP7_75t_L g1852 ( 
.A(n_1701),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1799),
.B(n_1758),
.Y(n_1853)
);

BUFx3_ASAP7_75t_L g1854 ( 
.A(n_1765),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1705),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1799),
.B(n_1758),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1810),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1762),
.B(n_1767),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1831),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1801),
.A2(n_1807),
.B1(n_1786),
.B2(n_1788),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1799),
.B(n_1759),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1752),
.B(n_1708),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1750),
.Y(n_1863)
);

BUFx3_ASAP7_75t_L g1864 ( 
.A(n_1765),
.Y(n_1864)
);

INVxp67_ASAP7_75t_SL g1865 ( 
.A(n_1750),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1801),
.A2(n_1793),
.B1(n_1803),
.B2(n_1833),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1708),
.B(n_1729),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1775),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1702),
.B(n_1726),
.Y(n_1869)
);

INVxp67_ASAP7_75t_L g1870 ( 
.A(n_1684),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1798),
.B(n_1736),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1694),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1680),
.B(n_1733),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1716),
.A2(n_1804),
.B1(n_1802),
.B2(n_1784),
.Y(n_1874)
);

HB1xp67_ASAP7_75t_L g1875 ( 
.A(n_1681),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1740),
.B(n_1721),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1684),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1682),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1700),
.B(n_1769),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1731),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1700),
.B(n_1769),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1683),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1695),
.B(n_1727),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1706),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1695),
.B(n_1698),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1698),
.B(n_1687),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1761),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1703),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1828),
.B(n_1725),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1742),
.Y(n_1890)
);

BUFx3_ASAP7_75t_L g1891 ( 
.A(n_1776),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1770),
.Y(n_1892)
);

NOR2x1_ASAP7_75t_L g1893 ( 
.A(n_1717),
.B(n_1748),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1738),
.B(n_1689),
.Y(n_1894)
);

AOI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1795),
.A2(n_1817),
.B1(n_1813),
.B2(n_1834),
.C(n_1830),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1687),
.B(n_1690),
.Y(n_1896)
);

AOI221x1_ASAP7_75t_L g1897 ( 
.A1(n_1819),
.A2(n_1806),
.B1(n_1722),
.B2(n_1756),
.C(n_1812),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1690),
.B(n_1809),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1782),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1728),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1768),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1809),
.B(n_1709),
.Y(n_1902)
);

BUFx2_ASAP7_75t_L g1903 ( 
.A(n_1766),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1730),
.B(n_1719),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1735),
.B(n_1732),
.Y(n_1905)
);

INVx2_ASAP7_75t_R g1906 ( 
.A(n_1704),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1745),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1737),
.B(n_1763),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1751),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1780),
.Y(n_1910)
);

INVx5_ASAP7_75t_L g1911 ( 
.A(n_1693),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1787),
.B(n_1826),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1790),
.B(n_1820),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1825),
.B(n_1715),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1822),
.B(n_1825),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1693),
.B(n_1801),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1749),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1836),
.B(n_1711),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1835),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1870),
.B(n_1808),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1836),
.B(n_1755),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1870),
.B(n_1797),
.Y(n_1922)
);

BUFx4f_ASAP7_75t_L g1923 ( 
.A(n_1876),
.Y(n_1923)
);

AND2x4_ASAP7_75t_SL g1924 ( 
.A(n_1876),
.B(n_1699),
.Y(n_1924)
);

AOI211xp5_ASAP7_75t_L g1925 ( 
.A1(n_1850),
.A2(n_1796),
.B(n_1789),
.C(n_1805),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1854),
.B(n_1720),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1860),
.A2(n_1804),
.B1(n_1827),
.B2(n_1802),
.Y(n_1927)
);

OAI33xp33_ASAP7_75t_L g1928 ( 
.A1(n_1914),
.A2(n_1743),
.A3(n_1772),
.B1(n_1815),
.B2(n_1832),
.B3(n_1823),
.Y(n_1928)
);

OAI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1897),
.A2(n_1827),
.B(n_1821),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1877),
.B(n_1783),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1836),
.B(n_1841),
.Y(n_1931)
);

BUFx2_ASAP7_75t_L g1932 ( 
.A(n_1854),
.Y(n_1932)
);

BUFx2_ASAP7_75t_L g1933 ( 
.A(n_1854),
.Y(n_1933)
);

NOR2x1_ASAP7_75t_L g1934 ( 
.A(n_1893),
.B(n_1773),
.Y(n_1934)
);

BUFx2_ASAP7_75t_SL g1935 ( 
.A(n_1892),
.Y(n_1935)
);

AOI211xp5_ASAP7_75t_L g1936 ( 
.A1(n_1850),
.A2(n_1739),
.B(n_1699),
.C(n_1794),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_R g1937 ( 
.A(n_1917),
.B(n_1746),
.Y(n_1937)
);

OAI221xp5_ASAP7_75t_L g1938 ( 
.A1(n_1860),
.A2(n_1821),
.B1(n_1818),
.B2(n_1814),
.C(n_1811),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1854),
.Y(n_1939)
);

AO21x2_ASAP7_75t_L g1940 ( 
.A1(n_1843),
.A2(n_1685),
.B(n_1771),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1877),
.B(n_1679),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1880),
.Y(n_1942)
);

BUFx2_ASAP7_75t_L g1943 ( 
.A(n_1864),
.Y(n_1943)
);

INVx3_ASAP7_75t_L g1944 ( 
.A(n_1869),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1842),
.Y(n_1945)
);

INVxp67_ASAP7_75t_L g1946 ( 
.A(n_1880),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1864),
.B(n_1720),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1841),
.B(n_1741),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1839),
.Y(n_1949)
);

NAND3xp33_ASAP7_75t_L g1950 ( 
.A(n_1897),
.B(n_1818),
.C(n_1814),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1852),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1842),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1874),
.A2(n_1811),
.B1(n_1800),
.B2(n_1791),
.Y(n_1953)
);

NAND3xp33_ASAP7_75t_L g1954 ( 
.A(n_1897),
.B(n_1800),
.C(n_1791),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1847),
.Y(n_1955)
);

INVxp67_ASAP7_75t_SL g1956 ( 
.A(n_1840),
.Y(n_1956)
);

AOI221xp5_ASAP7_75t_L g1957 ( 
.A1(n_1850),
.A2(n_1785),
.B1(n_1784),
.B2(n_1718),
.C(n_1716),
.Y(n_1957)
);

BUFx3_ASAP7_75t_L g1958 ( 
.A(n_1852),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1847),
.Y(n_1959)
);

AOI221xp5_ASAP7_75t_L g1960 ( 
.A1(n_1914),
.A2(n_1785),
.B1(n_1718),
.B2(n_1724),
.C(n_1741),
.Y(n_1960)
);

AOI22xp33_ASAP7_75t_L g1961 ( 
.A1(n_1866),
.A2(n_1724),
.B1(n_1714),
.B2(n_1699),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1848),
.Y(n_1962)
);

AOI221xp5_ASAP7_75t_L g1963 ( 
.A1(n_1888),
.A2(n_1679),
.B1(n_1699),
.B2(n_1754),
.C(n_1697),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1889),
.B(n_1713),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1864),
.B(n_1754),
.Y(n_1965)
);

OAI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1866),
.A2(n_1794),
.B1(n_1697),
.B2(n_1777),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1848),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1857),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1869),
.Y(n_1969)
);

OAI31xp33_ASAP7_75t_SL g1970 ( 
.A1(n_1893),
.A2(n_1774),
.A3(n_1778),
.B(n_1794),
.Y(n_1970)
);

OAI33xp33_ASAP7_75t_L g1971 ( 
.A1(n_1890),
.A2(n_1874),
.A3(n_1858),
.B1(n_1868),
.B2(n_1917),
.B3(n_1894),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1849),
.B(n_1697),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1852),
.Y(n_1973)
);

INVx3_ASAP7_75t_L g1974 ( 
.A(n_1869),
.Y(n_1974)
);

OAI321xp33_ASAP7_75t_L g1975 ( 
.A1(n_1895),
.A2(n_1697),
.A3(n_1794),
.B1(n_1714),
.B2(n_1792),
.C(n_1710),
.Y(n_1975)
);

BUFx2_ASAP7_75t_L g1976 ( 
.A(n_1864),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1841),
.B(n_1688),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1907),
.B(n_1688),
.Y(n_1978)
);

OAI221xp5_ASAP7_75t_L g1979 ( 
.A1(n_1895),
.A2(n_1900),
.B1(n_1888),
.B2(n_1868),
.C(n_1905),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1849),
.B(n_1855),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1876),
.B(n_1900),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1857),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1837),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1849),
.B(n_1855),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1837),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1889),
.B(n_1915),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1980),
.B(n_1844),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1951),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1931),
.B(n_1944),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1955),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1931),
.B(n_1861),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1980),
.B(n_1844),
.Y(n_1992)
);

OA21x2_ASAP7_75t_L g1993 ( 
.A1(n_1955),
.A2(n_1843),
.B(n_1845),
.Y(n_1993)
);

BUFx2_ASAP7_75t_L g1994 ( 
.A(n_1944),
.Y(n_1994)
);

OAI33xp33_ASAP7_75t_L g1995 ( 
.A1(n_1964),
.A2(n_1890),
.A3(n_1858),
.B1(n_1894),
.B2(n_1859),
.B3(n_1863),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1986),
.B(n_1846),
.Y(n_1996)
);

HB1xp67_ASAP7_75t_L g1997 ( 
.A(n_1973),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1959),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1959),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1956),
.B(n_1846),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1983),
.B(n_1846),
.Y(n_2001)
);

INVx3_ASAP7_75t_L g2002 ( 
.A(n_1944),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1983),
.B(n_1867),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1962),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1969),
.B(n_1861),
.Y(n_2005)
);

INVxp67_ASAP7_75t_L g2006 ( 
.A(n_1981),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1985),
.B(n_1984),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1962),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1919),
.Y(n_2009)
);

OR2x2_ASAP7_75t_L g2010 ( 
.A(n_1984),
.B(n_1844),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1958),
.B(n_1853),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1967),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1969),
.B(n_1853),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1985),
.B(n_1867),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1967),
.B(n_1867),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1968),
.Y(n_2016)
);

BUFx3_ASAP7_75t_L g2017 ( 
.A(n_1924),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1958),
.B(n_1853),
.Y(n_2018)
);

AND2x4_ASAP7_75t_L g2019 ( 
.A(n_1974),
.B(n_1911),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1974),
.B(n_1856),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1968),
.B(n_1863),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1940),
.B(n_1856),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1940),
.B(n_1851),
.Y(n_2023)
);

INVxp67_ASAP7_75t_L g2024 ( 
.A(n_1948),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1982),
.B(n_1865),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1982),
.Y(n_2026)
);

INVx1_ASAP7_75t_SL g2027 ( 
.A(n_1935),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1945),
.B(n_1865),
.Y(n_2028)
);

OR2x2_ASAP7_75t_L g2029 ( 
.A(n_1940),
.B(n_1884),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1921),
.B(n_1851),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1949),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1952),
.B(n_1859),
.Y(n_2032)
);

BUFx2_ASAP7_75t_L g2033 ( 
.A(n_1932),
.Y(n_2033)
);

OR2x2_ASAP7_75t_L g2034 ( 
.A(n_1949),
.B(n_1884),
.Y(n_2034)
);

NAND4xp25_ASAP7_75t_SL g2035 ( 
.A(n_1979),
.B(n_1925),
.C(n_1936),
.D(n_1960),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_2031),
.Y(n_2036)
);

INVxp67_ASAP7_75t_L g2037 ( 
.A(n_2030),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2006),
.B(n_1946),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2032),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1991),
.B(n_2024),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_1987),
.B(n_1941),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_2031),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2032),
.Y(n_2043)
);

OR2x2_ASAP7_75t_L g2044 ( 
.A(n_1987),
.B(n_1941),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1990),
.Y(n_2045)
);

INVx1_ASAP7_75t_SL g2046 ( 
.A(n_2017),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1990),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1998),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1998),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_2006),
.B(n_1996),
.Y(n_2050)
);

OAI322xp33_ASAP7_75t_L g2051 ( 
.A1(n_2029),
.A2(n_1930),
.A3(n_1953),
.B1(n_1950),
.B2(n_1954),
.C1(n_1938),
.C2(n_1894),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1991),
.B(n_1932),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_1987),
.B(n_1871),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1996),
.B(n_2024),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1999),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_2031),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1999),
.Y(n_2057)
);

INVx2_ASAP7_75t_SL g2058 ( 
.A(n_2033),
.Y(n_2058)
);

OR2x2_ASAP7_75t_L g2059 ( 
.A(n_1992),
.B(n_2010),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1991),
.B(n_1933),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1989),
.B(n_1933),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_1992),
.B(n_1871),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_1992),
.B(n_1871),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2004),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2030),
.B(n_1918),
.Y(n_2065)
);

INVxp67_ASAP7_75t_L g2066 ( 
.A(n_2030),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2004),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2031),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2008),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2008),
.Y(n_2070)
);

AOI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_2035),
.A2(n_1876),
.B1(n_1873),
.B2(n_1929),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2012),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1988),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2012),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_2010),
.B(n_1884),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2031),
.Y(n_2076)
);

INVx2_ASAP7_75t_SL g2077 ( 
.A(n_2033),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1989),
.B(n_1939),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2016),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_2010),
.B(n_1972),
.Y(n_2080)
);

INVx1_ASAP7_75t_SL g2081 ( 
.A(n_2017),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2028),
.B(n_1918),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2028),
.B(n_1948),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2016),
.Y(n_2084)
);

INVxp67_ASAP7_75t_L g2085 ( 
.A(n_2001),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_2029),
.B(n_1972),
.Y(n_2086)
);

BUFx2_ASAP7_75t_L g2087 ( 
.A(n_2033),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2023),
.B(n_1887),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2026),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_L g2090 ( 
.A(n_2071),
.B(n_2035),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2082),
.B(n_2065),
.Y(n_2091)
);

NAND4xp75_ASAP7_75t_L g2092 ( 
.A(n_2058),
.B(n_1934),
.C(n_1957),
.D(n_2023),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2055),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2050),
.B(n_2023),
.Y(n_2094)
);

OR2x2_ASAP7_75t_L g2095 ( 
.A(n_2041),
.B(n_2029),
.Y(n_2095)
);

INVx2_ASAP7_75t_SL g2096 ( 
.A(n_2087),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2038),
.B(n_2000),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2083),
.B(n_2000),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2055),
.Y(n_2099)
);

OAI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_2046),
.A2(n_1923),
.B1(n_1908),
.B2(n_1876),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2040),
.B(n_2022),
.Y(n_2101)
);

OR2x2_ASAP7_75t_L g2102 ( 
.A(n_2041),
.B(n_2001),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2087),
.Y(n_2103)
);

NAND3xp33_ASAP7_75t_L g2104 ( 
.A(n_2054),
.B(n_1963),
.C(n_1970),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2039),
.B(n_2022),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_2058),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2040),
.B(n_2022),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2052),
.B(n_2005),
.Y(n_2108)
);

INVxp67_ASAP7_75t_L g2109 ( 
.A(n_2073),
.Y(n_2109)
);

BUFx2_ASAP7_75t_L g2110 ( 
.A(n_2077),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2057),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2043),
.B(n_2025),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2085),
.B(n_2025),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2057),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2088),
.B(n_1942),
.Y(n_2115)
);

NOR2xp33_ASAP7_75t_L g2116 ( 
.A(n_2051),
.B(n_1977),
.Y(n_2116)
);

AND4x1_ASAP7_75t_L g2117 ( 
.A(n_2061),
.B(n_1995),
.C(n_1961),
.D(n_1971),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2037),
.B(n_2066),
.Y(n_2118)
);

CKINVDCx5p33_ASAP7_75t_R g2119 ( 
.A(n_2081),
.Y(n_2119)
);

AND2x4_ASAP7_75t_SL g2120 ( 
.A(n_2052),
.B(n_1926),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2060),
.B(n_2005),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2044),
.B(n_1942),
.Y(n_2122)
);

A2O1A1Ixp33_ASAP7_75t_L g2123 ( 
.A1(n_2077),
.A2(n_1975),
.B(n_1923),
.C(n_1905),
.Y(n_2123)
);

AND2x4_ASAP7_75t_L g2124 ( 
.A(n_2060),
.B(n_2019),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2044),
.B(n_1915),
.Y(n_2125)
);

NAND2xp33_ASAP7_75t_R g2126 ( 
.A(n_2086),
.B(n_1937),
.Y(n_2126)
);

INVx1_ASAP7_75t_SL g2127 ( 
.A(n_2086),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2053),
.B(n_1915),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2036),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2053),
.B(n_2003),
.Y(n_2130)
);

INVx1_ASAP7_75t_SL g2131 ( 
.A(n_2080),
.Y(n_2131)
);

OR2x2_ASAP7_75t_L g2132 ( 
.A(n_2062),
.B(n_2003),
.Y(n_2132)
);

OR2x2_ASAP7_75t_L g2133 ( 
.A(n_2062),
.B(n_2014),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_2063),
.B(n_2014),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_2036),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2061),
.B(n_2005),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_2078),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2072),
.Y(n_2138)
);

AOI221xp5_ASAP7_75t_L g2139 ( 
.A1(n_2090),
.A2(n_1995),
.B1(n_1928),
.B2(n_1873),
.C(n_1905),
.Y(n_2139)
);

AOI321xp33_ASAP7_75t_L g2140 ( 
.A1(n_2116),
.A2(n_2123),
.A3(n_1927),
.B1(n_2100),
.B2(n_1873),
.C(n_2118),
.Y(n_2140)
);

AOI32xp33_ASAP7_75t_L g2141 ( 
.A1(n_2092),
.A2(n_1966),
.A3(n_1898),
.B1(n_1924),
.B2(n_2027),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2099),
.Y(n_2142)
);

AOI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_2104),
.A2(n_1906),
.B1(n_1898),
.B2(n_1883),
.Y(n_2143)
);

INVxp67_ASAP7_75t_L g2144 ( 
.A(n_2126),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_2110),
.Y(n_2145)
);

OR2x2_ASAP7_75t_L g2146 ( 
.A(n_2125),
.B(n_2063),
.Y(n_2146)
);

OAI22xp33_ASAP7_75t_L g2147 ( 
.A1(n_2119),
.A2(n_1923),
.B1(n_1903),
.B2(n_1908),
.Y(n_2147)
);

NAND3xp33_ASAP7_75t_L g2148 ( 
.A(n_2117),
.B(n_1922),
.C(n_1920),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2122),
.A2(n_1906),
.B1(n_1898),
.B2(n_1883),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2119),
.B(n_2078),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2109),
.B(n_2080),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2138),
.Y(n_2152)
);

AOI221xp5_ASAP7_75t_L g2153 ( 
.A1(n_2094),
.A2(n_1851),
.B1(n_2015),
.B2(n_1875),
.C(n_1878),
.Y(n_2153)
);

AOI21xp33_ASAP7_75t_L g2154 ( 
.A1(n_2096),
.A2(n_1910),
.B(n_2075),
.Y(n_2154)
);

NOR4xp25_ASAP7_75t_SL g2155 ( 
.A(n_2110),
.B(n_1994),
.C(n_1903),
.D(n_1976),
.Y(n_2155)
);

OAI21xp5_ASAP7_75t_SL g2156 ( 
.A1(n_2092),
.A2(n_1883),
.B(n_1910),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2097),
.B(n_2059),
.Y(n_2157)
);

AOI21xp5_ASAP7_75t_L g2158 ( 
.A1(n_2115),
.A2(n_2021),
.B(n_1978),
.Y(n_2158)
);

A2O1A1Ixp33_ASAP7_75t_L g2159 ( 
.A1(n_2137),
.A2(n_1903),
.B(n_1908),
.C(n_1896),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2120),
.B(n_1989),
.Y(n_2160)
);

OAI21xp33_ASAP7_75t_L g2161 ( 
.A1(n_2131),
.A2(n_1916),
.B(n_1896),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_SL g2162 ( 
.A(n_2137),
.B(n_2027),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2127),
.B(n_2075),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_2091),
.B(n_2015),
.Y(n_2164)
);

O2A1O1Ixp33_ASAP7_75t_L g2165 ( 
.A1(n_2096),
.A2(n_1875),
.B(n_1878),
.C(n_1882),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2128),
.B(n_1912),
.Y(n_2166)
);

OAI32xp33_ASAP7_75t_L g2167 ( 
.A1(n_2103),
.A2(n_2059),
.A3(n_2011),
.B1(n_2018),
.B2(n_1997),
.Y(n_2167)
);

NAND2xp33_ASAP7_75t_SL g2168 ( 
.A(n_2101),
.B(n_1977),
.Y(n_2168)
);

AOI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_2120),
.A2(n_1896),
.B1(n_1909),
.B2(n_1862),
.Y(n_2169)
);

NOR2xp33_ASAP7_75t_L g2170 ( 
.A(n_2098),
.B(n_2113),
.Y(n_2170)
);

AOI221xp5_ASAP7_75t_L g2171 ( 
.A1(n_2103),
.A2(n_2021),
.B1(n_1862),
.B2(n_1882),
.C(n_2079),
.Y(n_2171)
);

INVx1_ASAP7_75t_SL g2172 ( 
.A(n_2095),
.Y(n_2172)
);

OAI32xp33_ASAP7_75t_L g2173 ( 
.A1(n_2106),
.A2(n_2018),
.A3(n_2011),
.B1(n_1988),
.B2(n_1997),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2099),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2124),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2112),
.B(n_1912),
.Y(n_2176)
);

O2A1O1Ixp33_ASAP7_75t_L g2177 ( 
.A1(n_2106),
.A2(n_1882),
.B(n_1862),
.C(n_1872),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_2151),
.B(n_2102),
.Y(n_2178)
);

OAI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_2143),
.A2(n_2124),
.B1(n_2017),
.B2(n_2101),
.Y(n_2179)
);

NAND4xp25_ASAP7_75t_L g2180 ( 
.A(n_2140),
.B(n_2107),
.C(n_2095),
.D(n_2105),
.Y(n_2180)
);

AOI322xp5_ASAP7_75t_L g2181 ( 
.A1(n_2143),
.A2(n_2107),
.A3(n_2136),
.B1(n_2108),
.B2(n_2121),
.C1(n_2124),
.C2(n_2130),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2144),
.B(n_2136),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2142),
.Y(n_2183)
);

OAI21xp33_ASAP7_75t_L g2184 ( 
.A1(n_2156),
.A2(n_2102),
.B(n_2093),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2152),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2174),
.Y(n_2186)
);

OAI21xp33_ASAP7_75t_L g2187 ( 
.A1(n_2141),
.A2(n_2114),
.B(n_2138),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2148),
.B(n_2108),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2145),
.Y(n_2189)
);

OAI21xp5_ASAP7_75t_SL g2190 ( 
.A1(n_2139),
.A2(n_1881),
.B(n_1879),
.Y(n_2190)
);

OAI31xp33_ASAP7_75t_L g2191 ( 
.A1(n_2159),
.A2(n_1965),
.A3(n_1978),
.B(n_2121),
.Y(n_2191)
);

AOI221x1_ASAP7_75t_L g2192 ( 
.A1(n_2159),
.A2(n_2111),
.B1(n_2135),
.B2(n_2072),
.C(n_2089),
.Y(n_2192)
);

OAI21xp33_ASAP7_75t_L g2193 ( 
.A1(n_2170),
.A2(n_2149),
.B(n_2150),
.Y(n_2193)
);

AOI322xp5_ASAP7_75t_L g2194 ( 
.A1(n_2147),
.A2(n_1902),
.A3(n_1886),
.B1(n_2111),
.B2(n_1879),
.C1(n_1881),
.C2(n_1913),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_2162),
.B(n_2170),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2163),
.Y(n_2196)
);

INVx2_ASAP7_75t_SL g2197 ( 
.A(n_2175),
.Y(n_2197)
);

INVx2_ASAP7_75t_SL g2198 ( 
.A(n_2162),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2153),
.B(n_2132),
.Y(n_2199)
);

INVx1_ASAP7_75t_SL g2200 ( 
.A(n_2172),
.Y(n_2200)
);

INVxp33_ASAP7_75t_L g2201 ( 
.A(n_2165),
.Y(n_2201)
);

HB1xp67_ASAP7_75t_L g2202 ( 
.A(n_2157),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2176),
.B(n_2132),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2160),
.Y(n_2204)
);

AOI221xp5_ASAP7_75t_L g2205 ( 
.A1(n_2167),
.A2(n_2129),
.B1(n_2135),
.B2(n_1882),
.C(n_1885),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2147),
.B(n_2133),
.Y(n_2206)
);

INVxp67_ASAP7_75t_L g2207 ( 
.A(n_2195),
.Y(n_2207)
);

OR2x2_ASAP7_75t_L g2208 ( 
.A(n_2188),
.B(n_2146),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_2195),
.B(n_2149),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2182),
.B(n_2169),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2182),
.B(n_2155),
.Y(n_2211)
);

OAI21xp33_ASAP7_75t_SL g2212 ( 
.A1(n_2198),
.A2(n_2154),
.B(n_2171),
.Y(n_2212)
);

OR2x2_ASAP7_75t_L g2213 ( 
.A(n_2200),
.B(n_2164),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_2193),
.B(n_2168),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2198),
.B(n_2158),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2202),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2202),
.B(n_2161),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2204),
.B(n_2166),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2183),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2185),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2204),
.B(n_2173),
.Y(n_2221)
);

INVx2_ASAP7_75t_SL g2222 ( 
.A(n_2197),
.Y(n_2222)
);

NAND3xp33_ASAP7_75t_L g2223 ( 
.A(n_2192),
.B(n_2177),
.C(n_2129),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_SL g2224 ( 
.A(n_2191),
.B(n_1965),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2189),
.B(n_2133),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2186),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2197),
.Y(n_2227)
);

HB1xp67_ASAP7_75t_L g2228 ( 
.A(n_2178),
.Y(n_2228)
);

NOR2x1_ASAP7_75t_L g2229 ( 
.A(n_2190),
.B(n_2135),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2196),
.Y(n_2230)
);

NAND3xp33_ASAP7_75t_L g2231 ( 
.A(n_2209),
.B(n_2201),
.C(n_2187),
.Y(n_2231)
);

AOI21xp5_ASAP7_75t_L g2232 ( 
.A1(n_2207),
.A2(n_2201),
.B(n_2199),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_L g2233 ( 
.A(n_2228),
.B(n_2184),
.Y(n_2233)
);

AOI21xp5_ASAP7_75t_L g2234 ( 
.A1(n_2212),
.A2(n_2206),
.B(n_2179),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2216),
.Y(n_2235)
);

NOR3xp33_ASAP7_75t_L g2236 ( 
.A(n_2214),
.B(n_2216),
.C(n_2230),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2215),
.B(n_2181),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2222),
.Y(n_2238)
);

NAND3xp33_ASAP7_75t_SL g2239 ( 
.A(n_2215),
.B(n_2205),
.C(n_2211),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2222),
.B(n_2194),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2227),
.B(n_2180),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_L g2242 ( 
.A(n_2213),
.B(n_2203),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2227),
.B(n_1912),
.Y(n_2243)
);

NAND4xp25_ASAP7_75t_L g2244 ( 
.A(n_2213),
.B(n_1965),
.C(n_1978),
.D(n_1909),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2210),
.B(n_2134),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2219),
.Y(n_2246)
);

NOR3x1_ASAP7_75t_L g2247 ( 
.A(n_2231),
.B(n_2230),
.C(n_2217),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2237),
.B(n_2210),
.Y(n_2248)
);

AOI211xp5_ASAP7_75t_L g2249 ( 
.A1(n_2234),
.A2(n_2223),
.B(n_2211),
.C(n_2221),
.Y(n_2249)
);

AOI211xp5_ASAP7_75t_SL g2250 ( 
.A1(n_2232),
.A2(n_2221),
.B(n_2219),
.C(n_2226),
.Y(n_2250)
);

AOI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_2239),
.A2(n_2229),
.B(n_2208),
.Y(n_2251)
);

NAND4xp25_ASAP7_75t_L g2252 ( 
.A(n_2233),
.B(n_2208),
.C(n_2226),
.D(n_2220),
.Y(n_2252)
);

AOI22xp33_ASAP7_75t_SL g2253 ( 
.A1(n_2241),
.A2(n_2218),
.B1(n_2225),
.B2(n_2220),
.Y(n_2253)
);

AOI32xp33_ASAP7_75t_L g2254 ( 
.A1(n_2241),
.A2(n_2218),
.A3(n_2224),
.B1(n_1879),
.B2(n_1881),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_L g2255 ( 
.A(n_2242),
.B(n_1913),
.Y(n_2255)
);

AOI321xp33_ASAP7_75t_L g2256 ( 
.A1(n_2236),
.A2(n_1886),
.A3(n_1885),
.B1(n_1901),
.B2(n_1845),
.C(n_1843),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_L g2257 ( 
.A(n_2244),
.B(n_1913),
.Y(n_2257)
);

OAI211xp5_ASAP7_75t_SL g2258 ( 
.A1(n_2240),
.A2(n_2134),
.B(n_2011),
.C(n_2018),
.Y(n_2258)
);

NOR3x1_ASAP7_75t_L g2259 ( 
.A(n_2238),
.B(n_1994),
.C(n_1939),
.Y(n_2259)
);

NAND3xp33_ASAP7_75t_SL g2260 ( 
.A(n_2235),
.B(n_1976),
.C(n_1943),
.Y(n_2260)
);

AOI211xp5_ASAP7_75t_L g2261 ( 
.A1(n_2246),
.A2(n_1845),
.B(n_1886),
.C(n_1885),
.Y(n_2261)
);

AOI22xp5_ASAP7_75t_L g2262 ( 
.A1(n_2249),
.A2(n_2245),
.B1(n_2243),
.B2(n_2019),
.Y(n_2262)
);

AOI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_2248),
.A2(n_2258),
.B1(n_2251),
.B2(n_2255),
.Y(n_2263)
);

AOI211x1_ASAP7_75t_L g2264 ( 
.A1(n_2252),
.A2(n_2089),
.B(n_2084),
.C(n_2074),
.Y(n_2264)
);

INVx1_ASAP7_75t_SL g2265 ( 
.A(n_2253),
.Y(n_2265)
);

XNOR2xp5_ASAP7_75t_L g2266 ( 
.A(n_2260),
.B(n_1926),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2259),
.Y(n_2267)
);

INVxp67_ASAP7_75t_L g2268 ( 
.A(n_2250),
.Y(n_2268)
);

AOI22xp33_ASAP7_75t_L g2269 ( 
.A1(n_2257),
.A2(n_1906),
.B1(n_1901),
.B2(n_1872),
.Y(n_2269)
);

NAND2xp33_ASAP7_75t_L g2270 ( 
.A(n_2254),
.B(n_2074),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2256),
.B(n_2019),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2266),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2267),
.Y(n_2273)
);

NAND3xp33_ASAP7_75t_L g2274 ( 
.A(n_2268),
.B(n_2263),
.C(n_2270),
.Y(n_2274)
);

OA21x2_ASAP7_75t_L g2275 ( 
.A1(n_2268),
.A2(n_2247),
.B(n_2076),
.Y(n_2275)
);

NAND3x1_ASAP7_75t_L g2276 ( 
.A(n_2262),
.B(n_2261),
.C(n_2002),
.Y(n_2276)
);

AOI22x1_ASAP7_75t_L g2277 ( 
.A1(n_2265),
.A2(n_1994),
.B1(n_1838),
.B2(n_1904),
.Y(n_2277)
);

NAND4xp75_ASAP7_75t_L g2278 ( 
.A(n_2264),
.B(n_1993),
.C(n_2020),
.D(n_2013),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_2271),
.B(n_2042),
.Y(n_2279)
);

AOI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_2273),
.A2(n_2269),
.B1(n_2019),
.B2(n_1947),
.Y(n_2280)
);

NAND3xp33_ASAP7_75t_L g2281 ( 
.A(n_2275),
.B(n_2084),
.C(n_2045),
.Y(n_2281)
);

OAI322xp33_ASAP7_75t_L g2282 ( 
.A1(n_2274),
.A2(n_2064),
.A3(n_2070),
.B1(n_2069),
.B2(n_2048),
.C1(n_2047),
.C2(n_2067),
.Y(n_2282)
);

NOR3xp33_ASAP7_75t_SL g2283 ( 
.A(n_2275),
.B(n_2007),
.C(n_1899),
.Y(n_2283)
);

NOR4xp25_ASAP7_75t_L g2284 ( 
.A(n_2272),
.B(n_2049),
.C(n_2068),
.D(n_2076),
.Y(n_2284)
);

OAI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_2276),
.A2(n_2068),
.B1(n_2056),
.B2(n_2042),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2279),
.Y(n_2286)
);

NAND4xp25_ASAP7_75t_L g2287 ( 
.A(n_2279),
.B(n_1891),
.C(n_1926),
.D(n_1947),
.Y(n_2287)
);

INVx3_ASAP7_75t_SL g2288 ( 
.A(n_2286),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_2283),
.Y(n_2289)
);

INVx1_ASAP7_75t_SL g2290 ( 
.A(n_2280),
.Y(n_2290)
);

OAI211xp5_ASAP7_75t_SL g2291 ( 
.A1(n_2281),
.A2(n_2284),
.B(n_2285),
.C(n_2287),
.Y(n_2291)
);

BUFx2_ASAP7_75t_L g2292 ( 
.A(n_2288),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_2289),
.Y(n_2293)
);

INVx2_ASAP7_75t_SL g2294 ( 
.A(n_2292),
.Y(n_2294)
);

AO21x2_ASAP7_75t_L g2295 ( 
.A1(n_2293),
.A2(n_2291),
.B(n_2290),
.Y(n_2295)
);

HB1xp67_ASAP7_75t_L g2296 ( 
.A(n_2295),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2294),
.Y(n_2297)
);

HB1xp67_ASAP7_75t_L g2298 ( 
.A(n_2295),
.Y(n_2298)
);

INVx2_ASAP7_75t_SL g2299 ( 
.A(n_2297),
.Y(n_2299)
);

OAI21xp5_ASAP7_75t_L g2300 ( 
.A1(n_2296),
.A2(n_2277),
.B(n_2278),
.Y(n_2300)
);

AOI21xp33_ASAP7_75t_SL g2301 ( 
.A1(n_2299),
.A2(n_2298),
.B(n_2300),
.Y(n_2301)
);

OAI22xp5_ASAP7_75t_SL g2302 ( 
.A1(n_2299),
.A2(n_2277),
.B1(n_2282),
.B2(n_1838),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2302),
.A2(n_2056),
.B1(n_2002),
.B2(n_2019),
.Y(n_2303)
);

AOI221xp5_ASAP7_75t_L g2304 ( 
.A1(n_2303),
.A2(n_2301),
.B1(n_2002),
.B2(n_2007),
.C(n_2009),
.Y(n_2304)
);

AOI211xp5_ASAP7_75t_L g2305 ( 
.A1(n_2304),
.A2(n_1838),
.B(n_2034),
.C(n_1904),
.Y(n_2305)
);


endmodule