module fake_netlist_6_1648_n_669 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_669);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_669;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_327;
wire n_369;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_621;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_647;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_252;
wire n_228;
wire n_594;
wire n_565;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_608;
wire n_261;
wire n_527;
wire n_620;
wire n_420;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_655;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_47),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_21),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_120),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_2),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

BUFx10_ASAP7_75t_L g141 ( 
.A(n_38),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_5),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_113),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_27),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_17),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_20),
.B(n_2),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_18),
.Y(n_149)
);

NOR2xp67_ASAP7_75t_L g150 ( 
.A(n_3),
.B(n_130),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_18),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_58),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_50),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_28),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_87),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_61),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_33),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_51),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_60),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_12),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_119),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_46),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_63),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_16),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_101),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_99),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_30),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_77),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_59),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_14),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_82),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_137),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

OAI22x1_ASAP7_75t_R g188 ( 
.A1(n_180),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_137),
.Y(n_190)
);

AND2x4_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_22),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

BUFx8_ASAP7_75t_SL g193 ( 
.A(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_0),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_1),
.Y(n_198)
);

OAI21x1_ASAP7_75t_L g199 ( 
.A1(n_138),
.A2(n_143),
.B(n_140),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_4),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_131),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_4),
.B(n_5),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_149),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_6),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g206 ( 
.A(n_138),
.B(n_140),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_133),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_147),
.B(n_7),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_143),
.B(n_8),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_9),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_148),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_154),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_159),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_150),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_176),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_136),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_219),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_224),
.B(n_179),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_164),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_134),
.Y(n_238)
);

AND3x2_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_182),
.C(n_181),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_142),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_135),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_191),
.B(n_139),
.Y(n_243)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_224),
.B(n_145),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_205),
.A2(n_146),
.B1(n_177),
.B2(n_175),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_187),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_194),
.A2(n_153),
.B1(n_155),
.B2(n_171),
.Y(n_254)
);

AND2x6_ASAP7_75t_L g255 ( 
.A(n_205),
.B(n_156),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_214),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_200),
.A2(n_187),
.B1(n_217),
.B2(n_201),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_187),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_209),
.B(n_157),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_225),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_260),
.Y(n_266)
);

OR2x6_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_218),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_253),
.B(n_218),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_263),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_186),
.Y(n_270)
);

OAI221xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_211),
.B1(n_210),
.B2(n_183),
.C(n_190),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_201),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_235),
.A2(n_203),
.B1(n_190),
.B2(n_183),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_240),
.B(n_216),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_257),
.B(n_184),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_216),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_206),
.Y(n_279)
);

OR2x6_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_259),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_187),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_254),
.B(n_184),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_204),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_233),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_255),
.A2(n_203),
.B1(n_202),
.B2(n_166),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_185),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_232),
.Y(n_289)
);

AND2x6_ASAP7_75t_L g290 ( 
.A(n_232),
.B(n_160),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_234),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_255),
.A2(n_202),
.B1(n_199),
.B2(n_192),
.Y(n_292)
);

AO22x2_ASAP7_75t_L g293 ( 
.A1(n_226),
.A2(n_188),
.B1(n_215),
.B2(n_168),
.Y(n_293)
);

NOR3xp33_ASAP7_75t_L g294 ( 
.A(n_234),
.B(n_167),
.C(n_161),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_247),
.B(n_185),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_192),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_255),
.A2(n_202),
.B1(n_173),
.B2(n_178),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_233),
.B(n_196),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_250),
.A2(n_202),
.B1(n_199),
.B2(n_208),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_256),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_244),
.B(n_170),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_239),
.B(n_193),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_251),
.B(n_222),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_230),
.A2(n_208),
.B1(n_197),
.B2(n_189),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_262),
.B(n_189),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_244),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_230),
.A2(n_197),
.B1(n_222),
.B2(n_188),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_226),
.Y(n_311)
);

BUFx12f_ASAP7_75t_L g312 ( 
.A(n_267),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_265),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_270),
.B(n_215),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_283),
.B(n_228),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_286),
.A2(n_242),
.B1(n_231),
.B2(n_252),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_279),
.B(n_227),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_262),
.Y(n_319)
);

NAND2x1p5_ASAP7_75t_L g320 ( 
.A(n_266),
.B(n_227),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_288),
.A2(n_248),
.B(n_245),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_281),
.B(n_222),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_229),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_13),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_276),
.B(n_13),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_296),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_297),
.A2(n_237),
.B(n_229),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_295),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_23),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_298),
.B(n_24),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_311),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_286),
.B(n_25),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_275),
.B(n_14),
.Y(n_335)
);

NAND2x1_ASAP7_75t_L g336 ( 
.A(n_287),
.B(n_26),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_282),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_299),
.A2(n_71),
.B(n_128),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_277),
.A2(n_68),
.B(n_126),
.Y(n_339)
);

NAND3xp33_ASAP7_75t_L g340 ( 
.A(n_274),
.B(n_15),
.C(n_16),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_L g341 ( 
.A1(n_271),
.A2(n_15),
.B(n_17),
.C(n_19),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_264),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_269),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_306),
.A2(n_72),
.B(n_29),
.Y(n_344)
);

A2O1A1Ixp33_ASAP7_75t_L g345 ( 
.A1(n_274),
.A2(n_19),
.B(n_31),
.C(n_32),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_309),
.B(n_34),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_300),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_290),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_310),
.B(n_39),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_284),
.A2(n_40),
.B(n_41),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_308),
.A2(n_42),
.B(n_43),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_290),
.B(n_307),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_44),
.Y(n_354)
);

AO22x1_ASAP7_75t_L g355 ( 
.A1(n_294),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_307),
.A2(n_302),
.B(n_285),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_280),
.B(n_268),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_272),
.A2(n_52),
.B(n_53),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_272),
.A2(n_54),
.B(n_55),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_290),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_280),
.B(n_56),
.Y(n_361)
);

BUFx4f_ASAP7_75t_L g362 ( 
.A(n_280),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_268),
.B(n_57),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_305),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_334),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_314),
.A2(n_293),
.B(n_267),
.C(n_65),
.Y(n_366)
);

NAND2x1p5_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_62),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_333),
.Y(n_368)
);

OAI21x1_ASAP7_75t_L g369 ( 
.A1(n_356),
.A2(n_64),
.B(n_66),
.Y(n_369)
);

OAI21x1_ASAP7_75t_L g370 ( 
.A1(n_321),
.A2(n_67),
.B(n_75),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_329),
.B(n_293),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_316),
.B(n_267),
.Y(n_372)
);

OAI21x1_ASAP7_75t_L g373 ( 
.A1(n_328),
.A2(n_76),
.B(n_78),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_79),
.Y(n_374)
);

AO21x1_ASAP7_75t_L g375 ( 
.A1(n_330),
.A2(n_80),
.B(n_81),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_337),
.B(n_83),
.Y(n_376)
);

AOI211x1_ASAP7_75t_L g377 ( 
.A1(n_340),
.A2(n_84),
.B(n_88),
.C(n_90),
.Y(n_377)
);

NOR2x1_ASAP7_75t_SL g378 ( 
.A(n_360),
.B(n_92),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_326),
.B(n_93),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_312),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_323),
.A2(n_94),
.B(n_95),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_357),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_342),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_362),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_318),
.B(n_96),
.Y(n_386)
);

AO21x1_ASAP7_75t_L g387 ( 
.A1(n_330),
.A2(n_97),
.B(n_98),
.Y(n_387)
);

A2O1A1Ixp33_ASAP7_75t_L g388 ( 
.A1(n_334),
.A2(n_102),
.B(n_103),
.C(n_104),
.Y(n_388)
);

OA21x2_ASAP7_75t_L g389 ( 
.A1(n_323),
.A2(n_106),
.B(n_107),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_319),
.A2(n_108),
.B(n_109),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_318),
.A2(n_110),
.B(n_111),
.Y(n_391)
);

OA22x2_ASAP7_75t_L g392 ( 
.A1(n_350),
.A2(n_331),
.B1(n_335),
.B2(n_322),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_331),
.B(n_114),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_117),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_353),
.A2(n_118),
.B(n_121),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_320),
.B(n_123),
.Y(n_396)
);

AOI211x1_ASAP7_75t_L g397 ( 
.A1(n_352),
.A2(n_125),
.B(n_129),
.C(n_343),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_325),
.B(n_327),
.Y(n_398)
);

NAND2x1_ASAP7_75t_L g399 ( 
.A(n_347),
.B(n_349),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_317),
.B(n_347),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_313),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_320),
.B(n_362),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_341),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_354),
.B(n_346),
.Y(n_404)
);

AOI211x1_ASAP7_75t_L g405 ( 
.A1(n_355),
.A2(n_339),
.B(n_351),
.C(n_338),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_348),
.A2(n_344),
.B(n_345),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_358),
.A2(n_314),
.B1(n_334),
.B2(n_331),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_359),
.B(n_329),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_332),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_315),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_314),
.A2(n_334),
.B1(n_330),
.B2(n_331),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_382),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_365),
.B(n_411),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_L g414 ( 
.A1(n_411),
.A2(n_365),
.B1(n_371),
.B2(n_372),
.Y(n_414)
);

AO31x2_ASAP7_75t_L g415 ( 
.A1(n_407),
.A2(n_375),
.A3(n_387),
.B(n_406),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_408),
.A2(n_369),
.B(n_386),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_368),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_383),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_398),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_409),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_384),
.B(n_371),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_374),
.A2(n_400),
.B(n_407),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_398),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_385),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_410),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_364),
.B(n_380),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_364),
.Y(n_427)
);

AO32x2_ASAP7_75t_L g428 ( 
.A1(n_397),
.A2(n_392),
.A3(n_377),
.B1(n_405),
.B2(n_403),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_401),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_400),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_394),
.A2(n_393),
.B1(n_392),
.B2(n_404),
.Y(n_431)
);

AND2x6_ASAP7_75t_L g432 ( 
.A(n_393),
.B(n_396),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_399),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_366),
.B(n_376),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_386),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_381),
.A2(n_379),
.B(n_395),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_367),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_367),
.Y(n_438)
);

OAI21x1_ASAP7_75t_SL g439 ( 
.A1(n_378),
.A2(n_391),
.B(n_390),
.Y(n_439)
);

O2A1O1Ixp33_ASAP7_75t_SL g440 ( 
.A1(n_388),
.A2(n_389),
.B(n_370),
.C(n_373),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_382),
.Y(n_441)
);

AO21x2_ASAP7_75t_L g442 ( 
.A1(n_406),
.A2(n_393),
.B(n_386),
.Y(n_442)
);

OAI21x1_ASAP7_75t_SL g443 ( 
.A1(n_378),
.A2(n_387),
.B(n_375),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_365),
.B(n_314),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_368),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_386),
.A2(n_408),
.B(n_393),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_371),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_368),
.Y(n_449)
);

AO21x2_ASAP7_75t_L g450 ( 
.A1(n_406),
.A2(n_393),
.B(n_386),
.Y(n_450)
);

AO21x2_ASAP7_75t_L g451 ( 
.A1(n_406),
.A2(n_393),
.B(n_386),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_L g452 ( 
.A1(n_411),
.A2(n_314),
.B1(n_334),
.B2(n_407),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_368),
.Y(n_453)
);

AO21x1_ASAP7_75t_SL g454 ( 
.A1(n_393),
.A2(n_334),
.B(n_331),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_418),
.Y(n_455)
);

BUFx10_ASAP7_75t_L g456 ( 
.A(n_424),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_419),
.Y(n_457)
);

NOR2x1_ASAP7_75t_SL g458 ( 
.A(n_454),
.B(n_435),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_452),
.B(n_444),
.Y(n_460)
);

NAND2x1_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_439),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_420),
.B(n_434),
.Y(n_462)
);

BUFx10_ASAP7_75t_L g463 ( 
.A(n_444),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_417),
.Y(n_464)
);

AO21x2_ASAP7_75t_L g465 ( 
.A1(n_447),
.A2(n_422),
.B(n_443),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_448),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_445),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_441),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_446),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_441),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_415),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_449),
.Y(n_472)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_436),
.A2(n_431),
.B(n_416),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_427),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_421),
.B(n_448),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_430),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_429),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_413),
.B(n_414),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_425),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_433),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_433),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_420),
.A2(n_414),
.B1(n_432),
.B2(n_426),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_426),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_412),
.Y(n_485)
);

OAI21x1_ASAP7_75t_L g486 ( 
.A1(n_416),
.A2(n_438),
.B(n_440),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_438),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_428),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_428),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_432),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_415),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_455),
.Y(n_492)
);

INVxp67_ASAP7_75t_R g493 ( 
.A(n_484),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_432),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_460),
.B(n_428),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_462),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_415),
.Y(n_497)
);

OR2x6_ASAP7_75t_L g498 ( 
.A(n_461),
.B(n_432),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_457),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_463),
.B(n_442),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_462),
.B(n_442),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_459),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_459),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_456),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_479),
.B(n_450),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_466),
.B(n_450),
.Y(n_506)
);

AND2x2_ASAP7_75t_SL g507 ( 
.A(n_483),
.B(n_491),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_490),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_477),
.B(n_472),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_477),
.B(n_451),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_472),
.B(n_451),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_478),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_478),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_480),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_481),
.B(n_482),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_463),
.B(n_480),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_464),
.Y(n_517)
);

NOR2x1_ASAP7_75t_L g518 ( 
.A(n_465),
.B(n_461),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_463),
.B(n_476),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_464),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_488),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_463),
.B(n_467),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_489),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_456),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_467),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_469),
.B(n_476),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_465),
.B(n_471),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_489),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_468),
.B(n_470),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_499),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_R g532 ( 
.A(n_530),
.B(n_516),
.Y(n_532)
);

AND2x4_ASAP7_75t_SL g533 ( 
.A(n_516),
.B(n_456),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_499),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_496),
.B(n_474),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_496),
.B(n_465),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_519),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_495),
.B(n_473),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_502),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_520),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_495),
.B(n_473),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_504),
.B(n_456),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_505),
.B(n_469),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_520),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_504),
.B(n_485),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_497),
.B(n_487),
.Y(n_546)
);

NOR2x1_ASAP7_75t_L g547 ( 
.A(n_525),
.B(n_514),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_525),
.Y(n_548)
);

NAND3xp33_ASAP7_75t_L g549 ( 
.A(n_500),
.B(n_487),
.C(n_482),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_505),
.B(n_486),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_523),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_519),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_523),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_501),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_522),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_509),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_522),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_524),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_525),
.B(n_481),
.C(n_458),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_554),
.B(n_501),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_554),
.B(n_546),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_540),
.B(n_507),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_531),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_537),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_546),
.B(n_506),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_548),
.B(n_494),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_536),
.B(n_506),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_548),
.B(n_494),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_537),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_536),
.B(n_528),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_544),
.B(n_528),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_532),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_543),
.B(n_510),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_531),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_535),
.B(n_494),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_533),
.B(n_556),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_552),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_552),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_555),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_543),
.B(n_510),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_549),
.A2(n_518),
.B(n_507),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_533),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_555),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_547),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_542),
.B(n_494),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_551),
.B(n_507),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_557),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_553),
.B(n_511),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_550),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_534),
.B(n_511),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_538),
.B(n_529),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_589),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_589),
.B(n_538),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_570),
.B(n_550),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_572),
.B(n_545),
.Y(n_595)
);

NOR5xp2_ASAP7_75t_L g596 ( 
.A(n_572),
.B(n_559),
.C(n_558),
.D(n_557),
.E(n_492),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_564),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_569),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_577),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_563),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_566),
.B(n_513),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_578),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_579),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_567),
.B(n_541),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_561),
.B(n_571),
.Y(n_605)
);

NAND2x1_ASAP7_75t_L g606 ( 
.A(n_584),
.B(n_498),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_573),
.B(n_541),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_583),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_576),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_582),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_609),
.B(n_576),
.Y(n_611)
);

INVxp67_ASAP7_75t_SL g612 ( 
.A(n_592),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_597),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_592),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_598),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_599),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_602),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_603),
.Y(n_618)
);

A2O1A1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_596),
.A2(n_581),
.B(n_575),
.C(n_585),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_600),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_613),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_615),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_619),
.A2(n_595),
.B1(n_568),
.B2(n_566),
.Y(n_623)
);

NOR2x1_ASAP7_75t_SL g624 ( 
.A(n_614),
.B(n_605),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_616),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_617),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_620),
.B(n_594),
.Y(n_627)
);

AOI221xp5_ASAP7_75t_L g628 ( 
.A1(n_623),
.A2(n_619),
.B1(n_618),
.B2(n_581),
.C(n_612),
.Y(n_628)
);

OAI221xp5_ASAP7_75t_SL g629 ( 
.A1(n_621),
.A2(n_610),
.B1(n_612),
.B2(n_593),
.C(n_607),
.Y(n_629)
);

AOI221xp5_ASAP7_75t_L g630 ( 
.A1(n_622),
.A2(n_593),
.B1(n_608),
.B2(n_601),
.C(n_611),
.Y(n_630)
);

NAND3xp33_ASAP7_75t_L g631 ( 
.A(n_625),
.B(n_596),
.C(n_606),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_626),
.A2(n_627),
.B1(n_609),
.B2(n_611),
.Y(n_632)
);

NOR3xp33_ASAP7_75t_L g633 ( 
.A(n_624),
.B(n_508),
.C(n_568),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_628),
.B(n_604),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_631),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_633),
.B(n_560),
.Y(n_636)
);

NAND3xp33_ASAP7_75t_L g637 ( 
.A(n_629),
.B(n_587),
.C(n_562),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_635),
.Y(n_638)
);

NAND3xp33_ASAP7_75t_L g639 ( 
.A(n_637),
.B(n_630),
.C(n_632),
.Y(n_639)
);

NOR2x1_ASAP7_75t_L g640 ( 
.A(n_634),
.B(n_503),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_638),
.B(n_636),
.Y(n_641)
);

NAND3x2_ASAP7_75t_L g642 ( 
.A(n_639),
.B(n_586),
.C(n_565),
.Y(n_642)
);

NOR3xp33_ASAP7_75t_L g643 ( 
.A(n_640),
.B(n_508),
.C(n_514),
.Y(n_643)
);

NOR3xp33_ASAP7_75t_L g644 ( 
.A(n_641),
.B(n_508),
.C(n_521),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_643),
.B(n_591),
.Y(n_645)
);

XNOR2x1_ASAP7_75t_L g646 ( 
.A(n_642),
.B(n_498),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_641),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_SL g648 ( 
.A(n_641),
.B(n_527),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_641),
.B(n_580),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_647),
.A2(n_648),
.B(n_646),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_649),
.Y(n_651)
);

NAND3xp33_ASAP7_75t_L g652 ( 
.A(n_644),
.B(n_517),
.C(n_526),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_645),
.A2(n_580),
.B1(n_573),
.B2(n_588),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g654 ( 
.A(n_647),
.B(n_458),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_649),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_651),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_SL g657 ( 
.A1(n_655),
.A2(n_498),
.B1(n_508),
.B2(n_517),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_650),
.A2(n_574),
.B1(n_590),
.B2(n_558),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_654),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_656),
.A2(n_652),
.B(n_653),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_658),
.A2(n_493),
.B(n_521),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_659),
.A2(n_493),
.B(n_526),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_660),
.A2(n_657),
.B(n_527),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_662),
.A2(n_515),
.B1(n_492),
.B2(n_509),
.Y(n_664)
);

XOR2xp5_ASAP7_75t_L g665 ( 
.A(n_661),
.B(n_515),
.Y(n_665)
);

AOI221xp5_ASAP7_75t_L g666 ( 
.A1(n_663),
.A2(n_515),
.B1(n_513),
.B2(n_512),
.C(n_539),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_666),
.B(n_665),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_667),
.B(n_664),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_668),
.A2(n_515),
.B1(n_512),
.B2(n_534),
.Y(n_669)
);


endmodule