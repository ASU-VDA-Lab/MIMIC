module fake_jpeg_22894_n_284 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_149;
wire n_48;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_30),
.Y(n_47)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_38),
.B1(n_29),
.B2(n_18),
.Y(n_51)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_27),
.B1(n_29),
.B2(n_19),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_29),
.B1(n_38),
.B2(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_47),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_52),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_29),
.B1(n_32),
.B2(n_18),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_55),
.B1(n_50),
.B2(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_25),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_21),
.Y(n_84)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_62),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_25),
.C(n_23),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_18),
.B1(n_35),
.B2(n_38),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_38),
.B1(n_37),
.B2(n_35),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_35),
.B1(n_29),
.B2(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_32),
.B1(n_26),
.B2(n_24),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_0),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_84),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_31),
.B1(n_20),
.B2(n_26),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_86),
.B1(n_28),
.B2(n_70),
.Y(n_112)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_80),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_17),
.Y(n_96)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_82),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_85),
.B(n_49),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_24),
.B1(n_20),
.B2(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_92),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_54),
.C(n_49),
.Y(n_92)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_96),
.B(n_101),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_53),
.B(n_17),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_98),
.A2(n_110),
.B(n_83),
.Y(n_139)
);

OA22x2_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_40),
.B1(n_16),
.B2(n_17),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_73),
.B1(n_60),
.B2(n_65),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_77),
.Y(n_132)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_109),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_61),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_72),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_54),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_82),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_124),
.B1(n_138),
.B2(n_99),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_118),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_70),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_121),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_78),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_78),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_122),
.B(n_125),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_59),
.B1(n_79),
.B2(n_67),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_126),
.B(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_94),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_132),
.B(n_139),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_134),
.B1(n_136),
.B2(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_103),
.A2(n_67),
.B1(n_80),
.B2(n_83),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_99),
.B1(n_113),
.B2(n_101),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_126),
.B1(n_139),
.B2(n_121),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_105),
.B(n_113),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_143),
.A2(n_154),
.B(n_170),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_112),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_149),
.C(n_155),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_157),
.B1(n_164),
.B2(n_140),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_99),
.B1(n_107),
.B2(n_88),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_148),
.A2(n_150),
.B1(n_152),
.B2(n_123),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_88),
.C(n_97),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_97),
.B1(n_77),
.B2(n_87),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_94),
.B(n_17),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_40),
.C(n_108),
.Y(n_155)
);

AND2x4_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_40),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_SL g189 ( 
.A(n_156),
.B(n_165),
.C(n_168),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_124),
.A2(n_91),
.B1(n_106),
.B2(n_90),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_91),
.B1(n_95),
.B2(n_28),
.Y(n_164)
);

OA21x2_ASAP7_75t_SL g165 ( 
.A1(n_119),
.A2(n_17),
.B(n_1),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_119),
.B(n_17),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_114),
.Y(n_178)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_118),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_SL g168 ( 
.A1(n_120),
.A2(n_22),
.B(n_21),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_119),
.A2(n_16),
.B(n_48),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_116),
.B(n_0),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_SL g196 ( 
.A1(n_171),
.A2(n_0),
.B(n_22),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_196),
.B1(n_156),
.B2(n_160),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_135),
.Y(n_174)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_175),
.B(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_161),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_169),
.Y(n_179)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_182),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_191),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_151),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_136),
.C(n_125),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_144),
.C(n_154),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_11),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_209),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_148),
.Y(n_201)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_197),
.A2(n_160),
.B(n_143),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_211),
.B(n_216),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_215),
.C(n_181),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_195),
.A2(n_166),
.B1(n_147),
.B2(n_153),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_217),
.B1(n_175),
.B2(n_189),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_208),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_190),
.B(n_22),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_22),
.B(n_21),
.C(n_16),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_209),
.B(n_2),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_1),
.B(n_2),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_178),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_189),
.A2(n_1),
.B(n_2),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_206),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_203),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_201),
.A2(n_185),
.B1(n_184),
.B2(n_177),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_230),
.B1(n_229),
.B2(n_219),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_200),
.B(n_192),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_184),
.B1(n_176),
.B2(n_187),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_228),
.A2(n_216),
.B(n_204),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_211),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_198),
.A2(n_173),
.B1(n_48),
.B2(n_16),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_232),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_212),
.B(n_3),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_3),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_233),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_238),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_202),
.B(n_214),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_215),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_221),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_225),
.A2(n_230),
.B1(n_224),
.B2(n_227),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_218),
.B1(n_48),
.B2(n_6),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_234),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_233),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_254),
.Y(n_261)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_253),
.Y(n_260)
);

NOR3xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_234),
.C(n_208),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_242),
.B(n_221),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_256),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_258),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_4),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_249),
.A2(n_240),
.B(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_237),
.B(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_264),
.B(n_9),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_246),
.C(n_238),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_11),
.C(n_12),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_235),
.Y(n_268)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

AO21x1_ASAP7_75t_L g269 ( 
.A1(n_260),
.A2(n_5),
.B(n_6),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_265),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_11),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_273),
.B1(n_274),
.B2(n_262),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_261),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_271),
.Y(n_275)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_278),
.B(n_273),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_280),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_272),
.B1(n_262),
.B2(n_15),
.Y(n_280)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_13),
.C(n_14),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_281),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_15),
.Y(n_284)
);


endmodule