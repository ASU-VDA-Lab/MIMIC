module fake_netlist_5_1449_n_1227 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1227);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1227;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_1194;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_1178;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_523;
wire n_268;
wire n_315;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_1161;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_1222;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_525;
wire n_493;
wire n_397;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_1191;
wire n_1198;
wire n_721;
wire n_998;
wire n_1157;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_1120;
wire n_915;
wire n_719;
wire n_372;
wire n_443;
wire n_293;
wire n_677;
wire n_244;
wire n_173;
wire n_859;
wire n_864;
wire n_1110;
wire n_951;
wire n_1121;
wire n_1203;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_314;
wire n_247;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_1179;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_1048;
wire n_932;
wire n_612;
wire n_1001;
wire n_516;
wire n_498;
wire n_385;
wire n_212;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_1195;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_1090;
wire n_757;
wire n_947;
wire n_1200;
wire n_307;
wire n_633;
wire n_1192;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1185;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_1032;
wire n_929;
wire n_981;
wire n_941;
wire n_1143;
wire n_804;
wire n_867;
wire n_186;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_171;
wire n_1182;
wire n_756;
wire n_1145;
wire n_943;
wire n_524;
wire n_878;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_1049;
wire n_992;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_1163;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_1108;
wire n_908;
wire n_449;
wire n_325;
wire n_1100;
wire n_1207;
wire n_1214;
wire n_862;
wire n_1016;
wire n_724;
wire n_856;
wire n_546;
wire n_900;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_1169;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_1221;
wire n_654;
wire n_370;
wire n_1172;
wire n_1095;
wire n_1096;
wire n_976;
wire n_234;
wire n_343;
wire n_428;
wire n_379;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_1208;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_1168;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1201;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_995;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_1176;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_1149;
wire n_882;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_1225;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_1073;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_181;
wire n_436;
wire n_962;
wire n_1219;
wire n_1204;
wire n_1215;
wire n_1216;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_1171;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_1218;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1188;
wire n_1030;
wire n_1223;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_1165;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_1177;
wire n_680;
wire n_974;
wire n_432;
wire n_553;
wire n_395;
wire n_727;
wire n_901;
wire n_839;
wire n_311;
wire n_813;
wire n_1159;
wire n_1210;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_328;
wire n_214;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_1167;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_928;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_482;
wire n_342;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_1173;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_1193;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1122;
wire n_1111;
wire n_1197;
wire n_1211;
wire n_1226;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_1041;
wire n_989;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_834;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1187;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_1164;
wire n_420;
wire n_630;
wire n_1202;
wire n_489;
wire n_632;
wire n_699;
wire n_1174;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_1058;
wire n_846;
wire n_465;
wire n_838;
wire n_358;
wire n_874;
wire n_362;
wire n_876;
wire n_170;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_349;
wire n_585;
wire n_1106;
wire n_1190;
wire n_1224;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_1052;
wire n_963;
wire n_954;
wire n_627;
wire n_1116;
wire n_1212;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_1175;
wire n_861;
wire n_534;
wire n_948;
wire n_1183;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_1217;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_176;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_182;
wire n_1005;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_679;
wire n_425;
wire n_513;
wire n_237;
wire n_407;
wire n_527;
wire n_647;
wire n_710;
wire n_707;
wire n_795;
wire n_695;
wire n_832;
wire n_180;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1220;
wire n_1044;
wire n_1205;
wire n_346;
wire n_937;
wire n_1209;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1072;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_1027;
wire n_971;
wire n_490;
wire n_805;
wire n_1156;
wire n_910;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_233;
wire n_686;
wire n_572;
wire n_366;
wire n_205;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_1037;
wire n_1160;
wire n_202;
wire n_1080;
wire n_266;
wire n_1162;
wire n_491;
wire n_272;
wire n_1074;
wire n_427;
wire n_1199;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_1181;
wire n_1196;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_931;
wire n_870;
wire n_334;
wire n_599;
wire n_766;
wire n_952;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_1213;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_1004;
wire n_935;
wire n_1186;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_1184;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_1189;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_1180;
wire n_1206;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_1170;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_12),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_21),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_165),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_99),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_44),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_158),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_0),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_16),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_48),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_23),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_77),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_12),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_61),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_38),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_29),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_0),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_17),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_47),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_128),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_50),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_60),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_93),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_5),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_52),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_79),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_110),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_68),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_86),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_85),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_139),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_102),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_131),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_78),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_24),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_157),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_146),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_8),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_108),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_28),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_34),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_160),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_148),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_145),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_100),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_70),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_45),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_29),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_10),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_37),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_83),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_92),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_143),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_127),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_133),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_7),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_26),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_73),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_125),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_153),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_67),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_82),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_58),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_11),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_48),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_150),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_90),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_140),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_156),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_57),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_10),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_118),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_122),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_105),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_28),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_18),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_47),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_164),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_25),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_14),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_31),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_144),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_162),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_4),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_166),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_51),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_14),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_45),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_138),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_141),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_17),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_80),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_168),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_7),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_104),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_37),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_19),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_161),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_66),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_36),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_46),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_96),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_31),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_152),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_27),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_21),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_163),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_178),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_195),
.Y(n_293)
);

INVxp33_ASAP7_75t_SL g294 ( 
.A(n_179),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_220),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_180),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_172),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_196),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_199),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_196),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_201),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_224),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_234),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_206),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_267),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_290),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_224),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_198),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_198),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_170),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_170),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_170),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_217),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_182),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_170),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_170),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_283),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_228),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_222),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_283),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_223),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_179),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_228),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_240),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_281),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_255),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_229),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_186),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_193),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_281),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_231),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_175),
.Y(n_336)
);

BUFx6f_ASAP7_75t_SL g337 ( 
.A(n_240),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_194),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_255),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_232),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_258),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_247),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_259),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_282),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_266),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_254),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_279),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_282),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_262),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_284),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_184),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_187),
.B(n_1),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_266),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_263),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_264),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_174),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_184),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_176),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_171),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_239),
.B(n_1),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_188),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_189),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_191),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_191),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_181),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_240),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_190),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_197),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_255),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_202),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_204),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_210),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_226),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_183),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_200),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_236),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_280),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_241),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_280),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_243),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_299),
.B(n_187),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_185),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_322),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_322),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_311),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_367),
.B(n_185),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_313),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_297),
.B(n_192),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_297),
.B(n_192),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_313),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_316),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_298),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_316),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_300),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

NAND2x1_ASAP7_75t_L g401 ( 
.A(n_299),
.B(n_257),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_319),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_323),
.Y(n_403)
);

OR2x6_ASAP7_75t_L g404 ( 
.A(n_361),
.B(n_239),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_354),
.B(n_292),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_336),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_306),
.B(n_208),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_362),
.B(n_208),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_336),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_332),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_333),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_330),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_340),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_330),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_291),
.B(n_173),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_341),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_343),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_347),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_348),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_301),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_368),
.B(n_273),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_339),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_345),
.B(n_242),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_295),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_339),
.A2(n_242),
.B(n_249),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_369),
.B(n_250),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_304),
.B(n_177),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_370),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_300),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_381),
.B(n_175),
.Y(n_432)
);

AND2x2_ASAP7_75t_SL g433 ( 
.A(n_353),
.B(n_257),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_302),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_351),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_357),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_307),
.A2(n_248),
.B1(n_288),
.B2(n_270),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_358),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_372),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_373),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_374),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_L g444 ( 
.A(n_302),
.B(n_305),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_377),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_361),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_309),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_310),
.B(n_273),
.Y(n_449)
);

CKINVDCx8_ASAP7_75t_R g450 ( 
.A(n_358),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_338),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_439),
.B(n_364),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_443),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_417),
.A2(n_288),
.B1(n_286),
.B2(n_271),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_402),
.Y(n_455)
);

AND2x6_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_257),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_414),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_430),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_392),
.B(n_294),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_393),
.B(n_294),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_422),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_412),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_293),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_389),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_443),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_328),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_402),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_359),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_430),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_402),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_430),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_412),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_366),
.Y(n_473)
);

INVx6_ASAP7_75t_L g474 ( 
.A(n_430),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_405),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_405),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_405),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_414),
.Y(n_478)
);

BUFx10_ASAP7_75t_L g479 ( 
.A(n_417),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_424),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_433),
.B(n_256),
.C(n_252),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_425),
.B(n_305),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_429),
.B(n_375),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_425),
.B(n_433),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_424),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_443),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_SL g487 ( 
.A(n_439),
.B(n_380),
.Y(n_487)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_438),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_424),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_386),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_412),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_437),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_437),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_437),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_429),
.B(n_314),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_433),
.B(n_314),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_386),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_443),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_406),
.B(n_451),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_386),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_451),
.B(n_321),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_404),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_390),
.B(n_376),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_428),
.B(n_321),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_451),
.B(n_324),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_389),
.Y(n_506)
);

AND2x2_ASAP7_75t_SL g507 ( 
.A(n_444),
.B(n_257),
.Y(n_507)
);

OAI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_404),
.A2(n_380),
.B1(n_378),
.B2(n_365),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_414),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g510 ( 
.A1(n_404),
.A2(n_274),
.B1(n_289),
.B2(n_277),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_389),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_426),
.B(n_324),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_414),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_416),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_416),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_450),
.B(n_331),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_443),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_L g518 ( 
.A(n_383),
.B(n_331),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_450),
.B(n_335),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_422),
.Y(n_520)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_438),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_394),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_458),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_481),
.A2(n_404),
.B1(n_428),
.B2(n_382),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_484),
.B(n_404),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_462),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_471),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_458),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_474),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_512),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_481),
.A2(n_404),
.B1(n_428),
.B2(n_382),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_474),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_499),
.B(n_406),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_469),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_462),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_471),
.B(n_443),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_469),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_471),
.B(n_428),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_479),
.B(n_450),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_471),
.B(n_383),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_507),
.B(n_423),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_490),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_479),
.B(n_398),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_479),
.B(n_398),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_507),
.B(n_423),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_507),
.B(n_457),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_455),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_463),
.B(n_449),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_482),
.B(n_431),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_479),
.B(n_431),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_455),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_496),
.B(n_434),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_499),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_504),
.A2(n_427),
.B(n_449),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_474),
.B(n_382),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_462),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_472),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_466),
.B(n_406),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_459),
.B(n_434),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_474),
.Y(n_560)
);

NOR2xp67_ASAP7_75t_L g561 ( 
.A(n_503),
.B(n_436),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_467),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_460),
.B(n_335),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_467),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_472),
.B(n_440),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_490),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_468),
.B(n_473),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_461),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_470),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_461),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_510),
.B(n_448),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_472),
.Y(n_572)
);

NAND3xp33_ASAP7_75t_SL g573 ( 
.A(n_454),
.B(n_308),
.C(n_303),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_491),
.B(n_382),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_470),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_L g576 ( 
.A(n_456),
.B(n_255),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_508),
.B(n_342),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_491),
.B(n_440),
.Y(n_578)
);

AOI221xp5_ASAP7_75t_L g579 ( 
.A1(n_488),
.A2(n_238),
.B1(n_207),
.B2(n_245),
.C(n_230),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_L g580 ( 
.A(n_456),
.B(n_255),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_475),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_497),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_L g583 ( 
.A(n_456),
.B(n_255),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_508),
.B(n_342),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_475),
.Y(n_585)
);

NAND3xp33_ASAP7_75t_L g586 ( 
.A(n_483),
.B(n_350),
.C(n_346),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_476),
.Y(n_587)
);

BUFx5_ASAP7_75t_L g588 ( 
.A(n_456),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_476),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_491),
.B(n_440),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_502),
.B(n_448),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_502),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_509),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_509),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_497),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_500),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_495),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_509),
.B(n_514),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_509),
.B(n_416),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_477),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_500),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_501),
.B(n_346),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_505),
.B(n_350),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_518),
.A2(n_272),
.B1(n_356),
.B2(n_355),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_516),
.B(n_355),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_477),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_514),
.B(n_416),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_519),
.B(n_356),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_452),
.B(n_364),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_456),
.A2(n_409),
.B1(n_408),
.B2(n_427),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_520),
.B(n_408),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_456),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_456),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_522),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_522),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_487),
.B(n_365),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_480),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_514),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_480),
.Y(n_619)
);

O2A1O1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_485),
.A2(n_441),
.B(n_445),
.C(n_442),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_597),
.B(n_454),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_570),
.B(n_521),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_548),
.B(n_514),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_529),
.A2(n_506),
.B(n_464),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_553),
.A2(n_327),
.B1(n_329),
.B2(n_320),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_529),
.A2(n_506),
.B(n_464),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_525),
.A2(n_515),
.B(n_513),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_529),
.A2(n_506),
.B(n_464),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_541),
.A2(n_427),
.B(n_285),
.C(n_287),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_540),
.B(n_558),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_558),
.B(n_513),
.Y(n_631)
);

A2O1A1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_545),
.A2(n_268),
.B(n_515),
.C(n_408),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_533),
.B(n_485),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_611),
.B(n_378),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_533),
.B(n_489),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_527),
.B(n_489),
.Y(n_636)
);

OAI321xp33_ASAP7_75t_L g637 ( 
.A1(n_579),
.A2(n_289),
.A3(n_274),
.B1(n_277),
.B2(n_413),
.C(n_435),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_527),
.B(n_492),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_565),
.B(n_411),
.Y(n_639)
);

NOR2x1p5_ASAP7_75t_SL g640 ( 
.A(n_588),
.B(n_492),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_565),
.B(n_411),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_568),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_527),
.B(n_493),
.Y(n_643)
);

NOR2x1p5_ASAP7_75t_L g644 ( 
.A(n_573),
.B(n_334),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_619),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_619),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_532),
.A2(n_506),
.B(n_464),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_571),
.A2(n_493),
.B1(n_494),
.B2(n_257),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_532),
.B(n_494),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_532),
.B(n_453),
.Y(n_650)
);

AO21x1_ASAP7_75t_L g651 ( 
.A1(n_546),
.A2(n_409),
.B(n_408),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_560),
.A2(n_511),
.B(n_465),
.Y(n_652)
);

AOI21xp33_ASAP7_75t_L g653 ( 
.A1(n_554),
.A2(n_401),
.B(n_441),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_560),
.A2(n_511),
.B(n_465),
.Y(n_654)
);

AOI21x1_ASAP7_75t_L g655 ( 
.A1(n_538),
.A2(n_536),
.B(n_574),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_560),
.A2(n_555),
.B(n_572),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_593),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_617),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_530),
.B(n_567),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_572),
.A2(n_511),
.B(n_465),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_523),
.A2(n_511),
.B(n_409),
.Y(n_661)
);

O2A1O1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_552),
.A2(n_442),
.B(n_445),
.C(n_413),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_535),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_605),
.A2(n_409),
.B(n_218),
.C(n_235),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_549),
.A2(n_418),
.B(n_435),
.C(n_415),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_594),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_567),
.B(n_344),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_543),
.B(n_349),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_578),
.A2(n_465),
.B(n_453),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_590),
.A2(n_465),
.B(n_453),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_617),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_549),
.A2(n_419),
.B(n_421),
.C(n_415),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_608),
.A2(n_253),
.B1(n_498),
.B2(n_486),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_550),
.B(n_396),
.Y(n_674)
);

O2A1O1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_523),
.A2(n_421),
.B(n_420),
.C(n_419),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_535),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_598),
.A2(n_486),
.B(n_453),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_591),
.B(n_453),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_559),
.B(n_325),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_610),
.A2(n_498),
.B(n_486),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_528),
.A2(n_498),
.B(n_486),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_547),
.Y(n_682)
);

CKINVDCx11_ASAP7_75t_R g683 ( 
.A(n_535),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_528),
.A2(n_498),
.B(n_486),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_565),
.A2(n_517),
.B1(n_498),
.B2(n_278),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_604),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_591),
.B(n_517),
.Y(n_687)
);

AOI33xp33_ASAP7_75t_L g688 ( 
.A1(n_611),
.A2(n_418),
.A3(n_420),
.B1(n_432),
.B2(n_407),
.B3(n_410),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_534),
.B(n_537),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_547),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_551),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_534),
.B(n_517),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_537),
.B(n_517),
.Y(n_693)
);

A2O1A1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_571),
.A2(n_432),
.B(n_446),
.C(n_401),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_602),
.B(n_352),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_556),
.A2(n_517),
.B1(n_203),
.B2(n_237),
.Y(n_696)
);

CKINVDCx16_ASAP7_75t_R g697 ( 
.A(n_526),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_551),
.A2(n_388),
.B(n_387),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_599),
.A2(n_478),
.B(n_446),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_535),
.Y(n_700)
);

NOR3xp33_ASAP7_75t_L g701 ( 
.A(n_586),
.B(n_432),
.C(n_446),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_544),
.B(n_296),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_563),
.B(n_337),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_524),
.A2(n_270),
.B1(n_286),
.B2(n_271),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_542),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_607),
.A2(n_557),
.B(n_618),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_618),
.A2(n_478),
.B(n_397),
.Y(n_707)
);

AOI21x1_ASAP7_75t_L g708 ( 
.A1(n_562),
.A2(n_388),
.B(n_387),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_620),
.A2(n_531),
.B(n_592),
.C(n_564),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_526),
.B(n_535),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_577),
.A2(n_395),
.B(n_399),
.C(n_403),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_R g712 ( 
.A(n_592),
.B(n_275),
.Y(n_712)
);

INVxp67_ASAP7_75t_R g713 ( 
.A(n_561),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_542),
.B(n_395),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_562),
.A2(n_400),
.B(n_399),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_612),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_SL g717 ( 
.A(n_644),
.B(n_539),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_639),
.B(n_584),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_659),
.B(n_603),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_630),
.B(n_564),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_689),
.A2(n_260),
.B1(n_248),
.B2(n_613),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_642),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_645),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_661),
.A2(n_650),
.B(n_656),
.Y(n_724)
);

O2A1O1Ixp33_ASAP7_75t_SL g725 ( 
.A1(n_709),
.A2(n_616),
.B(n_609),
.C(n_575),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_623),
.B(n_569),
.Y(n_726)
);

A2O1A1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_679),
.A2(n_585),
.B(n_569),
.C(n_575),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_SL g728 ( 
.A(n_625),
.B(n_260),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_634),
.B(n_588),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_648),
.A2(n_612),
.B1(n_613),
.B2(n_585),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_697),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_658),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_667),
.B(n_581),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_661),
.A2(n_580),
.B(n_576),
.Y(n_734)
);

O2A1O1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_621),
.A2(n_580),
.B(n_576),
.C(n_583),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_695),
.B(n_581),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_705),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_652),
.A2(n_583),
.B(n_588),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_631),
.B(n_587),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_646),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_633),
.B(n_587),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_654),
.A2(n_588),
.B(n_589),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_622),
.B(n_588),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_680),
.A2(n_588),
.B(n_589),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_649),
.A2(n_588),
.B(n_600),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_671),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_635),
.B(n_600),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_639),
.B(n_606),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_641),
.Y(n_749)
);

AO32x1_ASAP7_75t_L g750 ( 
.A1(n_682),
.A2(n_606),
.A3(n_614),
.B1(n_615),
.B2(n_601),
.Y(n_750)
);

INVx5_ASAP7_75t_L g751 ( 
.A(n_663),
.Y(n_751)
);

OAI21x1_ASAP7_75t_L g752 ( 
.A1(n_677),
.A2(n_582),
.B(n_566),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_664),
.A2(n_615),
.B(n_614),
.C(n_601),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_686),
.B(n_588),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_641),
.B(n_596),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_637),
.A2(n_596),
.B(n_595),
.C(n_582),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_688),
.B(n_595),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_712),
.Y(n_758)
);

O2A1O1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_665),
.A2(n_566),
.B(n_403),
.C(n_400),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_690),
.B(n_394),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_668),
.B(n_337),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_691),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_624),
.A2(n_478),
.B(n_209),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_678),
.B(n_394),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_672),
.A2(n_275),
.B(n_276),
.C(n_315),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_704),
.A2(n_337),
.B1(n_276),
.B2(n_407),
.Y(n_766)
);

O2A1O1Ixp5_ASAP7_75t_SL g767 ( 
.A1(n_653),
.A2(n_410),
.B(n_384),
.C(n_255),
.Y(n_767)
);

OA21x2_ASAP7_75t_L g768 ( 
.A1(n_653),
.A2(n_397),
.B(n_233),
.Y(n_768)
);

O2A1O1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_662),
.A2(n_397),
.B(n_384),
.C(n_4),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_701),
.B(n_205),
.Y(n_770)
);

O2A1O1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_694),
.A2(n_384),
.B(n_3),
.C(n_6),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_683),
.Y(n_772)
);

BUFx12f_ASAP7_75t_L g773 ( 
.A(n_702),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_657),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_687),
.B(n_211),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_716),
.B(n_385),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_626),
.A2(n_647),
.B(n_628),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_716),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_676),
.A2(n_478),
.B(n_244),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_666),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_676),
.A2(n_478),
.B(n_227),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_734),
.A2(n_676),
.B(n_710),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_735),
.A2(n_706),
.B(n_632),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_719),
.B(n_674),
.Y(n_784)
);

OAI22x1_ASAP7_75t_L g785 ( 
.A1(n_718),
.A2(n_703),
.B1(n_704),
.B2(n_673),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_SL g786 ( 
.A1(n_720),
.A2(n_700),
.B(n_663),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_722),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_762),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_SL g789 ( 
.A(n_728),
.B(n_625),
.C(n_675),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_752),
.A2(n_655),
.B(n_627),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_736),
.B(n_716),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_724),
.A2(n_676),
.B(n_670),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_723),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_777),
.A2(n_669),
.B(n_660),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_731),
.Y(n_795)
);

AND3x4_ASAP7_75t_L g796 ( 
.A(n_718),
.B(n_713),
.C(n_711),
.Y(n_796)
);

BUFx5_ASAP7_75t_L g797 ( 
.A(n_776),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_738),
.A2(n_693),
.B(n_692),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_717),
.A2(n_629),
.B(n_699),
.C(n_684),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_720),
.B(n_714),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_725),
.A2(n_638),
.B(n_636),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_L g802 ( 
.A(n_761),
.B(n_696),
.C(n_715),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_726),
.A2(n_643),
.B(n_681),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_721),
.A2(n_715),
.B(n_714),
.C(n_698),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_744),
.A2(n_742),
.B(n_739),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_745),
.A2(n_708),
.B(n_698),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_733),
.B(n_663),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_741),
.A2(n_651),
.B(n_700),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_767),
.A2(n_707),
.B(n_685),
.Y(n_809)
);

AOI211x1_ASAP7_75t_L g810 ( 
.A1(n_721),
.A2(n_2),
.B(n_3),
.C(n_6),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_741),
.A2(n_700),
.B(n_478),
.Y(n_811)
);

BUFx10_ASAP7_75t_L g812 ( 
.A(n_772),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_771),
.A2(n_640),
.B(n_246),
.C(n_225),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_748),
.B(n_212),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_740),
.A2(n_251),
.B1(n_214),
.B2(n_215),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_749),
.B(n_53),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_780),
.Y(n_817)
);

OAI21x1_ASAP7_75t_L g818 ( 
.A1(n_764),
.A2(n_384),
.B(n_385),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_753),
.A2(n_261),
.B(n_216),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_758),
.B(n_213),
.Y(n_820)
);

AO31x2_ASAP7_75t_L g821 ( 
.A1(n_727),
.A2(n_2),
.A3(n_8),
.B(n_9),
.Y(n_821)
);

AOI221x1_ASAP7_75t_L g822 ( 
.A1(n_765),
.A2(n_385),
.B1(n_391),
.B2(n_389),
.C(n_15),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_764),
.A2(n_265),
.B(n_221),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_769),
.A2(n_219),
.B(n_385),
.C(n_389),
.Y(n_824)
);

OA22x2_ASAP7_75t_L g825 ( 
.A1(n_766),
.A2(n_748),
.B1(n_774),
.B2(n_754),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_760),
.A2(n_385),
.B(n_91),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_760),
.A2(n_385),
.B(n_89),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_773),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_778),
.B(n_54),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_778),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_746),
.B(n_55),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_756),
.A2(n_391),
.B(n_389),
.Y(n_832)
);

NAND2x1_ASAP7_75t_L g833 ( 
.A(n_776),
.B(n_391),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_751),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_SL g835 ( 
.A1(n_729),
.A2(n_94),
.B(n_169),
.C(n_167),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_766),
.B(n_9),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_789),
.A2(n_770),
.B1(n_743),
.B2(n_755),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_793),
.Y(n_838)
);

BUFx12f_ASAP7_75t_L g839 ( 
.A(n_812),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_790),
.Y(n_840)
);

BUFx4f_ASAP7_75t_SL g841 ( 
.A(n_812),
.Y(n_841)
);

BUFx8_ASAP7_75t_L g842 ( 
.A(n_828),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_826),
.Y(n_843)
);

OAI22xp33_ASAP7_75t_L g844 ( 
.A1(n_784),
.A2(n_775),
.B1(n_747),
.B2(n_757),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_818),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_834),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_796),
.A2(n_747),
.B1(n_730),
.B2(n_732),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_806),
.Y(n_848)
);

INVx5_ASAP7_75t_L g849 ( 
.A(n_831),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_836),
.A2(n_737),
.B1(n_768),
.B2(n_730),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_SL g851 ( 
.A1(n_802),
.A2(n_768),
.B1(n_751),
.B2(n_776),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_791),
.B(n_751),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_821),
.Y(n_853)
);

BUFx12f_ASAP7_75t_L g854 ( 
.A(n_830),
.Y(n_854)
);

BUFx12f_ASAP7_75t_L g855 ( 
.A(n_829),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_795),
.Y(n_856)
);

NAND2x1p5_ASAP7_75t_L g857 ( 
.A(n_827),
.B(n_751),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_821),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_795),
.Y(n_859)
);

INVx6_ASAP7_75t_L g860 ( 
.A(n_829),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_821),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_SL g862 ( 
.A1(n_785),
.A2(n_776),
.B1(n_763),
.B2(n_15),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_825),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_831),
.B(n_776),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_825),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_817),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_802),
.A2(n_759),
.B1(n_779),
.B2(n_781),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_788),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_807),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_823),
.A2(n_391),
.B1(n_750),
.B2(n_16),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_833),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_797),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_800),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_797),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_823),
.B(n_56),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_797),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_804),
.Y(n_877)
);

BUFx8_ASAP7_75t_L g878 ( 
.A(n_797),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_819),
.A2(n_391),
.B1(n_750),
.B2(n_18),
.Y(n_879)
);

OAI22xp33_ASAP7_75t_L g880 ( 
.A1(n_822),
.A2(n_391),
.B1(n_13),
.B2(n_19),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_816),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_SL g882 ( 
.A1(n_810),
.A2(n_11),
.B1(n_13),
.B2(n_20),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_797),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_808),
.Y(n_884)
);

AO22x1_ASAP7_75t_L g885 ( 
.A1(n_787),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_885)
);

CKINVDCx11_ASAP7_75t_R g886 ( 
.A(n_816),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_783),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_819),
.A2(n_750),
.B1(n_24),
.B2(n_25),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_820),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_814),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_786),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_805),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_832),
.Y(n_893)
);

INVx5_ASAP7_75t_L g894 ( 
.A(n_835),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_857),
.A2(n_794),
.B(n_792),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_848),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_861),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_853),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_843),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_848),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_863),
.B(n_782),
.Y(n_901)
);

CKINVDCx9p33_ASAP7_75t_R g902 ( 
.A(n_887),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_861),
.B(n_809),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_853),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_858),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_848),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_858),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_892),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_861),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_892),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_840),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_866),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_866),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_866),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_840),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_863),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_865),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_884),
.Y(n_918)
);

OAI21x1_ASAP7_75t_L g919 ( 
.A1(n_857),
.A2(n_798),
.B(n_801),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_840),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_SL g921 ( 
.A1(n_880),
.A2(n_824),
.B(n_813),
.C(n_799),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_840),
.Y(n_922)
);

NAND4xp25_ASAP7_75t_L g923 ( 
.A(n_862),
.B(n_815),
.C(n_803),
.D(n_809),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_865),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_877),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_840),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_877),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_887),
.B(n_832),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_840),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_884),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_838),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_843),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_928),
.B(n_838),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_899),
.Y(n_934)
);

AO32x2_ASAP7_75t_L g935 ( 
.A1(n_929),
.A2(n_882),
.A3(n_847),
.B1(n_869),
.B2(n_856),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_923),
.A2(n_882),
.B1(n_875),
.B2(n_890),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_923),
.A2(n_875),
.B1(n_885),
.B2(n_889),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_928),
.A2(n_862),
.B(n_849),
.C(n_881),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_898),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_928),
.B(n_869),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_901),
.A2(n_849),
.B(n_881),
.C(n_888),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_931),
.B(n_851),
.Y(n_942)
);

NOR2x1_ASAP7_75t_SL g943 ( 
.A(n_925),
.B(n_891),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_931),
.B(n_850),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_925),
.B(n_873),
.Y(n_945)
);

CKINVDCx6p67_ASAP7_75t_R g946 ( 
.A(n_902),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_912),
.B(n_893),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_912),
.Y(n_948)
);

OAI211xp5_ASAP7_75t_L g949 ( 
.A1(n_921),
.A2(n_886),
.B(n_879),
.C(n_870),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_913),
.B(n_893),
.Y(n_950)
);

AO32x1_ASAP7_75t_L g951 ( 
.A1(n_898),
.A2(n_845),
.A3(n_893),
.B1(n_867),
.B2(n_872),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_916),
.A2(n_859),
.B1(n_849),
.B2(n_881),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_916),
.B(n_854),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_904),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_913),
.Y(n_955)
);

OA21x2_ASAP7_75t_L g956 ( 
.A1(n_919),
.A2(n_845),
.B(n_837),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_914),
.B(n_872),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_914),
.B(n_872),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_901),
.A2(n_849),
.B(n_864),
.C(n_894),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_917),
.B(n_876),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_917),
.B(n_876),
.Y(n_961)
);

OAI21xp33_ASAP7_75t_SL g962 ( 
.A1(n_927),
.A2(n_873),
.B(n_891),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_924),
.A2(n_849),
.B1(n_860),
.B2(n_856),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_921),
.A2(n_844),
.B(n_852),
.C(n_891),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_899),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_924),
.B(n_854),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_901),
.A2(n_885),
.B1(n_855),
.B2(n_860),
.Y(n_967)
);

NAND3xp33_ASAP7_75t_L g968 ( 
.A(n_901),
.B(n_927),
.C(n_918),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_930),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_901),
.A2(n_849),
.B(n_864),
.C(n_894),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_969),
.Y(n_971)
);

INVxp67_ASAP7_75t_SL g972 ( 
.A(n_968),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_933),
.B(n_920),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_933),
.B(n_920),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_934),
.B(n_920),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_934),
.B(n_920),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_934),
.B(n_922),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_944),
.B(n_918),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_965),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_968),
.B(n_897),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_944),
.B(n_930),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_939),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_940),
.B(n_930),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_969),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_965),
.B(n_922),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_939),
.Y(n_986)
);

NAND2xp33_ASAP7_75t_L g987 ( 
.A(n_936),
.B(n_864),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_965),
.B(n_922),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_965),
.B(n_922),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_954),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_946),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_954),
.B(n_897),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_948),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_948),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_955),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_978),
.B(n_940),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_971),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_978),
.B(n_981),
.Y(n_998)
);

OA21x2_ASAP7_75t_L g999 ( 
.A1(n_972),
.A2(n_980),
.B(n_982),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_973),
.B(n_965),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_994),
.Y(n_1001)
);

OAI31xp33_ASAP7_75t_SL g1002 ( 
.A1(n_972),
.A2(n_949),
.A3(n_942),
.B(n_952),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_973),
.B(n_956),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_981),
.B(n_960),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_979),
.B(n_985),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_991),
.B(n_937),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_983),
.B(n_955),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_973),
.B(n_943),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_991),
.B(n_953),
.Y(n_1009)
);

AND2x4_ASAP7_75t_SL g1010 ( 
.A(n_991),
.B(n_946),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_979),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_974),
.B(n_956),
.Y(n_1012)
);

OAI33xp33_ASAP7_75t_L g1013 ( 
.A1(n_982),
.A2(n_945),
.A3(n_905),
.B1(n_907),
.B2(n_904),
.B3(n_964),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_974),
.B(n_956),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_974),
.B(n_943),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_983),
.B(n_903),
.Y(n_1016)
);

NAND4xp25_ASAP7_75t_L g1017 ( 
.A(n_1002),
.B(n_937),
.C(n_936),
.D(n_966),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_1005),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1001),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1008),
.B(n_985),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_997),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1008),
.B(n_985),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1015),
.B(n_988),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_1011),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_1015),
.B(n_988),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_998),
.B(n_980),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_998),
.B(n_980),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1018),
.B(n_1005),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1019),
.Y(n_1029)
);

AO31x2_ASAP7_75t_L g1030 ( 
.A1(n_1021),
.A2(n_991),
.A3(n_1009),
.B(n_997),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1021),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_1017),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_1024),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1020),
.B(n_1005),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1034),
.B(n_1020),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_1032),
.B(n_839),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_1029),
.B(n_841),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1029),
.Y(n_1038)
);

OAI211xp5_ASAP7_75t_L g1039 ( 
.A1(n_1036),
.A2(n_1002),
.B(n_1006),
.C(n_1033),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1038),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1036),
.B(n_1028),
.Y(n_1041)
);

AOI32xp33_ASAP7_75t_L g1042 ( 
.A1(n_1035),
.A2(n_987),
.A3(n_1028),
.B1(n_1033),
.B2(n_1010),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1037),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1035),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1036),
.A2(n_987),
.B(n_938),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1038),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1038),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1036),
.B(n_1034),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_1036),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_1039),
.A2(n_1041),
.B(n_1048),
.Y(n_1050)
);

AOI21xp33_ASAP7_75t_SL g1051 ( 
.A1(n_1049),
.A2(n_999),
.B(n_1024),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1040),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_1043),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_1049),
.B(n_839),
.Y(n_1054)
);

NAND2x1p5_ASAP7_75t_L g1055 ( 
.A(n_1046),
.B(n_991),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1044),
.B(n_1026),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1044),
.B(n_1026),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_1047),
.B(n_1027),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1045),
.A2(n_1010),
.B1(n_1027),
.B2(n_999),
.Y(n_1059)
);

OAI21xp33_ASAP7_75t_SL g1060 ( 
.A1(n_1042),
.A2(n_1031),
.B(n_1023),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1049),
.B(n_1022),
.Y(n_1061)
);

OAI221xp5_ASAP7_75t_SL g1062 ( 
.A1(n_1039),
.A2(n_967),
.B1(n_941),
.B2(n_1031),
.C(n_959),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_1039),
.A2(n_999),
.B(n_1013),
.C(n_1011),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_1039),
.A2(n_999),
.B(n_1013),
.C(n_1011),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_1044),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1065),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1050),
.B(n_1022),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1053),
.B(n_1023),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_1061),
.B(n_996),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_1052),
.B(n_1030),
.Y(n_1070)
);

OAI221xp5_ASAP7_75t_L g1071 ( 
.A1(n_1062),
.A2(n_967),
.B1(n_999),
.B2(n_970),
.C(n_996),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1054),
.B(n_1025),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1057),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_1058),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1056),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1055),
.B(n_1025),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1055),
.B(n_1030),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1060),
.B(n_1030),
.Y(n_1078)
);

XOR2x2_ASAP7_75t_L g1079 ( 
.A(n_1059),
.B(n_839),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1063),
.A2(n_1010),
.B1(n_842),
.B2(n_855),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1064),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_1051),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1050),
.B(n_1030),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_1065),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1084),
.B(n_1030),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_L g1086 ( 
.A(n_1066),
.B(n_842),
.C(n_846),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1074),
.B(n_1000),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1073),
.B(n_1001),
.Y(n_1088)
);

AOI21x1_ASAP7_75t_L g1089 ( 
.A1(n_1081),
.A2(n_1005),
.B(n_997),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1082),
.A2(n_1004),
.B(n_951),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1075),
.B(n_1000),
.Y(n_1091)
);

OAI32xp33_ASAP7_75t_L g1092 ( 
.A1(n_1083),
.A2(n_1003),
.A3(n_1014),
.B1(n_1012),
.B2(n_1016),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1068),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_L g1094 ( 
.A(n_1067),
.B(n_842),
.C(n_846),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1069),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_L g1096 ( 
.A(n_1072),
.B(n_1078),
.C(n_1076),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1077),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1080),
.A2(n_962),
.B(n_22),
.Y(n_1098)
);

NAND3xp33_ASAP7_75t_SL g1099 ( 
.A(n_1080),
.B(n_842),
.C(n_963),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_1079),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_SL g1101 ( 
.A(n_1071),
.B(n_1012),
.C(n_1003),
.Y(n_1101)
);

OAI21xp33_ASAP7_75t_L g1102 ( 
.A1(n_1087),
.A2(n_1070),
.B(n_1012),
.Y(n_1102)
);

NAND4xp75_ASAP7_75t_L g1103 ( 
.A(n_1093),
.B(n_1070),
.C(n_979),
.D(n_30),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_1095),
.B(n_1007),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1096),
.B(n_1003),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1100),
.A2(n_1004),
.B(n_951),
.Y(n_1106)
);

NAND4xp25_ASAP7_75t_L g1107 ( 
.A(n_1086),
.B(n_1094),
.C(n_1088),
.D(n_1091),
.Y(n_1107)
);

AOI211x1_ASAP7_75t_SL g1108 ( 
.A1(n_1101),
.A2(n_1098),
.B(n_1099),
.C(n_1085),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1097),
.B(n_1014),
.Y(n_1109)
);

AOI221xp5_ASAP7_75t_L g1110 ( 
.A1(n_1098),
.A2(n_1014),
.B1(n_942),
.B2(n_962),
.C(n_995),
.Y(n_1110)
);

NOR2x1_ASAP7_75t_R g1111 ( 
.A(n_1089),
.B(n_846),
.Y(n_1111)
);

AOI211xp5_ASAP7_75t_L g1112 ( 
.A1(n_1092),
.A2(n_26),
.B(n_27),
.C(n_30),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_R g1113 ( 
.A(n_1090),
.B(n_32),
.Y(n_1113)
);

AO221x1_ASAP7_75t_L g1114 ( 
.A1(n_1093),
.A2(n_899),
.B1(n_990),
.B2(n_986),
.C(n_871),
.Y(n_1114)
);

AOI221xp5_ASAP7_75t_L g1115 ( 
.A1(n_1096),
.A2(n_995),
.B1(n_993),
.B2(n_990),
.C(n_986),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_L g1116 ( 
.A(n_1100),
.B(n_868),
.C(n_1016),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1100),
.A2(n_1007),
.B1(n_993),
.B2(n_860),
.Y(n_1117)
);

NOR3x1_ASAP7_75t_L g1118 ( 
.A(n_1093),
.B(n_32),
.C(n_33),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1098),
.A2(n_932),
.B(n_34),
.C(n_35),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1100),
.A2(n_951),
.B(n_868),
.Y(n_1120)
);

AOI221xp5_ASAP7_75t_L g1121 ( 
.A1(n_1096),
.A2(n_994),
.B1(n_977),
.B2(n_976),
.C(n_975),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1095),
.B(n_33),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1087),
.B(n_35),
.Y(n_1123)
);

AOI221xp5_ASAP7_75t_L g1124 ( 
.A1(n_1096),
.A2(n_975),
.B1(n_976),
.B2(n_977),
.C(n_989),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_L g1125 ( 
.A(n_1100),
.B(n_868),
.C(n_894),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1118),
.B(n_36),
.Y(n_1126)
);

AOI222xp33_ASAP7_75t_L g1127 ( 
.A1(n_1115),
.A2(n_894),
.B1(n_39),
.B2(n_40),
.C1(n_41),
.C2(n_42),
.Y(n_1127)
);

OAI211xp5_ASAP7_75t_L g1128 ( 
.A1(n_1112),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1122),
.Y(n_1129)
);

AOI221xp5_ASAP7_75t_L g1130 ( 
.A1(n_1107),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.C(n_44),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1116),
.A2(n_860),
.B1(n_989),
.B2(n_988),
.Y(n_1131)
);

OAI21xp33_ASAP7_75t_SL g1132 ( 
.A1(n_1103),
.A2(n_989),
.B(n_975),
.Y(n_1132)
);

OAI222xp33_ASAP7_75t_R g1133 ( 
.A1(n_1108),
.A2(n_43),
.B1(n_46),
.B2(n_49),
.C1(n_50),
.C2(n_51),
.Y(n_1133)
);

NOR3xp33_ASAP7_75t_SL g1134 ( 
.A(n_1123),
.B(n_49),
.C(n_52),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1119),
.A2(n_864),
.B(n_895),
.Y(n_1135)
);

OAI221xp5_ASAP7_75t_L g1136 ( 
.A1(n_1121),
.A2(n_894),
.B1(n_932),
.B2(n_857),
.C(n_971),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1124),
.A2(n_1105),
.B1(n_1113),
.B2(n_1110),
.Y(n_1137)
);

AOI311xp33_ASAP7_75t_L g1138 ( 
.A1(n_1117),
.A2(n_905),
.A3(n_907),
.B(n_909),
.C(n_935),
.Y(n_1138)
);

AOI211xp5_ASAP7_75t_L g1139 ( 
.A1(n_1111),
.A2(n_977),
.B(n_976),
.C(n_899),
.Y(n_1139)
);

OAI211xp5_ASAP7_75t_L g1140 ( 
.A1(n_1102),
.A2(n_894),
.B(n_811),
.C(n_971),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1125),
.B(n_1109),
.C(n_1104),
.Y(n_1141)
);

OAI211xp5_ASAP7_75t_SL g1142 ( 
.A1(n_1106),
.A2(n_932),
.B(n_984),
.C(n_971),
.Y(n_1142)
);

NOR2x1_ASAP7_75t_L g1143 ( 
.A(n_1120),
.B(n_992),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_1114),
.Y(n_1144)
);

OA21x2_ASAP7_75t_L g1145 ( 
.A1(n_1103),
.A2(n_984),
.B(n_895),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1122),
.Y(n_1146)
);

AOI221xp5_ASAP7_75t_L g1147 ( 
.A1(n_1107),
.A2(n_984),
.B1(n_899),
.B2(n_843),
.C(n_926),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_SL g1148 ( 
.A1(n_1123),
.A2(n_902),
.B(n_935),
.Y(n_1148)
);

AOI221xp5_ASAP7_75t_L g1149 ( 
.A1(n_1107),
.A2(n_899),
.B1(n_843),
.B2(n_926),
.C(n_911),
.Y(n_1149)
);

INVxp33_ASAP7_75t_SL g1150 ( 
.A(n_1126),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1129),
.Y(n_1151)
);

NOR2xp67_ASAP7_75t_L g1152 ( 
.A(n_1128),
.B(n_59),
.Y(n_1152)
);

NOR2x1_ASAP7_75t_L g1153 ( 
.A(n_1146),
.B(n_992),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1132),
.A2(n_929),
.B1(n_899),
.B2(n_878),
.Y(n_1154)
);

OAI211xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1137),
.A2(n_926),
.B(n_915),
.C(n_911),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1134),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1141),
.B(n_62),
.Y(n_1157)
);

NOR2x1_ASAP7_75t_L g1158 ( 
.A(n_1144),
.B(n_1145),
.Y(n_1158)
);

NAND4xp75_ASAP7_75t_L g1159 ( 
.A(n_1130),
.B(n_956),
.C(n_929),
.D(n_961),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_L g1160 ( 
.A(n_1127),
.B(n_1133),
.C(n_1147),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1135),
.B(n_992),
.Y(n_1161)
);

NAND2x1p5_ASAP7_75t_L g1162 ( 
.A(n_1145),
.B(n_871),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1140),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1143),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1148),
.Y(n_1165)
);

NAND4xp75_ASAP7_75t_L g1166 ( 
.A(n_1149),
.B(n_961),
.C(n_960),
.D(n_958),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1142),
.Y(n_1167)
);

NOR2x1_ASAP7_75t_L g1168 ( 
.A(n_1136),
.B(n_63),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1131),
.B(n_64),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1139),
.A2(n_1138),
.B1(n_926),
.B2(n_911),
.Y(n_1170)
);

NOR2x1_ASAP7_75t_L g1171 ( 
.A(n_1126),
.B(n_65),
.Y(n_1171)
);

NAND4xp75_ASAP7_75t_L g1172 ( 
.A(n_1158),
.B(n_69),
.C(n_71),
.D(n_72),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_SL g1173 ( 
.A(n_1156),
.B(n_935),
.C(n_878),
.Y(n_1173)
);

AOI211xp5_ASAP7_75t_L g1174 ( 
.A1(n_1164),
.A2(n_899),
.B(n_843),
.C(n_871),
.Y(n_1174)
);

OAI211xp5_ASAP7_75t_SL g1175 ( 
.A1(n_1151),
.A2(n_74),
.B(n_75),
.C(n_76),
.Y(n_1175)
);

NAND4xp25_ASAP7_75t_L g1176 ( 
.A(n_1160),
.B(n_910),
.C(n_908),
.D(n_903),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1167),
.B(n_957),
.Y(n_1177)
);

NAND3x1_ASAP7_75t_L g1178 ( 
.A(n_1171),
.B(n_935),
.C(n_874),
.Y(n_1178)
);

NOR2x1p5_ASAP7_75t_L g1179 ( 
.A(n_1165),
.B(n_871),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_1157),
.B(n_878),
.C(n_843),
.Y(n_1180)
);

NAND4xp25_ASAP7_75t_L g1181 ( 
.A(n_1150),
.B(n_910),
.C(n_908),
.D(n_903),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1152),
.A2(n_951),
.B(n_895),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1153),
.Y(n_1183)
);

NOR3xp33_ASAP7_75t_L g1184 ( 
.A(n_1169),
.B(n_915),
.C(n_84),
.Y(n_1184)
);

AOI221xp5_ASAP7_75t_L g1185 ( 
.A1(n_1163),
.A2(n_915),
.B1(n_958),
.B2(n_957),
.C(n_908),
.Y(n_1185)
);

NOR2x1_ASAP7_75t_L g1186 ( 
.A(n_1168),
.B(n_81),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1183),
.A2(n_1154),
.B(n_1162),
.Y(n_1187)
);

AO22x2_ASAP7_75t_L g1188 ( 
.A1(n_1172),
.A2(n_1159),
.B1(n_1166),
.B2(n_1170),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1179),
.Y(n_1189)
);

NAND4xp25_ASAP7_75t_L g1190 ( 
.A(n_1186),
.B(n_1155),
.C(n_1161),
.D(n_97),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1177),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1184),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1180),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_SL g1194 ( 
.A1(n_1174),
.A2(n_1161),
.B1(n_935),
.B2(n_871),
.Y(n_1194)
);

AND3x1_ASAP7_75t_L g1195 ( 
.A(n_1185),
.B(n_1182),
.C(n_1175),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1176),
.A2(n_910),
.B(n_909),
.C(n_935),
.Y(n_1196)
);

NOR3x1_ASAP7_75t_L g1197 ( 
.A(n_1173),
.B(n_88),
.C(n_95),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1181),
.B(n_950),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1178),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1183),
.A2(n_951),
.B(n_883),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1183),
.Y(n_1201)
);

AO22x2_ASAP7_75t_L g1202 ( 
.A1(n_1201),
.A2(n_874),
.B1(n_906),
.B2(n_900),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1193),
.A2(n_878),
.B1(n_871),
.B2(n_874),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1199),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1199),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1188),
.A2(n_950),
.B1(n_947),
.B2(n_897),
.Y(n_1206)
);

OAI22x1_ASAP7_75t_L g1207 ( 
.A1(n_1191),
.A2(n_874),
.B1(n_101),
.B2(n_103),
.Y(n_1207)
);

AO22x2_ASAP7_75t_L g1208 ( 
.A1(n_1189),
.A2(n_906),
.B1(n_900),
.B2(n_896),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1197),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_SL g1210 ( 
.A1(n_1192),
.A2(n_1195),
.B1(n_1194),
.B2(n_1187),
.Y(n_1210)
);

INVxp67_ASAP7_75t_SL g1211 ( 
.A(n_1190),
.Y(n_1211)
);

AO22x2_ASAP7_75t_L g1212 ( 
.A1(n_1204),
.A2(n_1198),
.B1(n_1200),
.B2(n_1196),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1205),
.Y(n_1213)
);

XNOR2x1_ASAP7_75t_L g1214 ( 
.A(n_1209),
.B(n_98),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1210),
.A2(n_106),
.B(n_107),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1211),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1207),
.B(n_113),
.Y(n_1217)
);

XOR2x2_ASAP7_75t_L g1218 ( 
.A(n_1214),
.B(n_1203),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1213),
.A2(n_1206),
.B1(n_1202),
.B2(n_1208),
.Y(n_1219)
);

OAI22x1_ASAP7_75t_L g1220 ( 
.A1(n_1217),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1215),
.A2(n_906),
.B1(n_900),
.B2(n_896),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1219),
.A2(n_1216),
.B(n_1212),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1222),
.A2(n_1218),
.B(n_1220),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1223),
.A2(n_1221),
.B(n_126),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1224),
.Y(n_1225)
);

OAI221xp5_ASAP7_75t_R g1226 ( 
.A1(n_1225),
.A2(n_119),
.B1(n_130),
.B2(n_132),
.C(n_134),
.Y(n_1226)
);

AOI211xp5_ASAP7_75t_L g1227 ( 
.A1(n_1226),
.A2(n_135),
.B(n_136),
.C(n_137),
.Y(n_1227)
);


endmodule