module fake_netlist_6_191_n_1624 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1624);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1624;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_52),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_44),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_102),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_21),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_1),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_98),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_55),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_99),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_40),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_47),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_104),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_66),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_5),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_24),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_29),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_105),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_56),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_10),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_60),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_97),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_35),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_61),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_48),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_51),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_140),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_8),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_49),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_124),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_75),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_86),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_4),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_113),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_2),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_76),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_28),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_57),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_41),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_36),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_12),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_36),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_112),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_45),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_21),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_0),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_62),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_42),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_28),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_42),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_50),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_26),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_148),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_5),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_46),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_109),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_131),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_92),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_54),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_2),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_96),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_1),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_107),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_145),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_38),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_77),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_71),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_27),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_18),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_137),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_43),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_119),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_18),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_115),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_93),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_35),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_22),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_37),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_111),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_12),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_144),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_40),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_30),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_69),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_39),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_110),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_0),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_83),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_129),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_128),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_80),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_30),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_58),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_17),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_41),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_143),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_136),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_142),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_103),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_106),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_38),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_64),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_39),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_90),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_120),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_89),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_72),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_134),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_122),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_147),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_33),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_130),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_59),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_13),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_88),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_63),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_82),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_85),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_9),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_14),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_67),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_91),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_65),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_95),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_19),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_13),
.Y(n_283)
);

HB1xp67_ASAP7_75t_SL g284 ( 
.A(n_29),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_4),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_19),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_87),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_138),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_6),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_74),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_15),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_123),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_43),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_94),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_26),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_81),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_179),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_196),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_163),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_196),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_191),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_296),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_177),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_179),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_196),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_155),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_284),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_196),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_275),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_155),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_280),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_196),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_168),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_206),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_206),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_219),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_176),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_214),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_178),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_197),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_160),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_219),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_182),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_185),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_280),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_187),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_240),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_240),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_214),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_276),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_170),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_268),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_184),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_273),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_205),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_200),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_209),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_217),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_213),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_188),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_225),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_228),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_233),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_234),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_190),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_237),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_238),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_244),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_214),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_249),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_251),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_260),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_276),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_151),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_192),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_195),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_277),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_282),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_285),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_289),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_250),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_212),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_276),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_202),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_218),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_220),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_298),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_298),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_318),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_329),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

NOR2x1_ASAP7_75t_L g376 ( 
.A(n_334),
.B(n_269),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_304),
.B(n_269),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_302),
.B(n_164),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_300),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_317),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_335),
.B(n_269),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_300),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_350),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_305),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_319),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_350),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_323),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_311),
.B(n_164),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_313),
.B(n_204),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_308),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_312),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_312),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_334),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_325),
.B(n_204),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_336),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_336),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_314),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_299),
.B(n_180),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_355),
.B(n_184),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_355),
.B(n_149),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_314),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_306),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_338),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_315),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_315),
.A2(n_208),
.B(n_158),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_297),
.B(n_208),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_316),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_339),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_316),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_310),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_301),
.B(n_202),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_321),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_297),
.B(n_153),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_331),
.A2(n_295),
.B1(n_154),
.B2(n_203),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_342),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_322),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_322),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_324),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_327),
.B(n_157),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_327),
.B(n_167),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_328),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_303),
.B(n_215),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_328),
.B(n_175),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_332),
.B(n_181),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_332),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_333),
.B(n_186),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_342),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_333),
.B(n_194),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_402),
.B(n_309),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_402),
.B(n_335),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_370),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_377),
.B(n_366),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_370),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_392),
.B(n_326),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_370),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_373),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_396),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_396),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_398),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_377),
.B(n_341),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_377),
.B(n_346),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_369),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_371),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_427),
.B(n_392),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_372),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_427),
.B(n_356),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_372),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_380),
.B(n_357),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_380),
.B(n_363),
.Y(n_455)
);

OAI22xp33_ASAP7_75t_L g456 ( 
.A1(n_415),
.A2(n_364),
.B1(n_354),
.B2(n_301),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_373),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_373),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_381),
.B(n_367),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_374),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_417),
.B(n_366),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_375),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_375),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

AND3x2_ASAP7_75t_L g466 ( 
.A(n_378),
.B(n_330),
.C(n_210),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_375),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_382),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_396),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_378),
.B(n_368),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_398),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_375),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_417),
.B(n_157),
.Y(n_473)
);

NAND3xp33_ASAP7_75t_L g474 ( 
.A(n_406),
.B(n_364),
.C(n_320),
.Y(n_474)
);

INVxp33_ASAP7_75t_L g475 ( 
.A(n_418),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_410),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_387),
.B(n_354),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_396),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_385),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_R g480 ( 
.A(n_387),
.B(n_337),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_374),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_410),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_374),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_385),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_382),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_385),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_369),
.Y(n_488)
);

BUFx8_ASAP7_75t_SL g489 ( 
.A(n_389),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_374),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_410),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_418),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_381),
.B(n_340),
.Y(n_493)
);

OR2x6_ASAP7_75t_L g494 ( 
.A(n_369),
.B(n_343),
.Y(n_494)
);

NAND3xp33_ASAP7_75t_L g495 ( 
.A(n_406),
.B(n_189),
.C(n_183),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_399),
.Y(n_496)
);

AOI21x1_ASAP7_75t_L g497 ( 
.A1(n_383),
.A2(n_395),
.B(n_386),
.Y(n_497)
);

NAND3xp33_ASAP7_75t_SL g498 ( 
.A(n_415),
.B(n_169),
.C(n_168),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_388),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_417),
.B(n_343),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_389),
.B(n_149),
.Y(n_501)
);

NOR2x1p5_ASAP7_75t_L g502 ( 
.A(n_415),
.B(n_169),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_374),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_383),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_414),
.B(n_348),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_386),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_SL g507 ( 
.A1(n_390),
.A2(n_263),
.B1(n_290),
.B2(n_362),
.Y(n_507)
);

BUFx16f_ASAP7_75t_R g508 ( 
.A(n_416),
.Y(n_508)
);

INVx8_ASAP7_75t_L g509 ( 
.A(n_410),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_388),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_396),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_403),
.B(n_365),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_423),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_423),
.B(n_150),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_410),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_401),
.Y(n_516)
);

INVxp33_ASAP7_75t_L g517 ( 
.A(n_404),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_396),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_388),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_388),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_393),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_396),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_404),
.B(n_150),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_397),
.Y(n_524)
);

INVx5_ASAP7_75t_L g525 ( 
.A(n_391),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_396),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_393),
.Y(n_527)
);

BUFx6f_ASAP7_75t_SL g528 ( 
.A(n_410),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_403),
.B(n_266),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_393),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_395),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_409),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_391),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_409),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_425),
.B(n_365),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_391),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_409),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_393),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_401),
.Y(n_539)
);

AOI21x1_ASAP7_75t_L g540 ( 
.A1(n_376),
.A2(n_278),
.B(n_201),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_405),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_414),
.B(n_152),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_403),
.B(n_221),
.Y(n_543)
);

CKINVDCx6p67_ASAP7_75t_R g544 ( 
.A(n_416),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_391),
.Y(n_545)
);

AO21x2_ASAP7_75t_L g546 ( 
.A1(n_425),
.A2(n_267),
.B(n_216),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_407),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_424),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_391),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_425),
.B(n_223),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_428),
.A2(n_157),
.B1(n_360),
.B2(n_359),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_405),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_391),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_424),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_428),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_405),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_428),
.Y(n_557)
);

BUFx8_ASAP7_75t_SL g558 ( 
.A(n_429),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_407),
.A2(n_226),
.B1(n_193),
.B2(n_198),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_429),
.B(n_258),
.C(n_239),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_412),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_433),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_391),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_412),
.B(n_152),
.Y(n_564)
);

NOR2x1p5_ASAP7_75t_L g565 ( 
.A(n_419),
.B(n_171),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_391),
.Y(n_566)
);

AND3x1_ASAP7_75t_L g567 ( 
.A(n_419),
.B(n_361),
.C(n_360),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_394),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_429),
.A2(n_173),
.B1(n_294),
.B2(n_172),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_394),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_405),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_394),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_424),
.Y(n_573)
);

BUFx10_ASAP7_75t_L g574 ( 
.A(n_424),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_420),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_384),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_476),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_562),
.B(n_156),
.Y(n_578)
);

O2A1O1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_450),
.A2(n_432),
.B(n_420),
.C(n_431),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_494),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_459),
.B(n_517),
.Y(n_581)
);

A2O1A1Ixp33_ASAP7_75t_L g582 ( 
.A1(n_524),
.A2(n_433),
.B(n_431),
.C(n_231),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_555),
.B(n_424),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_480),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_445),
.A2(n_446),
.B1(n_437),
.B2(n_439),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_555),
.B(n_424),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_476),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_512),
.Y(n_588)
);

NAND3x1_ASAP7_75t_L g589 ( 
.A(n_505),
.B(n_347),
.C(n_344),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_482),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_460),
.B(n_400),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_546),
.A2(n_157),
.B1(n_214),
.B2(n_287),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_470),
.B(n_156),
.Y(n_593)
);

O2A1O1Ixp33_ASAP7_75t_L g594 ( 
.A1(n_557),
.A2(n_432),
.B(n_344),
.C(n_345),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_565),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_548),
.B(n_157),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_548),
.B(n_214),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_546),
.A2(n_214),
.B1(n_246),
.B2(n_236),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_482),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_481),
.B(n_400),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_509),
.B(n_214),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_491),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_452),
.B(n_159),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_448),
.Y(n_604)
);

O2A1O1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_529),
.A2(n_353),
.B(n_345),
.C(n_347),
.Y(n_605)
);

NOR2xp67_ASAP7_75t_L g606 ( 
.A(n_474),
.B(n_400),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_509),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_492),
.A2(n_283),
.B1(n_286),
.B2(n_171),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_535),
.B(n_159),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_512),
.B(n_349),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_448),
.Y(n_611)
);

OAI221xp5_ASAP7_75t_L g612 ( 
.A1(n_551),
.A2(n_259),
.B1(n_256),
.B2(n_241),
.C(n_292),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_491),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_490),
.B(n_394),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_546),
.A2(n_214),
.B1(n_281),
.B2(n_243),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_488),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_515),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_554),
.B(n_394),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_535),
.B(n_161),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_436),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_515),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_500),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_554),
.B(n_411),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_573),
.B(n_411),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_573),
.B(n_411),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_532),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_435),
.B(n_161),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_444),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_535),
.B(n_162),
.Y(n_629)
);

OR2x2_ASAP7_75t_SL g630 ( 
.A(n_498),
.B(n_351),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_456),
.B(n_162),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_471),
.B(n_411),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_509),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_496),
.B(n_411),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_516),
.B(n_411),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_SL g636 ( 
.A(n_559),
.B(n_283),
.C(n_271),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_438),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_440),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_539),
.B(n_411),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_543),
.B(n_165),
.Y(n_640)
);

OAI221xp5_ASAP7_75t_L g641 ( 
.A1(n_569),
.A2(n_351),
.B1(n_361),
.B2(n_359),
.C(n_358),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_547),
.B(n_413),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_574),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_561),
.B(n_413),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_574),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_550),
.A2(n_166),
.B1(n_294),
.B2(n_165),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_575),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_494),
.A2(n_166),
.B1(n_172),
.B2(n_288),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_544),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_447),
.B(n_413),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_434),
.B(n_173),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_532),
.A2(n_174),
.B1(n_291),
.B2(n_286),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_440),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_449),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_449),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_564),
.B(n_270),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_523),
.A2(n_265),
.B1(n_227),
.B2(n_229),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_451),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_500),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_534),
.A2(n_174),
.B1(n_291),
.B2(n_271),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_451),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_572),
.Y(n_662)
);

OAI22xp33_ASAP7_75t_L g663 ( 
.A1(n_475),
.A2(n_199),
.B1(n_211),
.B2(n_222),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_494),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_441),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_493),
.A2(n_528),
.B1(n_560),
.B2(n_502),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_453),
.B(n_413),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_542),
.B(n_270),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_453),
.B(n_413),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_558),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_464),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_528),
.A2(n_461),
.B1(n_514),
.B2(n_501),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_464),
.B(n_413),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_465),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_465),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_441),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_468),
.B(n_413),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_528),
.A2(n_272),
.B1(n_274),
.B2(n_279),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_468),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_544),
.B(n_352),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_485),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_485),
.B(n_413),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_504),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_567),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_495),
.B(n_272),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_572),
.Y(n_686)
);

BUFx5_ASAP7_75t_L g687 ( 
.A(n_537),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_454),
.B(n_274),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_537),
.A2(n_353),
.B1(n_358),
.B2(n_352),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_507),
.B(n_279),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_506),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_473),
.B(n_531),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_461),
.A2(n_254),
.B1(n_224),
.B2(n_232),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_466),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_531),
.B(n_430),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_572),
.B(n_430),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_483),
.B(n_503),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_483),
.B(n_430),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_477),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_455),
.B(n_207),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_457),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_483),
.B(n_430),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_503),
.B(n_426),
.Y(n_703)
);

NOR2x1p5_ASAP7_75t_L g704 ( 
.A(n_513),
.B(n_230),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_503),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_511),
.B(n_426),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_513),
.B(n_288),
.Y(n_707)
);

INVx4_ASAP7_75t_L g708 ( 
.A(n_442),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_511),
.B(n_518),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_497),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_558),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_442),
.B(n_384),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_497),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_511),
.B(n_426),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_442),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_518),
.B(n_426),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_518),
.B(n_422),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_536),
.B(n_422),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_473),
.A2(n_235),
.B1(n_242),
.B2(n_252),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_442),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_458),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_442),
.B(n_384),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_540),
.B(n_422),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_489),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_462),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_536),
.B(n_421),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_462),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_607),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_662),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_607),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_662),
.Y(n_731)
);

NOR2x1p5_ASAP7_75t_L g732 ( 
.A(n_680),
.B(n_508),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_585),
.B(n_463),
.Y(n_733)
);

INVxp67_ASAP7_75t_SL g734 ( 
.A(n_626),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_654),
.B(n_463),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_592),
.A2(n_492),
.B1(n_473),
.B2(n_552),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_655),
.B(n_467),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_686),
.Y(n_738)
);

AND2x6_ASAP7_75t_SL g739 ( 
.A(n_688),
.B(n_489),
.Y(n_739)
);

NOR2x1_ASAP7_75t_R g740 ( 
.A(n_724),
.B(n_245),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_588),
.B(n_540),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_658),
.B(n_661),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_592),
.A2(n_615),
.B1(n_598),
.B2(n_652),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_622),
.B(n_563),
.Y(n_744)
);

INVx6_ASAP7_75t_L g745 ( 
.A(n_610),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_584),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_671),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_649),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_581),
.B(n_533),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_604),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_674),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_SL g752 ( 
.A(n_603),
.B(n_261),
.C(n_248),
.Y(n_752)
);

NOR2x1p5_ASAP7_75t_L g753 ( 
.A(n_700),
.B(n_247),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_643),
.B(n_645),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_686),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_675),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_679),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_659),
.B(n_563),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_607),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_705),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_681),
.B(n_467),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_607),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_683),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_691),
.B(n_472),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_604),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_595),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_626),
.B(n_479),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_633),
.Y(n_768)
);

NOR3xp33_ASAP7_75t_L g769 ( 
.A(n_690),
.B(n_684),
.C(n_707),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_611),
.B(n_533),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_628),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_705),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_611),
.Y(n_773)
);

AO22x1_ASAP7_75t_L g774 ( 
.A1(n_603),
.A2(n_473),
.B1(n_253),
.B2(n_257),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_598),
.A2(n_473),
.B1(n_571),
.B2(n_541),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_590),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_583),
.A2(n_262),
.B1(n_264),
.B2(n_255),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_R g778 ( 
.A(n_699),
.B(n_53),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_670),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_647),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_580),
.Y(n_781)
);

INVx4_ASAP7_75t_L g782 ( 
.A(n_633),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_586),
.B(n_590),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_577),
.A2(n_566),
.B1(n_563),
.B2(n_443),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_672),
.A2(n_526),
.B1(n_469),
.B2(n_522),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_R g786 ( 
.A(n_694),
.B(n_70),
.Y(n_786)
);

NOR2x2_ASAP7_75t_L g787 ( 
.A(n_652),
.B(n_3),
.Y(n_787)
);

XNOR2xp5_ASAP7_75t_SL g788 ( 
.A(n_660),
.B(n_3),
.Y(n_788)
);

AND2x6_ASAP7_75t_SL g789 ( 
.A(n_688),
.B(n_6),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_616),
.B(n_533),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_633),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_587),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_630),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_610),
.Y(n_794)
);

OR2x4_ASAP7_75t_L g795 ( 
.A(n_651),
.B(n_443),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_599),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_616),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_602),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_621),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_580),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_704),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_613),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_617),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_706),
.A2(n_484),
.B(n_519),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_664),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_664),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_651),
.B(n_408),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_685),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_620),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_695),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_606),
.B(n_684),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_643),
.B(n_526),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_579),
.B(n_487),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_615),
.A2(n_660),
.B1(n_612),
.B2(n_713),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_711),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_714),
.A2(n_510),
.B(n_519),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_637),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_627),
.A2(n_566),
.B(n_571),
.C(n_541),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_578),
.Y(n_819)
);

O2A1O1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_582),
.A2(n_556),
.B(n_552),
.C(n_521),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_627),
.B(n_486),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_687),
.B(n_591),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_687),
.B(n_486),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_711),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_609),
.B(n_408),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_687),
.B(n_499),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_666),
.A2(n_566),
.B1(n_469),
.B2(n_478),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_619),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_687),
.B(n_499),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_687),
.B(n_510),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_715),
.Y(n_831)
);

AO22x1_ASAP7_75t_L g832 ( 
.A1(n_668),
.A2(n_556),
.B1(n_568),
.B2(n_570),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_638),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_645),
.B(n_443),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_696),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_600),
.B(n_520),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_715),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_618),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_668),
.B(n_526),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_593),
.A2(n_526),
.B1(n_522),
.B2(n_469),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_608),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_629),
.B(n_478),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_697),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_640),
.A2(n_526),
.B1(n_522),
.B2(n_469),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_633),
.B(n_469),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_636),
.Y(n_846)
);

AND2x2_ASAP7_75t_SL g847 ( 
.A(n_719),
.B(n_522),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_631),
.B(n_408),
.Y(n_848)
);

INVx5_ASAP7_75t_L g849 ( 
.A(n_715),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_R g850 ( 
.A(n_601),
.B(n_100),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_636),
.B(n_478),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_656),
.B(n_553),
.Y(n_852)
);

NOR2x2_ASAP7_75t_L g853 ( 
.A(n_589),
.B(n_7),
.Y(n_853)
);

INVx4_ASAP7_75t_L g854 ( 
.A(n_715),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_693),
.Y(n_855)
);

AND2x6_ASAP7_75t_SL g856 ( 
.A(n_663),
.B(n_8),
.Y(n_856)
);

OAI22xp33_ASAP7_75t_L g857 ( 
.A1(n_641),
.A2(n_663),
.B1(n_710),
.B2(n_614),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_623),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_624),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_646),
.B(n_553),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_653),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_689),
.B(n_478),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_648),
.B(n_553),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_597),
.B(n_478),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_625),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_650),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_720),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_665),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_678),
.B(n_408),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_667),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_597),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_719),
.B(n_384),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_689),
.A2(n_530),
.B1(n_521),
.B2(n_538),
.Y(n_873)
);

NAND2x1p5_ASAP7_75t_L g874 ( 
.A(n_708),
.B(n_570),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_657),
.B(n_384),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_R g876 ( 
.A(n_692),
.B(n_78),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_669),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_673),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_723),
.A2(n_538),
.B1(n_527),
.B2(n_530),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_720),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_676),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_677),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_594),
.B(n_527),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_682),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_632),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_701),
.Y(n_886)
);

NOR2x1_ASAP7_75t_L g887 ( 
.A(n_708),
.B(n_549),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_698),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_596),
.A2(n_421),
.B1(n_549),
.B2(n_568),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_721),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_720),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_605),
.A2(n_421),
.B(n_568),
.C(n_570),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_596),
.A2(n_568),
.B1(n_384),
.B2(n_576),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_743),
.A2(n_702),
.B1(n_703),
.B2(n_709),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_743),
.A2(n_644),
.B(n_639),
.C(n_634),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_849),
.A2(n_716),
.B(n_717),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_728),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_752),
.A2(n_635),
.B1(n_642),
.B2(n_725),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_804),
.A2(n_718),
.B(n_726),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_747),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_751),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_734),
.B(n_727),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_808),
.B(n_722),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_756),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_752),
.A2(n_722),
.B1(n_712),
.B2(n_545),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_757),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_811),
.B(n_750),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_734),
.B(n_10),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_763),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_765),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_849),
.A2(n_576),
.B(n_545),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_810),
.B(n_11),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_814),
.A2(n_545),
.B1(n_525),
.B2(n_15),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_885),
.B(n_838),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_858),
.B(n_11),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_859),
.B(n_14),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_773),
.B(n_16),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_865),
.B(n_16),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_843),
.B(n_525),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_811),
.B(n_576),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_749),
.A2(n_545),
.B(n_525),
.C(n_22),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_749),
.A2(n_525),
.B(n_20),
.C(n_23),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_SL g923 ( 
.A1(n_860),
.A2(n_132),
.B(n_127),
.C(n_126),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_771),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_728),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_746),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_809),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_742),
.B(n_17),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_728),
.Y(n_929)
);

BUFx2_ASAP7_75t_SL g930 ( 
.A(n_779),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_783),
.A2(n_121),
.B(n_117),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_839),
.A2(n_822),
.B(n_823),
.Y(n_932)
);

NAND3xp33_ASAP7_75t_SL g933 ( 
.A(n_846),
.B(n_20),
.C(n_23),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_826),
.A2(n_116),
.B(n_101),
.Y(n_934)
);

OA22x2_ASAP7_75t_L g935 ( 
.A1(n_788),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_935)
);

O2A1O1Ixp5_ASAP7_75t_L g936 ( 
.A1(n_860),
.A2(n_84),
.B(n_73),
.C(n_32),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_794),
.B(n_819),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_817),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_769),
.A2(n_25),
.B(n_31),
.C(n_32),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_829),
.A2(n_31),
.B(n_33),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_830),
.A2(n_34),
.B(n_37),
.Y(n_941)
);

NOR2xp67_ASAP7_75t_L g942 ( 
.A(n_748),
.B(n_34),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_835),
.B(n_888),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_773),
.B(n_797),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_866),
.B(n_870),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_877),
.B(n_878),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_801),
.B(n_828),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_766),
.B(n_780),
.Y(n_948)
);

O2A1O1Ixp5_ASAP7_75t_SL g949 ( 
.A1(n_785),
.A2(n_812),
.B(n_777),
.C(n_845),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_735),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_737),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_833),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_769),
.A2(n_814),
.B(n_863),
.C(n_852),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_736),
.A2(n_775),
.B1(n_847),
.B2(n_862),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_861),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_857),
.A2(n_793),
.B(n_869),
.C(n_797),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_R g957 ( 
.A(n_815),
.B(n_824),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_761),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_781),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_767),
.A2(n_733),
.B(n_834),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_857),
.A2(n_798),
.B(n_792),
.C(n_796),
.Y(n_961)
);

OR2x6_ASAP7_75t_L g962 ( 
.A(n_745),
.B(n_800),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_805),
.B(n_732),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_764),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_868),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_882),
.B(n_884),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_881),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_821),
.A2(n_836),
.B(n_847),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_790),
.B(n_770),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_754),
.A2(n_852),
.B(n_807),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_832),
.A2(n_887),
.B(n_813),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_855),
.B(n_790),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_736),
.A2(n_795),
.B1(n_879),
.B2(n_873),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_SL g974 ( 
.A1(n_863),
.A2(n_770),
.B(n_776),
.C(n_803),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_805),
.B(n_806),
.Y(n_975)
);

OAI21xp33_ASAP7_75t_L g976 ( 
.A1(n_841),
.A2(n_799),
.B(n_778),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_778),
.B(n_776),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_728),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_795),
.A2(n_879),
.B1(n_873),
.B2(n_871),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_741),
.A2(n_871),
.B1(n_848),
.B2(n_851),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_886),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_825),
.A2(n_842),
.B(n_741),
.C(n_851),
.Y(n_982)
);

NAND3xp33_ASAP7_75t_L g983 ( 
.A(n_842),
.B(n_802),
.C(n_774),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_820),
.A2(n_883),
.B(n_772),
.C(n_731),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_890),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_729),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_759),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_759),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_745),
.B(n_753),
.Y(n_989)
);

OAI22xp33_ASAP7_75t_L g990 ( 
.A1(n_745),
.A2(n_803),
.B1(n_738),
.B2(n_760),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_SL g991 ( 
.A1(n_831),
.A2(n_837),
.B(n_820),
.C(n_827),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_755),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_730),
.B(n_782),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_744),
.A2(n_758),
.B(n_864),
.C(n_818),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_874),
.A2(n_854),
.B(n_816),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_874),
.A2(n_854),
.B(n_816),
.Y(n_996)
);

OA22x2_ASAP7_75t_L g997 ( 
.A1(n_787),
.A2(n_856),
.B1(n_853),
.B2(n_789),
.Y(n_997)
);

CKINVDCx8_ASAP7_75t_R g998 ( 
.A(n_739),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_744),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_SL g1000 ( 
.A(n_786),
.B(n_850),
.C(n_876),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_758),
.B(n_740),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_872),
.A2(n_844),
.B1(n_840),
.B2(n_730),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_782),
.A2(n_759),
.B1(n_762),
.B2(n_768),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_831),
.B(n_837),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_804),
.A2(n_892),
.B(n_784),
.C(n_875),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_786),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_759),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_850),
.B(n_762),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_762),
.B(n_768),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_762),
.B(n_768),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_768),
.A2(n_791),
.B1(n_867),
.B2(n_880),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_891),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_889),
.A2(n_450),
.B(n_581),
.C(n_690),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_SL g1014 ( 
.A(n_791),
.B(n_893),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_808),
.B(n_581),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_734),
.B(n_810),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_808),
.B(n_581),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_910),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_SL g1019 ( 
.A1(n_953),
.A2(n_973),
.B(n_954),
.Y(n_1019)
);

O2A1O1Ixp5_ASAP7_75t_L g1020 ( 
.A1(n_972),
.A2(n_969),
.B(n_971),
.C(n_968),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_914),
.B(n_1015),
.Y(n_1021)
);

OA21x2_ASAP7_75t_L g1022 ( 
.A1(n_932),
.A2(n_1005),
.B(n_970),
.Y(n_1022)
);

BUFx5_ASAP7_75t_L g1023 ( 
.A(n_993),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_924),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_899),
.A2(n_996),
.B(n_995),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_975),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_R g1027 ( 
.A(n_926),
.B(n_1000),
.Y(n_1027)
);

INVx3_ASAP7_75t_SL g1028 ( 
.A(n_947),
.Y(n_1028)
);

CKINVDCx11_ASAP7_75t_R g1029 ( 
.A(n_998),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_1017),
.B(n_948),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_900),
.Y(n_1031)
);

AOI21x1_ASAP7_75t_L g1032 ( 
.A1(n_960),
.A2(n_894),
.B(n_896),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_959),
.Y(n_1033)
);

AO21x2_ASAP7_75t_L g1034 ( 
.A1(n_974),
.A2(n_1002),
.B(n_991),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_907),
.B(n_963),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_SL g1036 ( 
.A1(n_982),
.A2(n_994),
.B(n_923),
.C(n_922),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_901),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_943),
.B(n_945),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_939),
.A2(n_956),
.B(n_976),
.C(n_933),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_957),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1016),
.A2(n_954),
.B1(n_973),
.B2(n_913),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_943),
.B(n_945),
.Y(n_1042)
);

CKINVDCx11_ASAP7_75t_R g1043 ( 
.A(n_947),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1016),
.A2(n_894),
.B(n_966),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_904),
.Y(n_1045)
);

AO31x2_ASAP7_75t_L g1046 ( 
.A1(n_984),
.A2(n_913),
.A3(n_921),
.B(n_895),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_944),
.B(n_935),
.Y(n_1047)
);

NAND3x1_ASAP7_75t_L g1048 ( 
.A(n_1001),
.B(n_989),
.C(n_917),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_993),
.B(n_987),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_946),
.B(n_966),
.Y(n_1050)
);

AO31x2_ASAP7_75t_L g1051 ( 
.A1(n_979),
.A2(n_919),
.A3(n_915),
.B(n_918),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_930),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_946),
.B(n_950),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1013),
.A2(n_979),
.B(n_936),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_902),
.A2(n_1008),
.B(n_964),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_906),
.B(n_909),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_948),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_935),
.B(n_997),
.Y(n_1058)
);

OAI22x1_ASAP7_75t_L g1059 ( 
.A1(n_1006),
.A2(n_983),
.B1(n_977),
.B2(n_903),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_962),
.B(n_928),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_961),
.A2(n_912),
.B(n_951),
.C(n_958),
.Y(n_1061)
);

NOR2xp67_ASAP7_75t_SL g1062 ( 
.A(n_897),
.B(n_978),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_902),
.A2(n_1014),
.B(n_990),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_980),
.B(n_916),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_908),
.B(n_999),
.Y(n_1065)
);

O2A1O1Ixp5_ASAP7_75t_SL g1066 ( 
.A1(n_986),
.A2(n_937),
.B(n_1007),
.C(n_925),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1014),
.A2(n_898),
.B(n_1009),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_962),
.B(n_942),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_927),
.B(n_965),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_962),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_931),
.A2(n_920),
.B(n_1010),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_934),
.A2(n_1004),
.B(n_1011),
.Y(n_1072)
);

BUFx8_ASAP7_75t_SL g1073 ( 
.A(n_1012),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_938),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1003),
.A2(n_911),
.B(n_905),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_992),
.A2(n_925),
.B(n_929),
.Y(n_1076)
);

OR2x6_ASAP7_75t_L g1077 ( 
.A(n_897),
.B(n_978),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_952),
.B(n_955),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_967),
.B(n_981),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_940),
.A2(n_941),
.B(n_985),
.C(n_929),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_897),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_978),
.B(n_988),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_988),
.A2(n_968),
.B(n_932),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_924),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_968),
.A2(n_932),
.B(n_970),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_945),
.B(n_946),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_L g1087 ( 
.A(n_953),
.B(n_450),
.C(n_439),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_926),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_924),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_899),
.A2(n_996),
.B(n_995),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_897),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_953),
.A2(n_1013),
.B(n_603),
.C(n_743),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_945),
.B(n_946),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_953),
.A2(n_968),
.B(n_949),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_953),
.A2(n_968),
.B(n_949),
.Y(n_1095)
);

O2A1O1Ixp5_ASAP7_75t_SL g1096 ( 
.A1(n_972),
.A2(n_450),
.B(n_381),
.C(n_656),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_899),
.A2(n_996),
.B(n_995),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_953),
.A2(n_968),
.B(n_949),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_945),
.B(n_946),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_968),
.A2(n_932),
.B(n_970),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_914),
.B(n_321),
.Y(n_1101)
);

INVx3_ASAP7_75t_SL g1102 ( 
.A(n_926),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_910),
.Y(n_1103)
);

AOI221xp5_ASAP7_75t_L g1104 ( 
.A1(n_953),
.A2(n_450),
.B1(n_663),
.B2(n_456),
.C(n_402),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_968),
.A2(n_932),
.B(n_970),
.Y(n_1105)
);

AO22x2_ASAP7_75t_L g1106 ( 
.A1(n_913),
.A2(n_954),
.B1(n_973),
.B2(n_933),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_899),
.A2(n_996),
.B(n_995),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_926),
.Y(n_1108)
);

AO32x2_ASAP7_75t_L g1109 ( 
.A1(n_913),
.A2(n_954),
.A3(n_973),
.B1(n_979),
.B2(n_894),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_899),
.A2(n_996),
.B(n_995),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_971),
.A2(n_968),
.B(n_970),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_926),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_953),
.A2(n_968),
.B(n_949),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1016),
.A2(n_743),
.B1(n_814),
.B2(n_734),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_993),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_914),
.B(n_808),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_R g1117 ( 
.A(n_926),
.B(n_584),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_899),
.A2(n_996),
.B(n_995),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_945),
.B(n_946),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_924),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_897),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_945),
.B(n_946),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_968),
.A2(n_932),
.B(n_970),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_968),
.A2(n_932),
.B(n_970),
.Y(n_1124)
);

AND2x6_ASAP7_75t_L g1125 ( 
.A(n_993),
.B(n_897),
.Y(n_1125)
);

BUFx10_ASAP7_75t_L g1126 ( 
.A(n_1001),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_945),
.B(n_946),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1005),
.A2(n_953),
.A3(n_954),
.B(n_968),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_968),
.A2(n_932),
.B(n_970),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_924),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_907),
.B(n_517),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1016),
.A2(n_743),
.B1(n_814),
.B2(n_734),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_945),
.B(n_946),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_945),
.B(n_946),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_953),
.A2(n_968),
.B(n_949),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_926),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_910),
.Y(n_1137)
);

OAI22x1_ASAP7_75t_L g1138 ( 
.A1(n_972),
.A2(n_846),
.B1(n_732),
.B2(n_788),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_953),
.A2(n_968),
.B(n_949),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_993),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_968),
.A2(n_932),
.B(n_970),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_897),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_945),
.B(n_946),
.Y(n_1143)
);

AOI221xp5_ASAP7_75t_L g1144 ( 
.A1(n_1104),
.A2(n_1087),
.B1(n_1041),
.B2(n_1039),
.C(n_1092),
.Y(n_1144)
);

OR2x6_ASAP7_75t_L g1145 ( 
.A(n_1019),
.B(n_1063),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_1029),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1056),
.Y(n_1147)
);

AOI221xp5_ASAP7_75t_L g1148 ( 
.A1(n_1087),
.A2(n_1041),
.B1(n_1106),
.B2(n_1054),
.C(n_1021),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1038),
.A2(n_1042),
.B1(n_1050),
.B2(n_1143),
.Y(n_1149)
);

AOI22x1_ASAP7_75t_L g1150 ( 
.A1(n_1059),
.A2(n_1044),
.B1(n_1138),
.B2(n_1106),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1086),
.A2(n_1143),
.B1(n_1093),
.B2(n_1099),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_1055),
.B(n_1067),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1083),
.A2(n_1097),
.B(n_1110),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1088),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1031),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1086),
.A2(n_1119),
.B1(n_1099),
.B2(n_1134),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1025),
.A2(n_1107),
.B(n_1118),
.Y(n_1157)
);

AOI221xp5_ASAP7_75t_L g1158 ( 
.A1(n_1054),
.A2(n_1132),
.B1(n_1114),
.B2(n_1093),
.C(n_1119),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1122),
.B(n_1127),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1114),
.A2(n_1132),
.B(n_1134),
.C(n_1133),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1070),
.B(n_1057),
.Y(n_1161)
);

AO21x2_ASAP7_75t_L g1162 ( 
.A1(n_1123),
.A2(n_1141),
.B(n_1124),
.Y(n_1162)
);

BUFx3_ASAP7_75t_L g1163 ( 
.A(n_1073),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1133),
.B(n_1053),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_1125),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1035),
.B(n_1058),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1120),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1047),
.A2(n_1064),
.B1(n_1116),
.B2(n_1094),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1142),
.B(n_1062),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_1129),
.A2(n_1080),
.A3(n_1061),
.B(n_1075),
.Y(n_1170)
);

OA21x2_ASAP7_75t_L g1171 ( 
.A1(n_1094),
.A2(n_1139),
.B(n_1095),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1111),
.A2(n_1032),
.B(n_1072),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1071),
.A2(n_1076),
.B(n_1020),
.Y(n_1173)
);

INVxp67_ASAP7_75t_SL g1174 ( 
.A(n_1022),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1066),
.A2(n_1135),
.B(n_1098),
.Y(n_1175)
);

OA21x2_ASAP7_75t_L g1176 ( 
.A1(n_1113),
.A2(n_1139),
.B(n_1064),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1108),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1113),
.A2(n_1096),
.B(n_1022),
.Y(n_1178)
);

AO21x2_ASAP7_75t_L g1179 ( 
.A1(n_1034),
.A2(n_1036),
.B(n_1065),
.Y(n_1179)
);

AO21x1_ASAP7_75t_L g1180 ( 
.A1(n_1060),
.A2(n_1082),
.B(n_1130),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1101),
.A2(n_1030),
.B1(n_1026),
.B2(n_1048),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1024),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1079),
.A2(n_1078),
.B(n_1069),
.Y(n_1183)
);

CKINVDCx11_ASAP7_75t_R g1184 ( 
.A(n_1112),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_1037),
.A2(n_1084),
.B(n_1045),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1089),
.A2(n_1049),
.B(n_1074),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1034),
.A2(n_1109),
.A3(n_1051),
.B(n_1128),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_1103),
.B(n_1018),
.Y(n_1188)
);

OAI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1028),
.A2(n_1052),
.B1(n_1137),
.B2(n_1068),
.C(n_1102),
.Y(n_1189)
);

OA21x2_ASAP7_75t_L g1190 ( 
.A1(n_1109),
.A2(n_1128),
.B(n_1051),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1049),
.A2(n_1140),
.B(n_1115),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1077),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1027),
.A2(n_1043),
.B1(n_1126),
.B2(n_1115),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1140),
.A2(n_1128),
.B(n_1046),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1125),
.A2(n_1121),
.B(n_1040),
.Y(n_1195)
);

OA21x2_ASAP7_75t_L g1196 ( 
.A1(n_1109),
.A2(n_1051),
.B(n_1046),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1046),
.A2(n_1023),
.B(n_1125),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1023),
.A2(n_1125),
.B(n_1077),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1142),
.B(n_1033),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1142),
.A2(n_1136),
.B1(n_1081),
.B2(n_1091),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1023),
.A2(n_1091),
.B(n_1126),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1023),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1117),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1092),
.A2(n_1100),
.A3(n_1105),
.B(n_1085),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1092),
.A2(n_450),
.B(n_953),
.C(n_1039),
.Y(n_1205)
);

NOR2x1_ASAP7_75t_R g1206 ( 
.A(n_1029),
.B(n_724),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1104),
.A2(n_1087),
.B1(n_935),
.B2(n_1106),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_1131),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1083),
.A2(n_1090),
.B(n_1025),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1035),
.B(n_1058),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1026),
.B(n_1021),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_R g1212 ( 
.A(n_1112),
.B(n_926),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1056),
.Y(n_1213)
);

AOI222xp33_ASAP7_75t_L g1214 ( 
.A1(n_1104),
.A2(n_418),
.B1(n_450),
.B2(n_191),
.C1(n_163),
.C2(n_690),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1104),
.A2(n_743),
.B(n_1092),
.C(n_953),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1104),
.A2(n_1087),
.B1(n_935),
.B2(n_1106),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1038),
.B(n_1042),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_1112),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_SL g1219 ( 
.A1(n_1138),
.A2(n_492),
.B1(n_418),
.B2(n_507),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1083),
.A2(n_1090),
.B(n_1025),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_1094),
.A2(n_1098),
.B(n_1095),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1021),
.B(n_321),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1073),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1083),
.A2(n_1090),
.B(n_1025),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1131),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1083),
.A2(n_1090),
.B(n_1025),
.Y(n_1226)
);

OA21x2_ASAP7_75t_L g1227 ( 
.A1(n_1094),
.A2(n_1098),
.B(n_1095),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1031),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1083),
.A2(n_1090),
.B(n_1025),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1088),
.Y(n_1230)
);

OAI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1104),
.A2(n_935),
.B1(n_1042),
.B2(n_1038),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1056),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1033),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1131),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1033),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1125),
.Y(n_1236)
);

OA21x2_ASAP7_75t_L g1237 ( 
.A1(n_1094),
.A2(n_1098),
.B(n_1095),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1083),
.A2(n_1090),
.B(n_1025),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1056),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1056),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1104),
.A2(n_1087),
.B1(n_935),
.B2(n_1106),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1033),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1033),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1142),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1087),
.A2(n_439),
.B(n_1092),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_1112),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1092),
.A2(n_1100),
.A3(n_1105),
.B(n_1085),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1087),
.A2(n_935),
.B1(n_418),
.B2(n_492),
.Y(n_1248)
);

OR2x6_ASAP7_75t_L g1249 ( 
.A(n_1019),
.B(n_1063),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1056),
.Y(n_1250)
);

INVx6_ASAP7_75t_L g1251 ( 
.A(n_1142),
.Y(n_1251)
);

OAI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1104),
.A2(n_935),
.B1(n_1042),
.B2(n_1038),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1094),
.A2(n_1098),
.B(n_1095),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1038),
.B(n_1042),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1051),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1159),
.B(n_1217),
.Y(n_1256)
);

INVxp67_ASAP7_75t_L g1257 ( 
.A(n_1211),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1185),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_SL g1259 ( 
.A1(n_1149),
.A2(n_1215),
.B(n_1254),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1166),
.B(n_1210),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1184),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1248),
.A2(n_1241),
.B1(n_1216),
.B2(n_1207),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1159),
.B(n_1164),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1208),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1147),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1213),
.B(n_1232),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1239),
.B(n_1240),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1255),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1182),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_1194),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1151),
.B(n_1156),
.Y(n_1271)
);

NOR2xp67_ASAP7_75t_L g1272 ( 
.A(n_1203),
.B(n_1189),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1225),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1248),
.A2(n_1241),
.B1(n_1216),
.B2(n_1207),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1188),
.Y(n_1275)
);

BUFx2_ASAP7_75t_SL g1276 ( 
.A(n_1218),
.Y(n_1276)
);

AOI21x1_ASAP7_75t_SL g1277 ( 
.A1(n_1161),
.A2(n_1150),
.B(n_1214),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1199),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1231),
.B(n_1252),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1245),
.A2(n_1215),
.B(n_1162),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1173),
.A2(n_1148),
.B(n_1174),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1168),
.A2(n_1193),
.B1(n_1252),
.B2(n_1231),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1205),
.A2(n_1181),
.B(n_1144),
.C(n_1222),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1168),
.A2(n_1193),
.B1(n_1219),
.B2(n_1222),
.Y(n_1284)
);

AOI21x1_ASAP7_75t_SL g1285 ( 
.A1(n_1205),
.A2(n_1179),
.B(n_1180),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1250),
.B(n_1234),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1228),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1218),
.A2(n_1246),
.B1(n_1203),
.B2(n_1146),
.Y(n_1288)
);

NOR2xp67_ASAP7_75t_L g1289 ( 
.A(n_1233),
.B(n_1235),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1144),
.A2(n_1160),
.B(n_1249),
.C(n_1145),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1155),
.Y(n_1291)
);

NOR2x1_ASAP7_75t_SL g1292 ( 
.A(n_1145),
.B(n_1249),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1184),
.Y(n_1293)
);

OAI31xp33_ASAP7_75t_L g1294 ( 
.A1(n_1160),
.A2(n_1200),
.A3(n_1199),
.B(n_1242),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1167),
.B(n_1176),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1148),
.A2(n_1158),
.B1(n_1243),
.B2(n_1195),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1212),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1202),
.B(n_1198),
.Y(n_1298)
);

BUFx12f_ASAP7_75t_L g1299 ( 
.A(n_1154),
.Y(n_1299)
);

NOR2xp67_ASAP7_75t_L g1300 ( 
.A(n_1177),
.B(n_1230),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1169),
.A2(n_1244),
.B(n_1201),
.Y(n_1301)
);

A2O1A1Ixp33_ASAP7_75t_SL g1302 ( 
.A1(n_1202),
.A2(n_1201),
.B(n_1236),
.C(n_1165),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1204),
.Y(n_1303)
);

OA21x2_ASAP7_75t_L g1304 ( 
.A1(n_1157),
.A2(n_1209),
.B(n_1153),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1197),
.B(n_1192),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1251),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1176),
.B(n_1246),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1186),
.B(n_1183),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1165),
.A2(n_1236),
.B1(n_1169),
.B2(n_1251),
.Y(n_1309)
);

OR2x6_ASAP7_75t_L g1310 ( 
.A(n_1152),
.B(n_1191),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_R g1311 ( 
.A(n_1244),
.B(n_1163),
.Y(n_1311)
);

NOR2xp67_ASAP7_75t_L g1312 ( 
.A(n_1163),
.B(n_1223),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1223),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1220),
.B(n_1224),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1212),
.B(n_1171),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1221),
.B(n_1227),
.Y(n_1316)
);

OA21x2_ASAP7_75t_L g1317 ( 
.A1(n_1226),
.A2(n_1229),
.B(n_1238),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1237),
.B(n_1253),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1170),
.A2(n_1196),
.B(n_1253),
.C(n_1237),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1253),
.A2(n_1196),
.B1(n_1190),
.B2(n_1206),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1187),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1187),
.B(n_1247),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1166),
.B(n_1210),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1166),
.B(n_1210),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1175),
.A2(n_1178),
.B(n_1172),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_SL g1326 ( 
.A1(n_1149),
.A2(n_1092),
.B(n_953),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1166),
.B(n_1210),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1316),
.B(n_1318),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1305),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1262),
.A2(n_1274),
.B1(n_1282),
.B2(n_1284),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1258),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1321),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1295),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1279),
.A2(n_1296),
.B1(n_1271),
.B2(n_1280),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1322),
.B(n_1319),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1298),
.B(n_1305),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1303),
.B(n_1307),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1270),
.Y(n_1338)
);

BUFx12f_ASAP7_75t_L g1339 ( 
.A(n_1261),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1270),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1268),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1298),
.B(n_1305),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1310),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1310),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1310),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1308),
.Y(n_1346)
);

AO21x2_ASAP7_75t_L g1347 ( 
.A1(n_1320),
.A2(n_1315),
.B(n_1326),
.Y(n_1347)
);

OA21x2_ASAP7_75t_L g1348 ( 
.A1(n_1269),
.A2(n_1291),
.B(n_1298),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1281),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1283),
.A2(n_1290),
.B(n_1259),
.Y(n_1350)
);

OR2x6_ASAP7_75t_L g1351 ( 
.A(n_1314),
.B(n_1301),
.Y(n_1351)
);

AO21x2_ASAP7_75t_L g1352 ( 
.A1(n_1302),
.A2(n_1292),
.B(n_1285),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1281),
.B(n_1325),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1314),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1325),
.B(n_1287),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1265),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1278),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1304),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1317),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1263),
.B(n_1256),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1337),
.B(n_1257),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1333),
.B(n_1265),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1331),
.Y(n_1363)
);

AO22x1_ASAP7_75t_L g1364 ( 
.A1(n_1350),
.A2(n_1309),
.B1(n_1278),
.B2(n_1261),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1328),
.B(n_1257),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1328),
.B(n_1260),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1328),
.B(n_1327),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1337),
.B(n_1286),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1346),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1336),
.B(n_1323),
.Y(n_1370)
);

INVxp67_ASAP7_75t_L g1371 ( 
.A(n_1346),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1343),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1336),
.B(n_1324),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1348),
.Y(n_1374)
);

NOR2x1_ASAP7_75t_R g1375 ( 
.A(n_1339),
.B(n_1293),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1336),
.B(n_1266),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1331),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1336),
.B(n_1267),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1343),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1348),
.Y(n_1380)
);

NOR2xp67_ASAP7_75t_SL g1381 ( 
.A(n_1350),
.B(n_1293),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1348),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1348),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1337),
.B(n_1275),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1348),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1355),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1372),
.Y(n_1387)
);

NAND4xp25_ASAP7_75t_L g1388 ( 
.A(n_1384),
.B(n_1330),
.C(n_1334),
.D(n_1360),
.Y(n_1388)
);

OAI33xp33_ASAP7_75t_L g1389 ( 
.A1(n_1362),
.A2(n_1360),
.A3(n_1335),
.B1(n_1341),
.B2(n_1338),
.B3(n_1340),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1384),
.A2(n_1330),
.B1(n_1334),
.B2(n_1272),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_R g1391 ( 
.A(n_1384),
.B(n_1297),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1361),
.B(n_1335),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1381),
.A2(n_1294),
.B(n_1362),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1368),
.B(n_1356),
.Y(n_1394)
);

OAI221xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1368),
.A2(n_1335),
.B1(n_1349),
.B2(n_1351),
.C(n_1344),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1375),
.B(n_1297),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1382),
.Y(n_1397)
);

AOI211xp5_ASAP7_75t_L g1398 ( 
.A1(n_1381),
.A2(n_1288),
.B(n_1349),
.C(n_1344),
.Y(n_1398)
);

OAI33xp33_ASAP7_75t_L g1399 ( 
.A1(n_1361),
.A2(n_1341),
.A3(n_1338),
.B1(n_1340),
.B2(n_1333),
.B3(n_1332),
.Y(n_1399)
);

NOR2x1p5_ASAP7_75t_L g1400 ( 
.A(n_1375),
.B(n_1339),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1368),
.B(n_1339),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1381),
.A2(n_1347),
.B1(n_1345),
.B2(n_1343),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1372),
.Y(n_1403)
);

OAI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1361),
.A2(n_1345),
.B1(n_1344),
.B2(n_1276),
.C(n_1264),
.Y(n_1404)
);

AO21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1380),
.A2(n_1341),
.B(n_1340),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1363),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1372),
.A2(n_1349),
.B(n_1277),
.C(n_1345),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1377),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1372),
.B(n_1329),
.Y(n_1409)
);

OAI321xp33_ASAP7_75t_L g1410 ( 
.A1(n_1369),
.A2(n_1351),
.A3(n_1354),
.B1(n_1338),
.B2(n_1353),
.C(n_1333),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1369),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1379),
.B(n_1357),
.Y(n_1412)
);

OA21x2_ASAP7_75t_L g1413 ( 
.A1(n_1380),
.A2(n_1383),
.B(n_1385),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1370),
.A2(n_1347),
.B1(n_1342),
.B2(n_1336),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1363),
.Y(n_1415)
);

OAI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1379),
.A2(n_1273),
.B1(n_1289),
.B2(n_1351),
.C(n_1354),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1386),
.B(n_1347),
.Y(n_1417)
);

AOI221xp5_ASAP7_75t_L g1418 ( 
.A1(n_1364),
.A2(n_1366),
.B1(n_1367),
.B2(n_1365),
.C(n_1347),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1371),
.Y(n_1419)
);

OAI31xp33_ASAP7_75t_L g1420 ( 
.A1(n_1379),
.A2(n_1354),
.A3(n_1306),
.B(n_1313),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1376),
.B(n_1336),
.Y(n_1421)
);

AO21x2_ASAP7_75t_L g1422 ( 
.A1(n_1383),
.A2(n_1358),
.B(n_1359),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1413),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1403),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1405),
.B(n_1386),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1405),
.B(n_1386),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1408),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1408),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1406),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1413),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1413),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1421),
.B(n_1386),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1392),
.B(n_1365),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1415),
.Y(n_1434)
);

NAND3xp33_ASAP7_75t_L g1435 ( 
.A(n_1390),
.B(n_1364),
.C(n_1374),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1411),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1388),
.B(n_1370),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1419),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1422),
.Y(n_1439)
);

INVx4_ASAP7_75t_SL g1440 ( 
.A(n_1387),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1392),
.B(n_1365),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1403),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1399),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1422),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1394),
.B(n_1371),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1422),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1407),
.A2(n_1351),
.B(n_1352),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1397),
.Y(n_1448)
);

INVx4_ASAP7_75t_L g1449 ( 
.A(n_1403),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1427),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1437),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1427),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1429),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1425),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1440),
.B(n_1421),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1428),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1428),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1429),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1425),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1424),
.Y(n_1460)
);

AND3x2_ASAP7_75t_L g1461 ( 
.A(n_1442),
.B(n_1398),
.C(n_1396),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1434),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1424),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1434),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1437),
.B(n_1367),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1436),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1443),
.B(n_1367),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1436),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1440),
.B(n_1400),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1440),
.B(n_1409),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1440),
.B(n_1409),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1438),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1425),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1443),
.B(n_1370),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1440),
.B(n_1409),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1438),
.B(n_1373),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1445),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1435),
.B(n_1339),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1445),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1448),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1433),
.B(n_1417),
.Y(n_1481)
);

NAND2xp33_ASAP7_75t_L g1482 ( 
.A(n_1435),
.B(n_1393),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1440),
.B(n_1412),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1442),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1442),
.B(n_1418),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1441),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1448),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1432),
.B(n_1414),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1432),
.B(n_1401),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1426),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1474),
.B(n_1441),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1467),
.B(n_1373),
.Y(n_1492)
);

INVxp67_ASAP7_75t_L g1493 ( 
.A(n_1463),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1450),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1463),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1460),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1454),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1484),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1469),
.B(n_1449),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1482),
.B(n_1373),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1450),
.Y(n_1501)
);

INVx4_ASAP7_75t_L g1502 ( 
.A(n_1469),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1452),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1469),
.B(n_1449),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1452),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1483),
.B(n_1449),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1456),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1479),
.B(n_1449),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1456),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1478),
.B(n_1391),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1483),
.B(n_1449),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1482),
.B(n_1376),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1483),
.B(n_1426),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1470),
.B(n_1426),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1454),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1477),
.B(n_1479),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1461),
.B(n_1376),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1457),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1486),
.B(n_1472),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1457),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1462),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1470),
.B(n_1471),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1485),
.B(n_1378),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1462),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1464),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1494),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1491),
.B(n_1492),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1513),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1510),
.B(n_1451),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1495),
.B(n_1493),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1522),
.B(n_1471),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1522),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1494),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1501),
.Y(n_1534)
);

AOI222xp33_ASAP7_75t_L g1535 ( 
.A1(n_1496),
.A2(n_1485),
.B1(n_1389),
.B2(n_1466),
.C1(n_1468),
.C2(n_1488),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1501),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1491),
.B(n_1466),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1503),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1511),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1513),
.B(n_1475),
.Y(n_1540)
);

AO21x2_ASAP7_75t_L g1541 ( 
.A1(n_1521),
.A2(n_1447),
.B(n_1430),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1498),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1503),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1505),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1514),
.B(n_1475),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1517),
.A2(n_1407),
.B(n_1468),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1514),
.B(n_1455),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1505),
.Y(n_1548)
);

NOR2xp67_ASAP7_75t_SL g1549 ( 
.A(n_1502),
.B(n_1299),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1502),
.B(n_1455),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1526),
.Y(n_1551)
);

OAI21xp33_ASAP7_75t_L g1552 ( 
.A1(n_1532),
.A2(n_1498),
.B(n_1516),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1547),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1531),
.B(n_1502),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1526),
.Y(n_1555)
);

AOI322xp5_ASAP7_75t_L g1556 ( 
.A1(n_1542),
.A2(n_1512),
.A3(n_1500),
.B1(n_1523),
.B2(n_1488),
.C1(n_1465),
.C2(n_1511),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1530),
.Y(n_1557)
);

OAI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1546),
.A2(n_1410),
.B1(n_1416),
.B2(n_1404),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1539),
.B(n_1506),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1529),
.A2(n_1299),
.B1(n_1313),
.B2(n_1506),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1528),
.B(n_1506),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1533),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1550),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1535),
.A2(n_1504),
.B1(n_1499),
.B2(n_1402),
.Y(n_1564)
);

AOI221xp5_ASAP7_75t_L g1565 ( 
.A1(n_1528),
.A2(n_1525),
.B1(n_1524),
.B2(n_1521),
.C(n_1509),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1531),
.B(n_1499),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1538),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1533),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1527),
.B(n_1519),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1554),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1568),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1566),
.B(n_1540),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1557),
.B(n_1549),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1568),
.Y(n_1574)
);

NOR2x1p5_ASAP7_75t_L g1575 ( 
.A(n_1559),
.B(n_1550),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1553),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1563),
.B(n_1540),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1557),
.B(n_1545),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1551),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_1561),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_SL g1581 ( 
.A1(n_1570),
.A2(n_1560),
.B1(n_1567),
.B2(n_1564),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1571),
.Y(n_1582)
);

AOI322xp5_ASAP7_75t_L g1583 ( 
.A1(n_1574),
.A2(n_1558),
.A3(n_1552),
.B1(n_1567),
.B2(n_1565),
.C1(n_1562),
.C2(n_1555),
.Y(n_1583)
);

AOI211xp5_ASAP7_75t_L g1584 ( 
.A1(n_1573),
.A2(n_1549),
.B(n_1569),
.C(n_1504),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1572),
.A2(n_1541),
.B1(n_1545),
.B2(n_1547),
.Y(n_1585)
);

AOI21xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1578),
.A2(n_1541),
.B(n_1537),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_SL g1587 ( 
.A1(n_1573),
.A2(n_1556),
.B(n_1548),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1577),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1575),
.Y(n_1589)
);

OAI21xp33_ASAP7_75t_L g1590 ( 
.A1(n_1570),
.A2(n_1527),
.B(n_1537),
.Y(n_1590)
);

O2A1O1Ixp33_ASAP7_75t_L g1591 ( 
.A1(n_1580),
.A2(n_1541),
.B(n_1544),
.C(n_1543),
.Y(n_1591)
);

NAND2xp33_ASAP7_75t_R g1592 ( 
.A(n_1588),
.B(n_1311),
.Y(n_1592)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1593 ( 
.A1(n_1590),
.A2(n_1576),
.B(n_1579),
.C(n_1543),
.D(n_1536),
.Y(n_1593)
);

AOI221xp5_ASAP7_75t_L g1594 ( 
.A1(n_1587),
.A2(n_1580),
.B1(n_1534),
.B2(n_1536),
.C(n_1525),
.Y(n_1594)
);

OAI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1585),
.A2(n_1508),
.B1(n_1519),
.B2(n_1490),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1581),
.A2(n_1497),
.B1(n_1515),
.B2(n_1534),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1596),
.Y(n_1597)
);

NOR2x1_ASAP7_75t_L g1598 ( 
.A(n_1595),
.B(n_1591),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1594),
.B(n_1589),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1592),
.B(n_1584),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1593),
.B(n_1582),
.Y(n_1601)
);

NOR3xp33_ASAP7_75t_L g1602 ( 
.A(n_1595),
.B(n_1586),
.C(n_1583),
.Y(n_1602)
);

AOI211xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1601),
.A2(n_1312),
.B(n_1508),
.C(n_1524),
.Y(n_1603)
);

OAI211xp5_ASAP7_75t_L g1604 ( 
.A1(n_1602),
.A2(n_1311),
.B(n_1300),
.C(n_1497),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1600),
.B(n_1489),
.Y(n_1605)
);

O2A1O1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1598),
.A2(n_1520),
.B(n_1518),
.C(n_1507),
.Y(n_1606)
);

OAI221xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1599),
.A2(n_1515),
.B1(n_1518),
.B2(n_1520),
.C(n_1509),
.Y(n_1607)
);

OAI221xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1604),
.A2(n_1597),
.B1(n_1507),
.B2(n_1420),
.C(n_1459),
.Y(n_1608)
);

NAND2xp33_ASAP7_75t_R g1609 ( 
.A(n_1605),
.B(n_1489),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1603),
.B(n_1459),
.Y(n_1610)
);

NAND5xp2_ASAP7_75t_L g1611 ( 
.A(n_1608),
.B(n_1606),
.C(n_1607),
.D(n_1395),
.E(n_1464),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1611),
.A2(n_1609),
.B1(n_1610),
.B2(n_1473),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1612),
.Y(n_1613)
);

XNOR2xp5_ASAP7_75t_L g1614 ( 
.A(n_1613),
.B(n_1473),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1614),
.B(n_1490),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1615),
.Y(n_1616)
);

XNOR2xp5_ASAP7_75t_L g1617 ( 
.A(n_1615),
.B(n_1306),
.Y(n_1617)
);

OAI22xp33_ASAP7_75t_SL g1618 ( 
.A1(n_1616),
.A2(n_1453),
.B1(n_1458),
.B2(n_1487),
.Y(n_1618)
);

XNOR2x1_ASAP7_75t_L g1619 ( 
.A(n_1617),
.B(n_1481),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1619),
.B(n_1480),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1618),
.B(n_1480),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1620),
.A2(n_1487),
.B(n_1476),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1622),
.A2(n_1621),
.B1(n_1431),
.B2(n_1423),
.Y(n_1623)
);

AOI211xp5_ASAP7_75t_L g1624 ( 
.A1(n_1623),
.A2(n_1439),
.B(n_1444),
.C(n_1446),
.Y(n_1624)
);


endmodule