module fake_jpeg_3449_n_525 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_3),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_47),
.Y(n_130)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_50),
.Y(n_146)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_53),
.Y(n_147)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_55),
.Y(n_136)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_58),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_59),
.Y(n_148)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_34),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_66),
.A2(n_75),
.B1(n_96),
.B2(n_33),
.Y(n_144)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_35),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_15),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_15),
.Y(n_112)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_94),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_7),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_39),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_97),
.B(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_25),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_101),
.B(n_112),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_46),
.A2(n_39),
.B1(n_33),
.B2(n_38),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_103),
.A2(n_119),
.B1(n_32),
.B2(n_26),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_24),
.B1(n_44),
.B2(n_43),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_106),
.B(n_122),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_47),
.A2(n_39),
.B1(n_33),
.B2(n_37),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_24),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_63),
.B(n_45),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_68),
.B(n_45),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_85),
.B(n_41),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_144),
.A2(n_19),
.B1(n_31),
.B2(n_25),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_60),
.Y(n_203)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_138),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_158),
.B(n_164),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_98),
.A2(n_53),
.B1(n_48),
.B2(n_54),
.Y(n_159)
);

AO21x1_ASAP7_75t_SL g233 ( 
.A1(n_159),
.A2(n_61),
.B(n_50),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_103),
.A2(n_69),
.B1(n_59),
.B2(n_58),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_160),
.A2(n_195),
.B1(n_197),
.B2(n_200),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_165),
.Y(n_206)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_125),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_135),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_171),
.B(n_183),
.Y(n_222)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_173),
.A2(n_180),
.B1(n_201),
.B2(n_21),
.Y(n_225)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_182),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_179),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_98),
.A2(n_44),
.B1(n_31),
.B2(n_43),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

BUFx2_ASAP7_75t_SL g211 ( 
.A(n_181),
.Y(n_211)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_99),
.B(n_83),
.C(n_70),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_189),
.Y(n_235)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_194),
.Y(n_210)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_192),
.Y(n_208)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_105),
.A2(n_33),
.B1(n_37),
.B2(n_41),
.Y(n_195)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_198),
.Y(n_238)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_203),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_109),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_119),
.A2(n_23),
.B1(n_21),
.B2(n_29),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_202),
.A2(n_117),
.B1(n_120),
.B2(n_68),
.Y(n_237)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_102),
.A3(n_129),
.B1(n_139),
.B2(n_133),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_169),
.B(n_177),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_209),
.A2(n_218),
.B(n_176),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_145),
.B(n_116),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_118),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_176),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_23),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_173),
.A2(n_160),
.B1(n_175),
.B2(n_147),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_232),
.B1(n_234),
.B2(n_202),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_174),
.A2(n_147),
.B1(n_130),
.B2(n_155),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_233),
.A2(n_170),
.B1(n_179),
.B2(n_131),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_162),
.A2(n_130),
.B1(n_148),
.B2(n_136),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_218),
.A2(n_163),
.B(n_161),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_239),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_240),
.B(n_267),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_216),
.A2(n_155),
.B1(n_148),
.B2(n_182),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_256),
.B1(n_228),
.B2(n_234),
.Y(n_271)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_242),
.Y(n_274)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_222),
.B(n_194),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_249),
.Y(n_278)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_190),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_251),
.Y(n_286)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_227),
.Y(n_253)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_253),
.Y(n_295)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_213),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_257),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_216),
.A2(n_193),
.B1(n_186),
.B2(n_188),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_266),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_268),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_209),
.B(n_183),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_262),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_206),
.A2(n_172),
.B1(n_168),
.B2(n_199),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_263),
.B1(n_227),
.B2(n_236),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_206),
.B(n_189),
.C(n_187),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_215),
.A2(n_179),
.B(n_185),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_264),
.A2(n_210),
.B(n_235),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_205),
.A2(n_170),
.B(n_167),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_237),
.B(n_207),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_204),
.B(n_181),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_204),
.B(n_157),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_223),
.B(n_114),
.C(n_192),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_267),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_271),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_272),
.A2(n_281),
.B(n_298),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_244),
.A2(n_233),
.B1(n_207),
.B2(n_225),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_275),
.A2(n_245),
.B1(n_235),
.B2(n_231),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_277),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_SL g281 ( 
.A(n_251),
.B(n_215),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_267),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_230),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_285),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_232),
.B1(n_233),
.B2(n_217),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_288),
.A2(n_248),
.B1(n_240),
.B2(n_261),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_257),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_293),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_266),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_253),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_253),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_259),
.A2(n_217),
.B(n_230),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_264),
.B(n_239),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_299),
.A2(n_300),
.B(n_306),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_SL g300 ( 
.A(n_275),
.B(n_260),
.C(n_256),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_303),
.B(n_312),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_246),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_309),
.C(n_327),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_249),
.C(n_262),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_274),
.Y(n_310)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_310),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_279),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_279),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_314),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_290),
.Y(n_314)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_315),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_316),
.A2(n_319),
.B1(n_288),
.B2(n_287),
.Y(n_333)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_289),
.Y(n_317)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_317),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_269),
.B(n_268),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_287),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_280),
.A2(n_240),
.B1(n_245),
.B2(n_241),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_278),
.B(n_254),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_320),
.B(n_321),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_255),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_331),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_242),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_324),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_286),
.B(n_243),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_325),
.A2(n_328),
.B1(n_276),
.B2(n_295),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_231),
.C(n_238),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_280),
.A2(n_245),
.B1(n_250),
.B2(n_247),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_278),
.B(n_238),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_329),
.B(n_312),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_208),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_330),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_290),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_338),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_333),
.A2(n_348),
.B1(n_354),
.B2(n_361),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_306),
.A2(n_298),
.B(n_294),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g376 ( 
.A(n_335),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_337),
.B(n_353),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_281),
.Y(n_338)
);

XOR2x1_ASAP7_75t_SL g341 ( 
.A(n_299),
.B(n_270),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_341),
.A2(n_331),
.B1(n_314),
.B2(n_304),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_303),
.B(n_291),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_350),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_307),
.B(n_273),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_355),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_293),
.C(n_284),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_327),
.C(n_313),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_326),
.A2(n_272),
.B1(n_271),
.B2(n_277),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_315),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_305),
.A2(n_311),
.B(n_325),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_363),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_297),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_352),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_326),
.A2(n_273),
.B1(n_276),
.B2(n_296),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_309),
.B(n_296),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_295),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_358),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_308),
.B(n_229),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_212),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_326),
.A2(n_282),
.B1(n_289),
.B2(n_220),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_311),
.A2(n_304),
.B(n_302),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_370),
.Y(n_399)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_339),
.Y(n_367)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_367),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_352),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_368),
.B(n_382),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_300),
.C(n_308),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_369),
.B(n_374),
.C(n_375),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_356),
.A2(n_302),
.B1(n_316),
.B2(n_320),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_371),
.A2(n_387),
.B1(n_392),
.B2(n_334),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_329),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_373),
.B(n_184),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_321),
.C(n_324),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_332),
.B(n_338),
.C(n_347),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_339),
.Y(n_377)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_377),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_346),
.B(n_323),
.Y(n_381)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_349),
.C(n_342),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_229),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_352),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_383),
.B(n_385),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_310),
.C(n_301),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_389),
.C(n_341),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_229),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_333),
.A2(n_328),
.B1(n_317),
.B2(n_282),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_386),
.A2(n_393),
.B1(n_334),
.B2(n_220),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_356),
.A2(n_220),
.B1(n_224),
.B2(n_236),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_388),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_336),
.B(n_226),
.C(n_212),
.Y(n_389)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_391),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_363),
.A2(n_342),
.B1(n_348),
.B2(n_359),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_335),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_395),
.B(n_397),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_403),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_370),
.A2(n_359),
.B1(n_350),
.B2(n_353),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_401),
.Y(n_426)
);

OAI21xp33_ASAP7_75t_L g403 ( 
.A1(n_376),
.A2(n_362),
.B(n_354),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_392),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_420),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_362),
.C(n_360),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_410),
.C(n_415),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_371),
.A2(n_366),
.B1(n_379),
.B2(n_390),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_345),
.Y(n_409)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_409),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_360),
.C(n_345),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_411),
.A2(n_418),
.B1(n_387),
.B2(n_379),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_390),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_365),
.B(n_224),
.Y(n_413)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_413),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_364),
.B(n_221),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_416),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_373),
.B(n_208),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_417),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_372),
.A2(n_226),
.B1(n_221),
.B2(n_211),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_226),
.C(n_178),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_375),
.C(n_381),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_393),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_427),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_397),
.Y(n_425)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_425),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_402),
.B(n_401),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_419),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_384),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_429),
.B(n_430),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_394),
.B(n_389),
.C(n_376),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_433),
.A2(n_37),
.B1(n_29),
.B2(n_41),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_434),
.A2(n_431),
.B1(n_426),
.B2(n_433),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_379),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_436),
.A2(n_437),
.B(n_443),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g437 ( 
.A1(n_414),
.A2(n_400),
.B(n_396),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_394),
.B(n_386),
.C(n_154),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_441),
.C(n_415),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_399),
.B(n_198),
.C(n_166),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_442),
.B(n_398),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_405),
.B(n_10),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_445),
.B(n_455),
.Y(n_466)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_449),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_395),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_424),
.B(n_408),
.C(n_411),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_452),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_403),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_432),
.A2(n_418),
.B(n_420),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_453),
.A2(n_457),
.B(n_427),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_454),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_113),
.C(n_87),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_425),
.A2(n_92),
.B(n_89),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_88),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_458),
.B(n_459),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_428),
.B(n_90),
.C(n_95),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_211),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_200),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_32),
.C(n_26),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_461),
.B(n_439),
.C(n_435),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_431),
.A2(n_120),
.B1(n_64),
.B2(n_62),
.Y(n_462)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_462),
.Y(n_478)
);

MAJx2_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_26),
.C(n_8),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_477),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_464),
.B(n_444),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_468),
.B(n_469),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_448),
.B(n_421),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_470),
.A2(n_479),
.B1(n_461),
.B2(n_462),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_445),
.A2(n_441),
.B(n_434),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_473),
.A2(n_123),
.B(n_30),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_450),
.B(n_443),
.C(n_32),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_474),
.B(n_475),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_451),
.B(n_67),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_9),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_476),
.B(n_456),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_485),
.B(n_486),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_472),
.B(n_455),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_467),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_487),
.B(n_488),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_474),
.B(n_458),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_465),
.B(n_449),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_489),
.B(n_490),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_481),
.B(n_447),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_481),
.B(n_459),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_491),
.A2(n_495),
.B(n_6),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_492),
.A2(n_482),
.B1(n_483),
.B2(n_493),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_478),
.A2(n_460),
.B1(n_123),
.B2(n_6),
.Y(n_493)
);

INVxp33_ASAP7_75t_L g498 ( 
.A(n_493),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_30),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_466),
.B(n_5),
.Y(n_495)
);

FAx1_ASAP7_75t_SL g496 ( 
.A(n_484),
.B(n_465),
.CI(n_477),
.CON(n_496),
.SN(n_496)
);

AO21x1_ASAP7_75t_L g512 ( 
.A1(n_496),
.A2(n_10),
.B(n_1),
.Y(n_512)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_497),
.Y(n_508)
);

O2A1O1Ixp33_ASAP7_75t_SL g499 ( 
.A1(n_492),
.A2(n_482),
.B(n_480),
.C(n_479),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_499),
.A2(n_0),
.B(n_1),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_500),
.Y(n_511)
);

OAI21x1_ASAP7_75t_SL g513 ( 
.A1(n_501),
.A2(n_0),
.B(n_1),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_482),
.B(n_30),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_503),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_487),
.A2(n_6),
.B(n_15),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_506),
.A2(n_10),
.B(n_1),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_507),
.B(n_510),
.Y(n_518)
);

OAI21xp33_ASAP7_75t_L g510 ( 
.A1(n_505),
.A2(n_504),
.B(n_502),
.Y(n_510)
);

AO21x1_ASAP7_75t_L g517 ( 
.A1(n_512),
.A2(n_513),
.B(n_514),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_508),
.B(n_497),
.C(n_498),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_515),
.B(n_519),
.Y(n_521)
);

AOI321xp33_ASAP7_75t_L g516 ( 
.A1(n_509),
.A2(n_496),
.A3(n_499),
.B1(n_30),
.B2(n_4),
.C(n_2),
.Y(n_516)
);

NAND2x1p5_ASAP7_75t_SL g522 ( 
.A(n_516),
.B(n_1),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_511),
.B(n_0),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_518),
.B(n_30),
.C(n_2),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_520),
.B(n_522),
.Y(n_523)
);

O2A1O1Ixp33_ASAP7_75t_SL g524 ( 
.A1(n_523),
.A2(n_521),
.B(n_517),
.C(n_4),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_2),
.B(n_4),
.Y(n_525)
);


endmodule