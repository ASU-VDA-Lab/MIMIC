module fake_jpeg_16080_n_212 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_212);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_11),
.B(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_44),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_35),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_28),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_32),
.A2(n_0),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_60),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_16),
.B(n_2),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_65),
.Y(n_83)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_16),
.B(n_3),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_38),
.B1(n_30),
.B2(n_27),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_77),
.B1(n_84),
.B2(n_86),
.Y(n_107)
);

OAI22x1_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_24),
.B1(n_8),
.B2(n_9),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_71),
.A2(n_74),
.B1(n_75),
.B2(n_87),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_39),
.A2(n_21),
.B1(n_33),
.B2(n_31),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_38),
.B1(n_30),
.B2(n_27),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_22),
.B1(n_17),
.B2(n_25),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_90),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_40),
.A2(n_25),
.B1(n_22),
.B2(n_17),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_41),
.A2(n_33),
.B1(n_31),
.B2(n_23),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_23),
.B1(n_21),
.B2(n_19),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_43),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_19),
.B1(n_9),
.B2(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_92),
.B(n_91),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_4),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_57),
.B1(n_60),
.B2(n_51),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_4),
.B(n_9),
.C(n_11),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_101),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_46),
.A2(n_4),
.B1(n_12),
.B2(n_13),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_103),
.B(n_94),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_44),
.A2(n_13),
.B1(n_53),
.B2(n_51),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_115),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_109),
.Y(n_136)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_100),
.B(n_88),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_111),
.B(n_126),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_84),
.B(n_88),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_96),
.B1(n_102),
.B2(n_81),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_120),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_99),
.B1(n_92),
.B2(n_70),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_122),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_73),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_80),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_70),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_126),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_129),
.B1(n_128),
.B2(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_72),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_91),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_128),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_95),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_134),
.B1(n_132),
.B2(n_131),
.Y(n_154)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_151),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_140),
.A2(n_153),
.B(n_133),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_81),
.B1(n_102),
.B2(n_67),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_142),
.A2(n_146),
.B1(n_130),
.B2(n_135),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_67),
.B1(n_107),
.B2(n_111),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_156),
.B1(n_109),
.B2(n_133),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_105),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_127),
.B(n_107),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_144),
.B(n_149),
.C(n_148),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_115),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_164),
.B1(n_168),
.B2(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_113),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_172),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_148),
.B(n_142),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

AO221x1_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_166),
.B1(n_169),
.B2(n_141),
.C(n_149),
.Y(n_183)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_150),
.B1(n_156),
.B2(n_146),
.Y(n_168)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_173),
.B(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_147),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_156),
.Y(n_173)
);

NOR4xp25_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_157),
.C(n_152),
.D(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_162),
.B(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_174),
.B(n_154),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_181),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_183),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_155),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_171),
.B1(n_161),
.B2(n_175),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_159),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_165),
.C(n_184),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_189),
.B1(n_169),
.B2(n_166),
.Y(n_194)
);

OAI22x1_ASAP7_75t_SL g189 ( 
.A1(n_168),
.A2(n_139),
.B1(n_145),
.B2(n_144),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_194),
.A2(n_197),
.B1(n_188),
.B2(n_186),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_180),
.Y(n_201)
);

XOR2x2_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_165),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_188),
.B1(n_177),
.B2(n_181),
.Y(n_197)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_183),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_198),
.A2(n_201),
.B(n_176),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_200),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_192),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_180),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_203),
.A2(n_193),
.B(n_182),
.Y(n_206)
);

OAI221xp5_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_190),
.B1(n_197),
.B2(n_185),
.C(n_191),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_178),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_206),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_207),
.B(n_208),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_182),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_206),
.C(n_204),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_210),
.Y(n_212)
);


endmodule