module real_aes_7081_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g154 ( .A1(n_0), .A2(n_155), .B(n_156), .C(n_160), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_1), .B(n_149), .Y(n_162) );
INVx1_ASAP7_75t_L g106 ( .A(n_2), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_3), .B(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_4), .A2(n_143), .B(n_440), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_5), .A2(n_123), .B(n_140), .C(n_484), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_6), .A2(n_143), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_7), .B(n_149), .Y(n_446) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_8), .A2(n_115), .B(n_237), .Y(n_236) );
AND2x6_ASAP7_75t_L g140 ( .A(n_9), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_10), .A2(n_123), .B(n_140), .C(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g537 ( .A(n_11), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_12), .B(n_38), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_13), .B(n_159), .Y(n_486) );
INVx1_ASAP7_75t_L g120 ( .A(n_14), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_15), .B(n_134), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_16), .A2(n_135), .B(n_495), .C(n_497), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_17), .B(n_149), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_18), .B(n_177), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_19), .A2(n_123), .B(n_169), .C(n_176), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_20), .A2(n_158), .B(n_211), .C(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_21), .B(n_159), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_22), .B(n_159), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_23), .Y(n_464) );
INVx1_ASAP7_75t_L g434 ( .A(n_24), .Y(n_434) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_25), .A2(n_123), .B(n_176), .C(n_240), .Y(n_239) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_26), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_27), .Y(n_482) );
INVx1_ASAP7_75t_L g458 ( .A(n_28), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_29), .A2(n_143), .B(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g125 ( .A(n_30), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_31), .A2(n_138), .B(n_192), .C(n_193), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_32), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_33), .A2(n_158), .B(n_443), .C(n_445), .Y(n_442) );
INVxp67_ASAP7_75t_L g459 ( .A(n_34), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_35), .B(n_242), .Y(n_241) );
CKINVDCx14_ASAP7_75t_R g441 ( .A(n_36), .Y(n_441) );
A2O1A1Ixp33_ASAP7_75t_L g432 ( .A1(n_37), .A2(n_123), .B(n_176), .C(n_433), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_39), .A2(n_160), .B(n_535), .C(n_536), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_40), .B(n_167), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_41), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_42), .B(n_134), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_43), .B(n_143), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_44), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_45), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_46), .A2(n_138), .B(n_192), .C(n_220), .Y(n_219) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_47), .A2(n_66), .B1(n_101), .B2(n_684), .C1(n_688), .C2(n_689), .Y(n_100) );
INVx1_ASAP7_75t_L g157 ( .A(n_48), .Y(n_157) );
INVx1_ASAP7_75t_L g221 ( .A(n_49), .Y(n_221) );
INVx1_ASAP7_75t_L g502 ( .A(n_50), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_51), .B(n_143), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_52), .Y(n_181) );
CKINVDCx14_ASAP7_75t_R g533 ( .A(n_53), .Y(n_533) );
INVx1_ASAP7_75t_L g141 ( .A(n_54), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_55), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_56), .B(n_149), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_57), .A2(n_130), .B(n_175), .C(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g119 ( .A(n_58), .Y(n_119) );
INVx1_ASAP7_75t_SL g444 ( .A(n_59), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_60), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_61), .B(n_134), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_62), .B(n_149), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_63), .B(n_135), .Y(n_208) );
INVx1_ASAP7_75t_L g467 ( .A(n_64), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g152 ( .A(n_65), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_66), .Y(n_688) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_67), .A2(n_99), .B1(n_691), .B2(n_700), .C1(n_711), .C2(n_717), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g702 ( .A1(n_67), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_67), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_68), .B(n_171), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g122 ( .A1(n_69), .A2(n_123), .B(n_128), .C(n_138), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_70), .Y(n_230) );
INVx1_ASAP7_75t_L g695 ( .A(n_71), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_72), .A2(n_143), .B(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_73), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_74), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_75), .A2(n_143), .B(n_492), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_76), .A2(n_167), .B(n_454), .Y(n_453) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_77), .Y(n_431) );
INVx1_ASAP7_75t_L g493 ( .A(n_78), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_79), .B(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_80), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_81), .A2(n_143), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g496 ( .A(n_82), .Y(n_496) );
INVx2_ASAP7_75t_L g117 ( .A(n_83), .Y(n_117) );
INVx1_ASAP7_75t_L g485 ( .A(n_84), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_85), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_86), .B(n_159), .Y(n_209) );
OR2x2_ASAP7_75t_L g104 ( .A(n_87), .B(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g421 ( .A(n_87), .Y(n_421) );
OR2x2_ASAP7_75t_L g699 ( .A(n_87), .B(n_690), .Y(n_699) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_88), .A2(n_123), .B(n_138), .C(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_89), .B(n_143), .Y(n_190) );
INVx1_ASAP7_75t_L g194 ( .A(n_90), .Y(n_194) );
INVxp67_ASAP7_75t_L g233 ( .A(n_91), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_92), .B(n_115), .Y(n_538) );
INVx1_ASAP7_75t_L g129 ( .A(n_93), .Y(n_129) );
INVx1_ASAP7_75t_L g204 ( .A(n_94), .Y(n_204) );
INVx2_ASAP7_75t_L g505 ( .A(n_95), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_96), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g223 ( .A(n_97), .B(n_179), .Y(n_223) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI22xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_108), .B1(n_418), .B2(n_422), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g686 ( .A(n_103), .Y(n_686) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OR2x2_ASAP7_75t_L g420 ( .A(n_105), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g690 ( .A(n_105), .Y(n_690) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g685 ( .A(n_108), .Y(n_685) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_108), .Y(n_703) );
OR3x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_326), .C(n_375), .Y(n_108) );
NAND5xp2_ASAP7_75t_L g109 ( .A(n_110), .B(n_260), .C(n_289), .D(n_297), .E(n_312), .Y(n_109) );
O2A1O1Ixp33_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_183), .B(n_199), .C(n_244), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_163), .Y(n_111) );
AND2x2_ASAP7_75t_L g255 ( .A(n_112), .B(n_252), .Y(n_255) );
AND2x2_ASAP7_75t_L g288 ( .A(n_112), .B(n_164), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_112), .B(n_187), .Y(n_381) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_148), .Y(n_112) );
INVx2_ASAP7_75t_L g186 ( .A(n_113), .Y(n_186) );
BUFx2_ASAP7_75t_L g355 ( .A(n_113), .Y(n_355) );
AO21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_121), .B(n_146), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_114), .B(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g149 ( .A(n_114), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_114), .B(n_198), .Y(n_197) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_114), .A2(n_203), .B(n_213), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_114), .B(n_437), .Y(n_436) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_114), .A2(n_463), .B(n_470), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_114), .B(n_488), .Y(n_487) );
INVx4_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_115), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_115), .A2(n_238), .B(n_239), .Y(n_237) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g215 ( .A(n_116), .Y(n_215) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
AND2x2_ASAP7_75t_SL g179 ( .A(n_117), .B(n_118), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_142), .Y(n_121) );
INVx5_ASAP7_75t_L g153 ( .A(n_123), .Y(n_153) );
AND2x6_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_124), .Y(n_137) );
BUFx3_ASAP7_75t_L g161 ( .A(n_124), .Y(n_161) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g145 ( .A(n_125), .Y(n_145) );
INVx1_ASAP7_75t_L g212 ( .A(n_125), .Y(n_212) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_127), .Y(n_132) );
INVx3_ASAP7_75t_L g135 ( .A(n_127), .Y(n_135) );
AND2x2_ASAP7_75t_L g144 ( .A(n_127), .B(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_127), .Y(n_159) );
INVx1_ASAP7_75t_L g242 ( .A(n_127), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B(n_133), .C(n_136), .Y(n_128) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp33_ASAP7_75t_L g457 ( .A1(n_131), .A2(n_134), .B1(n_458), .B2(n_459), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_131), .B(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_131), .B(n_505), .Y(n_504) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
INVx2_ASAP7_75t_L g155 ( .A(n_134), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_134), .B(n_233), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g433 ( .A1(n_134), .A2(n_174), .B(n_434), .C(n_435), .Y(n_433) );
INVx5_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_135), .B(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx3_ASAP7_75t_L g445 ( .A(n_137), .Y(n_445) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
O2A1O1Ixp33_ASAP7_75t_SL g151 ( .A1(n_139), .A2(n_152), .B(n_153), .C(n_154), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_139), .A2(n_153), .B(n_230), .C(n_231), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g440 ( .A1(n_139), .A2(n_153), .B(n_441), .C(n_442), .Y(n_440) );
O2A1O1Ixp33_ASAP7_75t_SL g454 ( .A1(n_139), .A2(n_153), .B(n_455), .C(n_456), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_SL g492 ( .A1(n_139), .A2(n_153), .B(n_493), .C(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g501 ( .A1(n_139), .A2(n_153), .B(n_502), .C(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_139), .A2(n_153), .B(n_533), .C(n_534), .Y(n_532) );
INVx4_ASAP7_75t_SL g139 ( .A(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g143 ( .A(n_140), .B(n_144), .Y(n_143) );
BUFx3_ASAP7_75t_L g176 ( .A(n_140), .Y(n_176) );
NAND2x1p5_ASAP7_75t_L g205 ( .A(n_140), .B(n_144), .Y(n_205) );
BUFx2_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
INVx1_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
AND2x2_ASAP7_75t_L g163 ( .A(n_148), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g253 ( .A(n_148), .Y(n_253) );
AND2x2_ASAP7_75t_L g339 ( .A(n_148), .B(n_252), .Y(n_339) );
AND2x2_ASAP7_75t_L g394 ( .A(n_148), .B(n_186), .Y(n_394) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_162), .Y(n_148) );
INVx2_ASAP7_75t_L g192 ( .A(n_153), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_158), .B(n_444), .Y(n_443) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g535 ( .A(n_159), .Y(n_535) );
INVx2_ASAP7_75t_L g469 ( .A(n_160), .Y(n_469) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_161), .Y(n_196) );
INVx1_ASAP7_75t_L g497 ( .A(n_161), .Y(n_497) );
INVx1_ASAP7_75t_L g311 ( .A(n_163), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_163), .B(n_187), .Y(n_358) );
INVx5_ASAP7_75t_L g252 ( .A(n_164), .Y(n_252) );
AND2x4_ASAP7_75t_L g273 ( .A(n_164), .B(n_253), .Y(n_273) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_164), .Y(n_295) );
AND2x2_ASAP7_75t_L g370 ( .A(n_164), .B(n_355), .Y(n_370) );
AND2x2_ASAP7_75t_L g373 ( .A(n_164), .B(n_188), .Y(n_373) );
OR2x6_ASAP7_75t_L g164 ( .A(n_165), .B(n_180), .Y(n_164) );
AOI21xp5_ASAP7_75t_SL g165 ( .A1(n_166), .A2(n_168), .B(n_177), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_172), .B(n_174), .Y(n_169) );
INVx2_ASAP7_75t_L g173 ( .A(n_171), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_173), .A2(n_194), .B(n_195), .C(n_196), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_173), .A2(n_196), .B(n_221), .C(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_173), .A2(n_467), .B(n_468), .C(n_469), .Y(n_466) );
O2A1O1Ixp5_ASAP7_75t_L g484 ( .A1(n_173), .A2(n_469), .B(n_485), .C(n_486), .Y(n_484) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_175), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_178), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g182 ( .A(n_179), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_179), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_179), .A2(n_218), .B(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g430 ( .A1(n_179), .A2(n_205), .B(n_431), .C(n_432), .Y(n_430) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_179), .A2(n_531), .B(n_538), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_182), .A2(n_481), .B(n_487), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_183), .B(n_253), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_183), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_187), .Y(n_184) );
AND2x2_ASAP7_75t_L g278 ( .A(n_185), .B(n_253), .Y(n_278) );
AND2x2_ASAP7_75t_L g296 ( .A(n_185), .B(n_188), .Y(n_296) );
INVx1_ASAP7_75t_L g316 ( .A(n_185), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_185), .B(n_252), .Y(n_361) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_185), .Y(n_403) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_186), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_187), .B(n_251), .Y(n_250) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_187), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_187), .A2(n_248), .B(n_309), .C(n_311), .Y(n_308) );
AND2x2_ASAP7_75t_L g315 ( .A(n_187), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g324 ( .A(n_187), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g328 ( .A(n_187), .B(n_252), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_187), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g343 ( .A(n_187), .B(n_253), .Y(n_343) );
AND2x2_ASAP7_75t_L g393 ( .A(n_187), .B(n_394), .Y(n_393) );
INVx5_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
BUFx2_ASAP7_75t_L g257 ( .A(n_188), .Y(n_257) );
AND2x2_ASAP7_75t_L g298 ( .A(n_188), .B(n_251), .Y(n_298) );
AND2x2_ASAP7_75t_L g310 ( .A(n_188), .B(n_285), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_188), .B(n_339), .Y(n_357) );
OR2x6_ASAP7_75t_L g188 ( .A(n_189), .B(n_197), .Y(n_188) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_224), .Y(n_199) );
INVx1_ASAP7_75t_L g246 ( .A(n_200), .Y(n_246) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_216), .Y(n_200) );
OR2x2_ASAP7_75t_L g248 ( .A(n_201), .B(n_216), .Y(n_248) );
NAND3xp33_ASAP7_75t_L g254 ( .A(n_201), .B(n_255), .C(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_201), .B(n_226), .Y(n_265) );
OR2x2_ASAP7_75t_L g280 ( .A(n_201), .B(n_268), .Y(n_280) );
AND2x2_ASAP7_75t_L g286 ( .A(n_201), .B(n_235), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_201), .B(n_417), .Y(n_416) );
INVx5_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_202), .B(n_226), .Y(n_283) );
AND2x2_ASAP7_75t_L g322 ( .A(n_202), .B(n_236), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_202), .B(n_235), .Y(n_350) );
OR2x2_ASAP7_75t_L g353 ( .A(n_202), .B(n_235), .Y(n_353) );
OAI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_206), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_205), .A2(n_464), .B(n_465), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_205), .A2(n_482), .B(n_483), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_210), .A2(n_241), .B(n_243), .Y(n_240) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g452 ( .A(n_215), .Y(n_452) );
INVx5_ASAP7_75t_SL g268 ( .A(n_216), .Y(n_268) );
OR2x2_ASAP7_75t_L g274 ( .A(n_216), .B(n_225), .Y(n_274) );
AND2x2_ASAP7_75t_L g290 ( .A(n_216), .B(n_291), .Y(n_290) );
AOI321xp33_ASAP7_75t_L g297 ( .A1(n_216), .A2(n_298), .A3(n_299), .B1(n_300), .B2(n_306), .C(n_308), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_216), .B(n_224), .Y(n_307) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_216), .Y(n_320) );
OR2x2_ASAP7_75t_L g367 ( .A(n_216), .B(n_265), .Y(n_367) );
AND2x2_ASAP7_75t_L g389 ( .A(n_216), .B(n_286), .Y(n_389) );
AND2x2_ASAP7_75t_L g408 ( .A(n_216), .B(n_226), .Y(n_408) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_223), .Y(n_216) );
INVx1_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_235), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_226), .B(n_235), .Y(n_249) );
AND2x2_ASAP7_75t_L g258 ( .A(n_226), .B(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g285 ( .A(n_226), .Y(n_285) );
AND2x2_ASAP7_75t_L g291 ( .A(n_226), .B(n_286), .Y(n_291) );
INVxp67_ASAP7_75t_L g321 ( .A(n_226), .Y(n_321) );
OR2x2_ASAP7_75t_L g363 ( .A(n_226), .B(n_268), .Y(n_363) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_234), .Y(n_226) );
OA21x2_ASAP7_75t_L g438 ( .A1(n_227), .A2(n_439), .B(n_446), .Y(n_438) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_227), .A2(n_491), .B(n_498), .Y(n_490) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_227), .A2(n_500), .B(n_506), .Y(n_499) );
OR2x2_ASAP7_75t_L g245 ( .A(n_235), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_SL g259 ( .A(n_235), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_235), .B(n_248), .Y(n_292) );
AND2x2_ASAP7_75t_L g341 ( .A(n_235), .B(n_285), .Y(n_341) );
AND2x2_ASAP7_75t_L g379 ( .A(n_235), .B(n_268), .Y(n_379) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_236), .B(n_268), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_247), .B(n_250), .C(n_254), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_245), .A2(n_247), .B1(n_372), .B2(n_374), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_247), .A2(n_270), .B1(n_325), .B2(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
INVx1_ASAP7_75t_SL g399 ( .A(n_248), .Y(n_399) );
INVx1_ASAP7_75t_SL g299 ( .A(n_249), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_251), .B(n_271), .Y(n_301) );
AOI222xp33_ASAP7_75t_L g312 ( .A1(n_251), .A2(n_292), .B1(n_299), .B2(n_313), .C1(n_317), .C2(n_323), .Y(n_312) );
AND2x2_ASAP7_75t_L g402 ( .A(n_251), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx2_ASAP7_75t_L g277 ( .A(n_252), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_252), .B(n_272), .Y(n_347) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_252), .Y(n_384) );
AND2x2_ASAP7_75t_L g387 ( .A(n_252), .B(n_296), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_252), .B(n_403), .Y(n_413) );
INVx1_ASAP7_75t_L g304 ( .A(n_253), .Y(n_304) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_253), .Y(n_332) );
O2A1O1Ixp33_ASAP7_75t_L g395 ( .A1(n_255), .A2(n_396), .B(n_397), .C(n_400), .Y(n_395) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NAND3xp33_ASAP7_75t_L g318 ( .A(n_257), .B(n_319), .C(n_322), .Y(n_318) );
OR2x2_ASAP7_75t_L g346 ( .A(n_257), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_257), .B(n_273), .Y(n_374) );
OR2x2_ASAP7_75t_L g279 ( .A(n_259), .B(n_280), .Y(n_279) );
AOI211xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_263), .B(n_269), .C(n_281), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_262), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g368 ( .A(n_263), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_264), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g282 ( .A(n_267), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_268), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g336 ( .A(n_268), .B(n_286), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_268), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_268), .B(n_285), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_274), .B1(n_275), .B2(n_279), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_271), .B(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_273), .B(n_315), .Y(n_314) );
OAI221xp5_ASAP7_75t_SL g337 ( .A1(n_274), .A2(n_338), .B1(n_340), .B2(n_342), .C(n_344), .Y(n_337) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g392 ( .A(n_277), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g405 ( .A(n_277), .B(n_394), .Y(n_405) );
INVx1_ASAP7_75t_L g325 ( .A(n_278), .Y(n_325) );
INVx1_ASAP7_75t_L g396 ( .A(n_279), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_280), .A2(n_363), .B(n_386), .Y(n_385) );
AOI21xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_284), .B(n_287), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OAI21xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_292), .B(n_293), .Y(n_289) );
INVx1_ASAP7_75t_L g329 ( .A(n_290), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_291), .A2(n_377), .B1(n_380), .B2(n_382), .C(n_385), .Y(n_376) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_299), .A2(n_389), .B1(n_390), .B2(n_392), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g365 ( .A(n_301), .Y(n_365) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NOR2xp67_ASAP7_75t_SL g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AND2x2_ASAP7_75t_L g369 ( .A(n_305), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g334 ( .A(n_310), .Y(n_334) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_315), .B(n_339), .Y(n_391) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_321), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g407 ( .A(n_322), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g414 ( .A(n_322), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI211xp5_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_329), .B(n_330), .C(n_364), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI211xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_337), .C(n_356), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g417 ( .A(n_341), .Y(n_417) );
AND2x2_ASAP7_75t_L g354 ( .A(n_343), .B(n_355), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_348), .B1(n_352), .B2(n_354), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
OR2x2_ASAP7_75t_L g362 ( .A(n_350), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g415 ( .A(n_351), .Y(n_415) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI31xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .A3(n_359), .B(n_362), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI211xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B(n_368), .C(n_371), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
CKINVDCx16_ASAP7_75t_R g372 ( .A(n_373), .Y(n_372) );
NAND5xp2_ASAP7_75t_L g375 ( .A(n_376), .B(n_388), .C(n_395), .D(n_409), .E(n_412), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_387), .A2(n_413), .B1(n_414), .B2(n_416), .Y(n_412) );
INVx1_ASAP7_75t_SL g411 ( .A(n_389), .Y(n_411) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_404), .B(n_406), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI22xp5_ASAP7_75t_SL g684 ( .A1(n_420), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_684) );
NOR2x2_ASAP7_75t_L g689 ( .A(n_421), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g687 ( .A(n_422), .Y(n_687) );
OR3x1_ASAP7_75t_L g422 ( .A(n_423), .B(n_595), .C(n_642), .Y(n_422) );
NAND3xp33_ASAP7_75t_SL g423 ( .A(n_424), .B(n_541), .C(n_566), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_479), .B1(n_507), .B2(n_510), .C(n_518), .Y(n_424) );
OAI21xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_447), .B(n_472), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_427), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_427), .B(n_523), .Y(n_639) );
AND2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_438), .Y(n_427) );
AND2x2_ASAP7_75t_L g509 ( .A(n_428), .B(n_478), .Y(n_509) );
AND2x2_ASAP7_75t_L g559 ( .A(n_428), .B(n_477), .Y(n_559) );
AND2x2_ASAP7_75t_L g580 ( .A(n_428), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g585 ( .A(n_428), .B(n_552), .Y(n_585) );
OR2x2_ASAP7_75t_L g593 ( .A(n_428), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g665 ( .A(n_428), .B(n_461), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_428), .B(n_614), .Y(n_679) );
INVx3_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g524 ( .A(n_429), .B(n_438), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_429), .B(n_461), .Y(n_525) );
AND2x4_ASAP7_75t_L g547 ( .A(n_429), .B(n_478), .Y(n_547) );
AND2x2_ASAP7_75t_L g577 ( .A(n_429), .B(n_449), .Y(n_577) );
AND2x2_ASAP7_75t_L g586 ( .A(n_429), .B(n_576), .Y(n_586) );
AND2x2_ASAP7_75t_L g602 ( .A(n_429), .B(n_462), .Y(n_602) );
OR2x2_ASAP7_75t_L g611 ( .A(n_429), .B(n_594), .Y(n_611) );
AND2x2_ASAP7_75t_L g617 ( .A(n_429), .B(n_552), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_429), .B(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g631 ( .A(n_429), .B(n_474), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_429), .B(n_520), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_429), .B(n_581), .Y(n_670) );
OR2x6_ASAP7_75t_L g429 ( .A(n_430), .B(n_436), .Y(n_429) );
INVx2_ASAP7_75t_L g478 ( .A(n_438), .Y(n_478) );
AND2x2_ASAP7_75t_L g576 ( .A(n_438), .B(n_461), .Y(n_576) );
AND2x2_ASAP7_75t_L g581 ( .A(n_438), .B(n_462), .Y(n_581) );
INVx1_ASAP7_75t_L g637 ( .A(n_438), .Y(n_637) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g546 ( .A(n_448), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_461), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_449), .B(n_509), .Y(n_508) );
BUFx3_ASAP7_75t_L g523 ( .A(n_449), .Y(n_523) );
OR2x2_ASAP7_75t_L g594 ( .A(n_449), .B(n_461), .Y(n_594) );
OR2x2_ASAP7_75t_L g655 ( .A(n_449), .B(n_562), .Y(n_655) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_453), .B(n_460), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_451), .A2(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g475 ( .A(n_453), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_460), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_461), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g614 ( .A(n_461), .B(n_474), .Y(n_614) );
INVx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
BUFx2_ASAP7_75t_L g553 ( .A(n_462), .Y(n_553) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_473), .A2(n_659), .B1(n_663), .B2(n_666), .C(n_667), .Y(n_658) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_477), .Y(n_473) );
INVx1_ASAP7_75t_SL g521 ( .A(n_474), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_474), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g653 ( .A(n_474), .B(n_509), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_477), .B(n_523), .Y(n_645) );
AND2x2_ASAP7_75t_L g552 ( .A(n_478), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_SL g556 ( .A(n_479), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_479), .B(n_562), .Y(n_592) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_489), .Y(n_479) );
AND2x2_ASAP7_75t_L g517 ( .A(n_480), .B(n_490), .Y(n_517) );
INVx4_ASAP7_75t_L g529 ( .A(n_480), .Y(n_529) );
BUFx3_ASAP7_75t_L g572 ( .A(n_480), .Y(n_572) );
AND3x2_ASAP7_75t_L g587 ( .A(n_480), .B(n_588), .C(n_589), .Y(n_587) );
AND2x2_ASAP7_75t_L g669 ( .A(n_489), .B(n_583), .Y(n_669) );
AND2x2_ASAP7_75t_L g677 ( .A(n_489), .B(n_562), .Y(n_677) );
INVx1_ASAP7_75t_SL g682 ( .A(n_489), .Y(n_682) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
INVx1_ASAP7_75t_SL g540 ( .A(n_490), .Y(n_540) );
AND2x2_ASAP7_75t_L g563 ( .A(n_490), .B(n_529), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_490), .B(n_513), .Y(n_565) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_490), .Y(n_605) );
OR2x2_ASAP7_75t_L g610 ( .A(n_490), .B(n_529), .Y(n_610) );
INVx2_ASAP7_75t_L g515 ( .A(n_499), .Y(n_515) );
AND2x2_ASAP7_75t_L g550 ( .A(n_499), .B(n_530), .Y(n_550) );
OR2x2_ASAP7_75t_L g570 ( .A(n_499), .B(n_530), .Y(n_570) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_499), .Y(n_590) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
AOI21xp33_ASAP7_75t_L g640 ( .A1(n_508), .A2(n_549), .B(n_641), .Y(n_640) );
AOI322xp5_ASAP7_75t_L g676 ( .A1(n_510), .A2(n_520), .A3(n_547), .B1(n_677), .B2(n_678), .C1(n_680), .C2(n_683), .Y(n_676) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_516), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_512), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_513), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g539 ( .A(n_514), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g607 ( .A(n_515), .B(n_529), .Y(n_607) );
AND2x2_ASAP7_75t_L g674 ( .A(n_515), .B(n_530), .Y(n_674) );
INVx1_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g615 ( .A(n_517), .B(n_569), .Y(n_615) );
AOI31xp33_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_522), .A3(n_525), .B(n_526), .Y(n_518) );
AND2x2_ASAP7_75t_L g574 ( .A(n_520), .B(n_552), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_520), .B(n_544), .Y(n_656) );
AND2x2_ASAP7_75t_L g675 ( .A(n_520), .B(n_580), .Y(n_675) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_523), .B(n_552), .Y(n_564) );
NAND2x1p5_ASAP7_75t_L g598 ( .A(n_523), .B(n_581), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_523), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_523), .B(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_524), .B(n_581), .Y(n_613) );
INVx1_ASAP7_75t_L g657 ( .A(n_524), .Y(n_657) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_539), .Y(n_527) );
INVxp67_ASAP7_75t_L g609 ( .A(n_528), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_529), .B(n_540), .Y(n_545) );
INVx1_ASAP7_75t_L g651 ( .A(n_529), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_529), .B(n_628), .Y(n_662) );
BUFx3_ASAP7_75t_L g562 ( .A(n_530), .Y(n_562) );
AND2x2_ASAP7_75t_L g588 ( .A(n_530), .B(n_540), .Y(n_588) );
INVx2_ASAP7_75t_L g628 ( .A(n_530), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_539), .B(n_661), .Y(n_660) );
AOI211xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_546), .B(n_548), .C(n_557), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AOI21xp33_ASAP7_75t_L g591 ( .A1(n_543), .A2(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_544), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_544), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g624 ( .A(n_545), .B(n_570), .Y(n_624) );
INVx3_ASAP7_75t_L g555 ( .A(n_547), .Y(n_555) );
OAI22xp5_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_551), .B1(n_554), .B2(n_556), .Y(n_548) );
OAI21xp5_ASAP7_75t_SL g573 ( .A1(n_550), .A2(n_574), .B(n_575), .Y(n_573) );
AND2x2_ASAP7_75t_L g599 ( .A(n_550), .B(n_563), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_550), .B(n_651), .Y(n_650) );
INVxp67_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g554 ( .A(n_553), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g623 ( .A(n_553), .Y(n_623) );
OAI21xp5_ASAP7_75t_SL g567 ( .A1(n_554), .A2(n_568), .B(n_573), .Y(n_567) );
OAI22xp33_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_560), .B1(n_564), .B2(n_565), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_559), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g583 ( .A(n_562), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_562), .B(n_605), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_578), .C(n_591), .Y(n_566) );
OAI22xp5_ASAP7_75t_SL g633 ( .A1(n_568), .A2(n_634), .B1(n_638), .B2(n_639), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g638 ( .A(n_570), .B(n_571), .Y(n_638) );
AND2x2_ASAP7_75t_L g646 ( .A(n_571), .B(n_627), .Y(n_646) );
CKINVDCx16_ASAP7_75t_R g571 ( .A(n_572), .Y(n_571) );
O2A1O1Ixp33_ASAP7_75t_SL g654 ( .A1(n_572), .A2(n_655), .B(n_656), .C(n_657), .Y(n_654) );
OR2x2_ASAP7_75t_L g681 ( .A(n_572), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
OAI21xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .B(n_584), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
O2A1O1Ixp33_ASAP7_75t_L g616 ( .A1(n_580), .A2(n_617), .B(n_618), .C(n_621), .Y(n_616) );
OAI21xp33_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_586), .B(n_587), .Y(n_584) );
AND2x2_ASAP7_75t_L g649 ( .A(n_588), .B(n_607), .Y(n_649) );
INVxp67_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g627 ( .A(n_590), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g632 ( .A(n_592), .Y(n_632) );
NAND3xp33_ASAP7_75t_SL g595 ( .A(n_596), .B(n_616), .C(n_629), .Y(n_595) );
AOI211xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_599), .B(n_600), .C(n_608), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_L g666 ( .A(n_603), .Y(n_666) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx1_ASAP7_75t_L g626 ( .A(n_605), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_605), .B(n_674), .Y(n_673) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_611), .C(n_612), .Y(n_608) );
INVx2_ASAP7_75t_SL g620 ( .A(n_610), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_611), .A2(n_622), .B1(n_624), .B2(n_625), .Y(n_621) );
OAI21xp33_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_614), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B(n_633), .C(n_640), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVxp33_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g683 ( .A(n_637), .Y(n_683) );
NAND4xp25_ASAP7_75t_L g642 ( .A(n_643), .B(n_658), .C(n_671), .D(n_676), .Y(n_642) );
AOI211xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B(n_647), .C(n_654), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_650), .B(n_652), .Y(n_647) );
AOI21xp33_ASAP7_75t_L g667 ( .A1(n_648), .A2(n_668), .B(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_655), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_675), .Y(n_671) );
INVxp67_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_697), .Y(n_692) );
NOR2xp33_ASAP7_75t_SL g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_SL g716 ( .A(n_694), .Y(n_716) );
INVx1_ASAP7_75t_L g715 ( .A(n_696), .Y(n_715) );
OA21x2_ASAP7_75t_L g718 ( .A1(n_696), .A2(n_716), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_699), .Y(n_708) );
BUFx2_ASAP7_75t_L g719 ( .A(n_699), .Y(n_719) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_706), .B(n_709), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_703), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_708), .B(n_710), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_712), .Y(n_711) );
CKINVDCx6p67_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_718), .Y(n_717) );
endmodule