module fake_jpeg_30296_n_493 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_493);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_493;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_14),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_54),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_85),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_56),
.Y(n_127)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_61),
.B(n_71),
.Y(n_129)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_16),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_74),
.Y(n_122)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_15),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_79),
.B(n_94),
.Y(n_147)
);

BUFx16f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_80),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_82),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_14),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

BUFx16f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_93),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_91),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_39),
.B(n_14),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_40),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_97),
.Y(n_123)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_100),
.Y(n_124)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_101),
.Y(n_143)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_40),
.B(n_0),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_37),
.B1(n_33),
.B2(n_30),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_105),
.A2(n_106),
.B1(n_118),
.B2(n_130),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_37),
.B1(n_33),
.B2(n_41),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_37),
.B1(n_33),
.B2(n_41),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_45),
.B1(n_42),
.B2(n_48),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_91),
.A2(n_33),
.B1(n_41),
.B2(n_20),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_52),
.B(n_22),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_45),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_98),
.A2(n_41),
.B1(n_36),
.B2(n_34),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_153),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_58),
.A2(n_42),
.B1(n_36),
.B2(n_34),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_60),
.A2(n_28),
.B1(n_4),
.B2(n_5),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_89),
.B(n_28),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_159),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_63),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_64),
.A2(n_68),
.B1(n_72),
.B2(n_92),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_95),
.B1(n_87),
.B2(n_97),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_77),
.B(n_3),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_90),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_66),
.B(n_13),
.Y(n_159)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_162),
.B(n_164),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_163),
.B(n_166),
.Y(n_244)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_107),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_165),
.B(n_169),
.Y(n_235)
);

HAxp5_ASAP7_75t_SL g166 ( 
.A(n_156),
.B(n_80),
.CON(n_166),
.SN(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_96),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_182),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_168),
.A2(n_109),
.B1(n_113),
.B2(n_126),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_110),
.B(n_62),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_170),
.B(n_179),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_69),
.B(n_74),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_176),
.A2(n_113),
.B(n_102),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_124),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_147),
.B(n_50),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_180),
.B(n_190),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g181 ( 
.A(n_135),
.B(n_88),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_181),
.B(n_176),
.C(n_214),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_129),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_117),
.B(n_81),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_193),
.Y(n_224)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_78),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_188),
.B(n_194),
.Y(n_232)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_146),
.B(n_108),
.Y(n_190)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_120),
.B(n_5),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_125),
.B(n_56),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_125),
.B(n_133),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_195),
.B(n_214),
.Y(n_257)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_196),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_128),
.A2(n_65),
.B1(n_7),
.B2(n_8),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_109),
.B1(n_103),
.B2(n_151),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_6),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_201),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

AO22x1_ASAP7_75t_SL g200 ( 
.A1(n_133),
.A2(n_138),
.B1(n_160),
.B2(n_152),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_200),
.B(n_202),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_155),
.B(n_6),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_7),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_116),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_203),
.B(n_206),
.Y(n_243)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_204),
.Y(n_227)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_132),
.B(n_7),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_212),
.Y(n_247)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_208),
.Y(n_241)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_209),
.Y(n_249)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_102),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_123),
.B(n_7),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_123),
.B(n_8),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_181),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_182),
.A2(n_119),
.B(n_123),
.C(n_132),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_219),
.B(n_258),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_225),
.A2(n_177),
.B1(n_199),
.B2(n_209),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_210),
.A2(n_122),
.B1(n_121),
.B2(n_127),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_230),
.A2(n_238),
.B(n_253),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_210),
.A2(n_127),
.B1(n_140),
.B2(n_116),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_231),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_178),
.A2(n_122),
.B1(n_121),
.B2(n_151),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_167),
.B(n_172),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_242),
.C(n_215),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_181),
.A2(n_114),
.B1(n_140),
.B2(n_103),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_259),
.B1(n_191),
.B2(n_171),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_227),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_296),
.Y(n_307)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_262),
.A2(n_279),
.B1(n_290),
.B2(n_230),
.Y(n_310)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_263),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_224),
.B(n_175),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_264),
.B(n_284),
.Y(n_319)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_267),
.Y(n_316)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_268),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_289),
.B1(n_291),
.B2(n_294),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_270),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_195),
.C(n_191),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_287),
.C(n_242),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_166),
.B1(n_200),
.B2(n_187),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_272),
.A2(n_219),
.B1(n_225),
.B2(n_220),
.Y(n_312)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_189),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_277),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_227),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_SL g328 ( 
.A(n_275),
.B(n_223),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_235),
.B(n_174),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_244),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_278),
.B(n_292),
.Y(n_327)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_280),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_217),
.B(n_200),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_285),
.Y(n_317)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_283),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_233),
.B(n_173),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_205),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_236),
.B(n_185),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_293),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_240),
.B(n_161),
.C(n_196),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_254),
.A2(n_192),
.B1(n_208),
.B2(n_213),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_232),
.A2(n_183),
.B1(n_137),
.B2(n_204),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_232),
.A2(n_137),
.B1(n_10),
.B2(n_11),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_229),
.B(n_9),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_257),
.B(n_9),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_238),
.A2(n_137),
.B1(n_11),
.B2(n_12),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_247),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_216),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_10),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_234),
.B(n_10),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_234),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_299),
.B(n_304),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_253),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_300),
.A2(n_328),
.B(n_275),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_248),
.B1(n_259),
.B2(n_244),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_302),
.A2(n_262),
.B1(n_272),
.B2(n_287),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_267),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_305),
.B(n_274),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_260),
.B(n_258),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_306),
.B(n_314),
.C(n_326),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_310),
.A2(n_312),
.B1(n_291),
.B2(n_288),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_276),
.A2(n_244),
.B(n_243),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_311),
.A2(n_322),
.B(n_323),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_229),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_261),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_329),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_288),
.A2(n_228),
.B(n_220),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_294),
.A2(n_228),
.B1(n_245),
.B2(n_221),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_271),
.B(n_256),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_296),
.Y(n_332)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_334),
.A2(n_350),
.B1(n_359),
.B2(n_362),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_303),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_335),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_336),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_305),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_349),
.C(n_358),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_264),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_339),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_351),
.Y(n_366)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_301),
.Y(n_342)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_303),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_343),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_319),
.B(n_297),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_344),
.B(n_321),
.Y(n_388)
);

INVxp33_ASAP7_75t_SL g345 ( 
.A(n_316),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_345),
.Y(n_389)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_301),
.Y(n_346)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_346),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_306),
.B(n_293),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_347),
.B(n_327),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_277),
.Y(n_348)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_312),
.A2(n_269),
.B1(n_284),
.B2(n_285),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_298),
.A2(n_286),
.B1(n_283),
.B2(n_282),
.Y(n_351)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_315),
.Y(n_353)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_266),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_354),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_270),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_355),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_309),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_361),
.Y(n_367)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_309),
.Y(n_357)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_307),
.B(n_311),
.C(n_322),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_298),
.A2(n_280),
.B1(n_273),
.B2(n_268),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_265),
.Y(n_360)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_313),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_300),
.A2(n_270),
.B1(n_218),
.B2(n_249),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_360),
.B(n_300),
.Y(n_369)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_369),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_307),
.C(n_300),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_358),
.C(n_352),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_308),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_337),
.A2(n_300),
.B(n_323),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_377),
.B(n_336),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_321),
.Y(n_378)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_378),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_334),
.A2(n_302),
.B1(n_325),
.B2(n_324),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_382),
.A2(n_384),
.B1(n_318),
.B2(n_328),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_350),
.A2(n_313),
.B1(n_325),
.B2(n_324),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_362),
.B(n_337),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_385),
.Y(n_393)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_388),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_335),
.B(n_343),
.Y(n_390)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_390),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_391),
.B(n_409),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_349),
.C(n_352),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_392),
.B(n_399),
.C(n_400),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_376),
.A2(n_341),
.B1(n_351),
.B2(n_361),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_395),
.A2(n_406),
.B1(n_408),
.B2(n_363),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_397),
.A2(n_385),
.B(n_369),
.Y(n_417)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_367),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_407),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_368),
.B(n_347),
.C(n_332),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_340),
.C(n_359),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_333),
.C(n_357),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_401),
.B(n_404),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_379),
.A2(n_344),
.B1(n_356),
.B2(n_346),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_403),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_388),
.B(n_342),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_367),
.B(n_318),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_376),
.A2(n_331),
.B1(n_353),
.B2(n_308),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_390),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_410),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_365),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_411),
.B(n_413),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_331),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_414),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_249),
.C(n_263),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

OAI21xp33_ASAP7_75t_L g415 ( 
.A1(n_402),
.A2(n_363),
.B(n_372),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_418),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_423),
.Y(n_437)
);

MAJx2_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_392),
.C(n_399),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_398),
.A2(n_382),
.B1(n_385),
.B2(n_371),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_419),
.A2(n_406),
.B1(n_408),
.B2(n_405),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_393),
.A2(n_385),
.B(n_372),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_420),
.A2(n_426),
.B(n_370),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_393),
.A2(n_377),
.B(n_366),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_378),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_427),
.B(n_428),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_395),
.A2(n_366),
.B1(n_386),
.B2(n_375),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_409),
.B(n_375),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_429),
.B(n_364),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_386),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_433),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_400),
.C(n_401),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_435),
.B(n_441),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_440),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_420),
.A2(n_387),
.B(n_413),
.Y(n_438)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_438),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_424),
.B(n_394),
.C(n_396),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_364),
.C(n_389),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_443),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_389),
.C(n_381),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_430),
.A2(n_381),
.B1(n_370),
.B2(n_365),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_444),
.B(n_433),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_445),
.A2(n_417),
.B(n_422),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_380),
.C(n_315),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_447),
.B(n_431),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_416),
.B(n_380),
.Y(n_448)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_448),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_452),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_437),
.A2(n_430),
.B1(n_419),
.B2(n_425),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_450),
.A2(n_462),
.B1(n_426),
.B2(n_439),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_446),
.A2(n_421),
.B1(n_434),
.B2(n_425),
.Y(n_451)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_427),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_422),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_454),
.Y(n_467)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_439),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_447),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_457),
.A2(n_442),
.B(n_429),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_441),
.A2(n_421),
.B1(n_428),
.B2(n_423),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_460),
.A2(n_461),
.B(n_459),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_463),
.A2(n_468),
.B(n_473),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_465),
.B(n_466),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_458),
.B(n_435),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_469),
.B(n_470),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_449),
.A2(n_241),
.B1(n_218),
.B2(n_251),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_457),
.A2(n_251),
.B(n_252),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_471),
.A2(n_452),
.B(n_454),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_453),
.A2(n_222),
.B(n_246),
.Y(n_473)
);

A2O1A1O1Ixp25_ASAP7_75t_L g481 ( 
.A1(n_477),
.A2(n_472),
.B(n_467),
.C(n_471),
.D(n_466),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_468),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_478),
.B(n_479),
.C(n_450),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_464),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_462),
.Y(n_480)
);

NOR3xp33_ASAP7_75t_L g484 ( 
.A(n_480),
.B(n_455),
.C(n_218),
.Y(n_484)
);

OAI21x1_ASAP7_75t_L g486 ( 
.A1(n_481),
.A2(n_483),
.B(n_485),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_482),
.B(n_484),
.Y(n_487)
);

AOI21x1_ASAP7_75t_SL g483 ( 
.A1(n_476),
.A2(n_455),
.B(n_241),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_475),
.A2(n_237),
.B(n_246),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_482),
.A2(n_474),
.B(n_237),
.Y(n_488)
);

BUFx24_ASAP7_75t_SL g489 ( 
.A(n_488),
.Y(n_489)
);

AO221x1_ASAP7_75t_L g490 ( 
.A1(n_487),
.A2(n_137),
.B1(n_252),
.B2(n_13),
.C(n_11),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_486),
.C(n_12),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_491),
.B(n_489),
.C(n_12),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_492),
.Y(n_493)
);


endmodule