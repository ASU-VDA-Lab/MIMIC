module real_jpeg_894_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_249;
wire n_83;
wire n_78;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_164;
wire n_48;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_213;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_4),
.A2(n_57),
.B1(n_58),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_4),
.A2(n_34),
.B1(n_36),
.B2(n_70),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_70),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_70),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_7),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_7),
.B(n_29),
.C(n_42),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_7),
.A2(n_38),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_7),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_7),
.B(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_7),
.B(n_27),
.C(n_34),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_7),
.B(n_58),
.C(n_74),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_7),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_7),
.B(n_62),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_7),
.B(n_73),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_8),
.A2(n_57),
.B1(n_58),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_8),
.A2(n_34),
.B1(n_36),
.B2(n_95),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_95),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_95),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_249),
.Y(n_11)
);

OAI21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_238),
.B(n_248),
.Y(n_12)
);

AOI21x1_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_207),
.B(n_235),
.Y(n_13)
);

OAI21x1_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_186),
.B(n_206),
.Y(n_14)
);

AOI21x1_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_164),
.B(n_185),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_111),
.Y(n_16)
);

AOI21xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_97),
.B(n_110),
.Y(n_17)
);

NAND3xp33_ASAP7_75t_SL g111 ( 
.A(n_18),
.B(n_112),
.C(n_113),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_84),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_19),
.B(n_84),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_65),
.C(n_80),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_20),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_50),
.B2(n_64),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_21),
.A2(n_22),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_21),
.A2(n_22),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_39),
.B2(n_49),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_23),
.B(n_49),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_23),
.A2(n_24),
.B1(n_71),
.B2(n_72),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_23),
.A2(n_24),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_23),
.A2(n_72),
.B(n_83),
.C(n_155),
.Y(n_158)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_24),
.B(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_24),
.B(n_71),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_24),
.B(n_55),
.C(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_24),
.A2(n_198),
.B(n_202),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_24),
.B(n_198),
.Y(n_202)
);

AO21x2_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_33),
.B(n_37),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_25),
.A2(n_33),
.B1(n_37),
.B2(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_25),
.A2(n_33),
.B1(n_218),
.B2(n_231),
.Y(n_230)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_25),
.A2(n_33),
.B(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_27),
.Y(n_32)
);

OA22x2_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_29),
.B1(n_42),
.B2(n_46),
.Y(n_47)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_29),
.B(n_123),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_33),
.Y(n_140)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_34),
.A2(n_36),
.B1(n_74),
.B2(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_34),
.B(n_134),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_39),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_39),
.A2(n_49),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_39),
.A2(n_49),
.B1(n_174),
.B2(n_181),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_39),
.A2(n_49),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_39),
.A2(n_49),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_39),
.A2(n_49),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_39),
.B(n_216),
.C(n_217),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_39),
.B(n_227),
.C(n_233),
.Y(n_247)
);

AO21x2_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_47),
.B(n_48),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_40),
.A2(n_47),
.B1(n_48),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_40),
.A2(n_47),
.B1(n_246),
.B2(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_47),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_53),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

AOI211xp5_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_72),
.B(n_82),
.C(n_83),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_49),
.A2(n_181),
.B(n_192),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_49),
.B(n_215),
.C(n_230),
.Y(n_241)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_54),
.A2(n_55),
.B1(n_108),
.B2(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_54),
.B(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_54),
.A2(n_55),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_54),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_54),
.A2(n_55),
.B1(n_121),
.B2(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_55),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_55),
.B(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_55),
.B(n_71),
.C(n_139),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_61),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_62),
.Y(n_63)
);

AO22x1_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_58),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_58),
.B(n_145),
.Y(n_144)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_61),
.B(n_94),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_80),
.B1(n_81),
.B2(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_72),
.B2(n_79),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_72),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_72),
.B1(n_93),
.B2(n_96),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_116),
.C(n_120),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_71),
.A2(n_72),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_71),
.A2(n_72),
.B1(n_132),
.B2(n_133),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_71),
.A2(n_72),
.B1(n_120),
.B2(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_72),
.B(n_93),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B(n_78),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_73),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_73),
.A2(n_76),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_76),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_78),
.Y(n_178)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_85),
.B(n_89),
.C(n_92),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_86),
.A2(n_87),
.B(n_90),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_86),
.A2(n_87),
.B(n_171),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_93),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_101),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.C(n_107),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_103),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_104),
.A2(n_105),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_127),
.B(n_163),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_124),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_124),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_157),
.B(n_162),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_151),
.B(n_156),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_141),
.B(n_150),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_135),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_153),
.Y(n_156)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_159),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_165),
.B(n_166),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_184),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_173),
.B1(n_182),
.B2(n_183),
.Y(n_169)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_182),
.C(n_184),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_181),
.Y(n_173)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_174),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_176),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_177),
.A2(n_180),
.B(n_201),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_188),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_188)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_196),
.B2(n_197),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_196),
.C(n_203),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_211),
.B1(n_212),
.B2(n_220),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_223),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_222),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_222),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_221),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_220),
.C(n_221),
.Y(n_234)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_219),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_215),
.A2(n_216),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_223),
.A2(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_234),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_234),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_233),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_230),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_247),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_239),
.B(n_247),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_244),
.C(n_245),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_253),
.Y(n_255)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);


endmodule