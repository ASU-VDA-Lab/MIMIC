module fake_ibex_1366_n_1223 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_195, n_163, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1223);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1223;

wire n_1084;
wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1148;
wire n_1011;
wire n_992;
wire n_1104;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_1196;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_1182;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_1143;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_510;
wire n_845;
wire n_972;
wire n_981;
wire n_1100;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_1080;
wire n_1162;
wire n_1199;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1044;
wire n_1018;
wire n_1106;
wire n_1129;
wire n_449;
wire n_1138;
wire n_547;
wire n_1134;
wire n_727;
wire n_1131;
wire n_1077;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_1174;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1217;
wire n_1045;
wire n_753;
wire n_645;
wire n_747;
wire n_500;
wire n_963;
wire n_1147;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_1189;
wire n_531;
wire n_647;
wire n_1187;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_280;
wire n_375;
wire n_340;
wire n_317;
wire n_708;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_1218;
wire n_1166;
wire n_1181;
wire n_1140;
wire n_326;
wire n_327;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_1144;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_1203;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_1109;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_671;
wire n_228;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_1193;
wire n_458;
wire n_244;
wire n_1053;
wire n_1112;
wire n_1207;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_1172;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_1169;
wire n_386;
wire n_549;
wire n_224;
wire n_1210;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_1201;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_1103;
wire n_1161;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1177;
wire n_1057;
wire n_1068;
wire n_496;
wire n_301;
wire n_325;
wire n_617;
wire n_434;
wire n_1184;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_1195;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_1141;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_1075;
wire n_719;
wire n_370;
wire n_431;
wire n_614;
wire n_1197;
wire n_574;
wire n_1168;
wire n_289;
wire n_716;
wire n_865;
wire n_1130;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_1179;
wire n_1192;
wire n_933;
wire n_1081;
wire n_215;
wire n_1153;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_1155;
wire n_750;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1191;
wire n_1101;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_1133;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_1178;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_1211;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_1214;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_1137;
wire n_1082;
wire n_222;
wire n_660;
wire n_1213;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_1070;
wire n_454;
wire n_980;
wire n_1074;
wire n_777;
wire n_1200;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_1180;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_1220;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_1028;
wire n_1012;
wire n_993;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_1183;
wire n_253;
wire n_208;
wire n_234;
wire n_1204;
wire n_300;
wire n_1151;
wire n_1135;
wire n_973;
wire n_1146;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_999;
wire n_1092;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_648;
wire n_229;
wire n_209;
wire n_472;
wire n_571;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1142;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_1215;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1173;
wire n_1069;
wire n_573;
wire n_1208;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_433;
wire n_262;
wire n_439;
wire n_299;
wire n_704;
wire n_949;
wire n_1007;
wire n_1171;
wire n_1126;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_1115;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_1219;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_1170;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_1049;
wire n_1086;
wire n_763;
wire n_1158;
wire n_745;
wire n_329;
wire n_1149;
wire n_447;
wire n_1176;
wire n_940;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_788;
wire n_1202;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_1160;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_1216;
wire n_1222;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_1033;
wire n_1118;
wire n_692;
wire n_627;
wire n_990;
wire n_1198;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_1167;
wire n_653;
wire n_1205;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_1059;
wire n_1019;
wire n_902;
wire n_332;
wire n_799;
wire n_1190;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_951;
wire n_272;
wire n_881;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_223;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1209;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_285;
wire n_247;
wire n_379;
wire n_288;
wire n_1128;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_807;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_1145;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_1164;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_866;
wire n_958;
wire n_1175;
wire n_485;
wire n_1139;
wire n_870;
wire n_1221;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_1212;
wire n_461;
wire n_575;
wire n_313;
wire n_1159;
wire n_1119;
wire n_903;
wire n_1154;
wire n_519;
wire n_345;
wire n_408;
wire n_1095;
wire n_361;
wire n_1085;
wire n_455;
wire n_1136;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_528;
wire n_1005;
wire n_1102;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_1194;
wire n_462;
wire n_1150;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_1165;
wire n_1185;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_816;
wire n_697;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_1058;
wire n_1105;
wire n_1163;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_1000;
wire n_984;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_1038;
wire n_1157;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_1186;
wire n_657;
wire n_764;
wire n_1156;
wire n_1206;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_947;
wire n_559;
wire n_425;
wire n_1050;

INVx1_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_22),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_133),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_84),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_63),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_136),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_0),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_178),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_2),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_122),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_179),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_167),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_94),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_87),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_98),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_45),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_62),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_139),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_89),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_142),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_72),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_53),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_6),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_112),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_32),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_143),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_144),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_59),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_91),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_82),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_83),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_150),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_38),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_113),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_102),
.Y(n_237)
);

INVxp67_ASAP7_75t_SL g238 ( 
.A(n_3),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_64),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_43),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_101),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_110),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_79),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_103),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_151),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_88),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_57),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_0),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_153),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_195),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_95),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_118),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_129),
.Y(n_255)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_119),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_2),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_48),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_125),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_92),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_196),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_24),
.Y(n_263)
);

INVxp33_ASAP7_75t_SL g264 ( 
.A(n_169),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_26),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_127),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_31),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_97),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_130),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_106),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_123),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_145),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_177),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_41),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_183),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_99),
.Y(n_276)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_131),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_3),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_68),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_21),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_51),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_176),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_21),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_65),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_135),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_172),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_73),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_50),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_171),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_13),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_141),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_137),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_148),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_19),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_56),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_78),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_198),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_116),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_149),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_185),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_20),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_47),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_197),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_37),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_9),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_190),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_74),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_23),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_181),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_199),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_140),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_187),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_128),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_189),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_154),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_104),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_146),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_25),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_80),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_40),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_155),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_109),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_108),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_147),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_193),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_33),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_18),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_134),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_52),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_37),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_76),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_15),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_14),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_163),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_191),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_22),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_71),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_121),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_69),
.B(n_192),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_170),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_6),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_100),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_13),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_156),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_19),
.B(n_115),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_60),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_188),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_39),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_66),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_17),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_107),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_12),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_114),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_235),
.B(n_1),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_350),
.B(n_207),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_209),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_246),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_246),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_246),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_314),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_L g362 ( 
.A(n_314),
.B(n_42),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_334),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_209),
.Y(n_364)
);

BUFx8_ASAP7_75t_L g365 ( 
.A(n_345),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_330),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_202),
.B(n_1),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_304),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_234),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_202),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_234),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_234),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_314),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_330),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_314),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_223),
.Y(n_376)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_225),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_304),
.Y(n_378)
);

CKINVDCx8_ASAP7_75t_R g379 ( 
.A(n_211),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_314),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_345),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_258),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_267),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_278),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_314),
.Y(n_385)
);

AND2x2_ASAP7_75t_SL g386 ( 
.A(n_345),
.B(n_44),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_314),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_208),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_269),
.B(n_4),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_234),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_280),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_208),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_283),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_215),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_269),
.B(n_4),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_215),
.B(n_5),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_312),
.Y(n_397)
);

OA21x2_ASAP7_75t_L g398 ( 
.A1(n_226),
.A2(n_67),
.B(n_194),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_326),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_226),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_245),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_245),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_338),
.B(n_5),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_312),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_289),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_290),
.Y(n_406)
);

NOR2x1_ASAP7_75t_L g407 ( 
.A(n_294),
.B(n_46),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_338),
.B(n_326),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_301),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_312),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_305),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_312),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_308),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_332),
.B(n_7),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_332),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_210),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_289),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_327),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_291),
.B(n_7),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_291),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_210),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_225),
.B(n_318),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_336),
.B(n_8),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_343),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_225),
.B(n_8),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_217),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_352),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_296),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_296),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_217),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_318),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_303),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_201),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_303),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_318),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_204),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_220),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_250),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_205),
.Y(n_439)
);

AND2x2_ASAP7_75t_SL g440 ( 
.A(n_206),
.B(n_49),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_213),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_311),
.B(n_9),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_311),
.B(n_10),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_320),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_220),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_320),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_323),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_216),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_323),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_300),
.Y(n_450)
);

BUFx8_ASAP7_75t_L g451 ( 
.A(n_331),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_218),
.B(n_10),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_219),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_300),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_331),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_337),
.B(n_11),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_265),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g458 ( 
.A(n_221),
.B(n_81),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_337),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_333),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_346),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_346),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_222),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_347),
.B(n_11),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_224),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_367),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_431),
.B(n_435),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_357),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_381),
.B(n_347),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_377),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_381),
.B(n_227),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_386),
.A2(n_264),
.B1(n_263),
.B2(n_341),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_367),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_415),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_431),
.B(n_238),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_369),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_367),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_381),
.B(n_228),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_408),
.B(n_229),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_396),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_377),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_433),
.B(n_233),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_377),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_357),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_439),
.B(n_237),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_396),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_431),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_422),
.B(n_214),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_396),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_435),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_415),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_441),
.B(n_239),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_358),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_358),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_399),
.B(n_435),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_464),
.B(n_240),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_361),
.B(n_241),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_368),
.B(n_214),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_364),
.B(n_230),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_369),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_369),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_369),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_448),
.B(n_242),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_365),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_464),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_365),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_464),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_386),
.A2(n_264),
.B1(n_351),
.B2(n_349),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_378),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g510 ( 
.A1(n_440),
.A2(n_348),
.B1(n_342),
.B2(n_340),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_371),
.Y(n_511)
);

AO22x1_ASAP7_75t_L g512 ( 
.A1(n_365),
.A2(n_364),
.B1(n_425),
.B2(n_389),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_409),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_389),
.A2(n_440),
.B1(n_458),
.B2(n_356),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_359),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_359),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_453),
.B(n_243),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_438),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_443),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_458),
.B(n_230),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_363),
.B(n_244),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_463),
.B(n_247),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_409),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_429),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_429),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_371),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_465),
.B(n_248),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_355),
.B(n_249),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_436),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_451),
.B(n_232),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_398),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_451),
.B(n_252),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_457),
.B(n_232),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_451),
.B(n_376),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_382),
.B(n_254),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_460),
.B(n_379),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_417),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_398),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_446),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_383),
.B(n_257),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_356),
.A2(n_253),
.B1(n_293),
.B2(n_297),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_384),
.B(n_260),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_455),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_417),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_455),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_455),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_461),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_391),
.B(n_261),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_461),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_388),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_393),
.B(n_293),
.Y(n_551)
);

INVxp33_ASAP7_75t_SL g552 ( 
.A(n_388),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_461),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_406),
.B(n_262),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_394),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_394),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_400),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_411),
.B(n_268),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_413),
.B(n_270),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_395),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_400),
.Y(n_561)
);

AND2x2_ASAP7_75t_SL g562 ( 
.A(n_403),
.B(n_271),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_418),
.B(n_297),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_401),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_371),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_424),
.B(n_427),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_401),
.B(n_273),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_402),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_354),
.B(n_310),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_402),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_370),
.B(n_276),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_398),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_405),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_405),
.A2(n_444),
.B1(n_459),
.B2(n_428),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_428),
.B(n_282),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_392),
.B(n_310),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_432),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_432),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_444),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_366),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_447),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_447),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_414),
.B(n_284),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_417),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_449),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_392),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_423),
.A2(n_353),
.B1(n_344),
.B2(n_277),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_459),
.B(n_285),
.Y(n_589)
);

NOR2x1p5_ASAP7_75t_L g590 ( 
.A(n_416),
.B(n_203),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_360),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_366),
.Y(n_592)
);

OR2x6_ASAP7_75t_L g593 ( 
.A(n_419),
.B(n_339),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_417),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_442),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_360),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_416),
.B(n_286),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_373),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_373),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_375),
.B(n_287),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_375),
.B(n_288),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_407),
.B(n_295),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_380),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_380),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_371),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_385),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_513),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_560),
.B(n_421),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_496),
.A2(n_452),
.B1(n_456),
.B2(n_419),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_560),
.B(n_421),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_595),
.B(n_385),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_504),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_523),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_557),
.Y(n_614)
);

BUFx4f_ASAP7_75t_L g615 ( 
.A(n_536),
.Y(n_615)
);

NAND2x1p5_ASAP7_75t_L g616 ( 
.A(n_506),
.B(n_456),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_543),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_534),
.B(n_558),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_514),
.A2(n_430),
.B1(n_454),
.B2(n_450),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_534),
.B(n_212),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_543),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_545),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_558),
.B(n_387),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_483),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_557),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_496),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_545),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_497),
.B(n_231),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_547),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_474),
.Y(n_630)
);

OR2x6_ASAP7_75t_SL g631 ( 
.A(n_491),
.B(n_426),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_559),
.B(n_387),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_547),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_518),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_520),
.A2(n_454),
.B1(n_450),
.B2(n_445),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_559),
.B(n_255),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_518),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_529),
.B(n_251),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_551),
.B(n_266),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_496),
.A2(n_362),
.B1(n_462),
.B2(n_420),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_529),
.B(n_272),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_580),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_490),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_553),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_467),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_490),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_509),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_496),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_467),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_487),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_555),
.Y(n_651)
);

BUFx4f_ASAP7_75t_L g652 ( 
.A(n_528),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_524),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_497),
.B(n_274),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_521),
.B(n_256),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_563),
.B(n_259),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_SL g657 ( 
.A1(n_592),
.A2(n_374),
.B1(n_445),
.B2(n_437),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_521),
.B(n_328),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_509),
.B(n_426),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_525),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_594),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_550),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_512),
.B(n_430),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_533),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_532),
.B(n_279),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_520),
.A2(n_437),
.B1(n_362),
.B2(n_309),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_568),
.Y(n_667)
);

NAND2x1p5_ASAP7_75t_L g668 ( 
.A(n_530),
.B(n_298),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_468),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_484),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_495),
.B(n_299),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_552),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_570),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_479),
.B(n_302),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_479),
.B(n_306),
.Y(n_675)
);

NOR2x2_ASAP7_75t_L g676 ( 
.A(n_541),
.B(n_374),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_515),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_579),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_602),
.B(n_307),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_602),
.B(n_317),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_472),
.A2(n_325),
.B1(n_329),
.B2(n_324),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_556),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_516),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_532),
.B(n_281),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_566),
.B(n_319),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_493),
.Y(n_686)
);

OR2x6_ASAP7_75t_L g687 ( 
.A(n_541),
.B(n_321),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_475),
.B(n_322),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_494),
.Y(n_689)
);

AND3x2_ASAP7_75t_SL g690 ( 
.A(n_587),
.B(n_12),
.C(n_14),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_562),
.B(n_292),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_561),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_SL g693 ( 
.A(n_588),
.B(n_315),
.C(n_335),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_564),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_573),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_582),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_544),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_531),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_577),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_466),
.B(n_236),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_510),
.A2(n_462),
.B1(n_434),
.B2(n_420),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_473),
.B(n_275),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_585),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_575),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_477),
.B(n_316),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_578),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_594),
.Y(n_707)
);

INVx5_ASAP7_75t_L g708 ( 
.A(n_537),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_581),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_531),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_538),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_584),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_488),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_480),
.B(n_420),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_586),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_575),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_486),
.B(n_434),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_470),
.B(n_434),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_489),
.B(n_505),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_475),
.B(n_434),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_481),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_588),
.B(n_462),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_507),
.B(n_462),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_576),
.Y(n_724)
);

NOR3xp33_ASAP7_75t_L g725 ( 
.A(n_587),
.B(n_15),
.C(n_16),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_498),
.B(n_16),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_539),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_687),
.A2(n_508),
.B1(n_510),
.B2(n_528),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_611),
.B(n_508),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_637),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_634),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_611),
.B(n_618),
.Y(n_732)
);

O2A1O1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_618),
.A2(n_597),
.B(n_519),
.C(n_583),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_634),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_647),
.B(n_590),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_612),
.B(n_569),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_674),
.B(n_471),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_643),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_698),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_659),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_664),
.B(n_499),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_679),
.A2(n_680),
.B(n_675),
.C(n_674),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_698),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_687),
.A2(n_722),
.B1(n_679),
.B2(n_680),
.Y(n_744)
);

INVx8_ASAP7_75t_L g745 ( 
.A(n_663),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_687),
.A2(n_589),
.B1(n_540),
.B2(n_542),
.Y(n_746)
);

OR2x6_ASAP7_75t_L g747 ( 
.A(n_663),
.B(n_626),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_671),
.A2(n_593),
.B1(n_548),
.B2(n_471),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_675),
.B(n_478),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_626),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_719),
.A2(n_538),
.B(n_572),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_719),
.B(n_478),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_671),
.A2(n_593),
.B1(n_589),
.B2(n_572),
.Y(n_753)
);

BUFx2_ASAP7_75t_L g754 ( 
.A(n_652),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_698),
.A2(n_469),
.B(n_601),
.Y(n_755)
);

OAI21x1_ASAP7_75t_L g756 ( 
.A1(n_714),
.A2(n_723),
.B(n_717),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_710),
.A2(n_469),
.B(n_601),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_613),
.B(n_482),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_652),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_716),
.Y(n_760)
);

INVx4_ASAP7_75t_L g761 ( 
.A(n_648),
.Y(n_761)
);

BUFx8_ASAP7_75t_L g762 ( 
.A(n_724),
.Y(n_762)
);

BUFx12f_ASAP7_75t_L g763 ( 
.A(n_642),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_716),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_672),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_692),
.B(n_482),
.Y(n_766)
);

INVx8_ASAP7_75t_L g767 ( 
.A(n_663),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_630),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_662),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_645),
.Y(n_770)
);

INVx4_ASAP7_75t_L g771 ( 
.A(n_648),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_608),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_610),
.B(n_535),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_694),
.B(n_485),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_666),
.B(n_701),
.C(n_725),
.Y(n_775)
);

INVx5_ASAP7_75t_L g776 ( 
.A(n_648),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_649),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_624),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_631),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_651),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_713),
.B(n_554),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_643),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_646),
.Y(n_783)
);

AOI222xp33_ASAP7_75t_L g784 ( 
.A1(n_657),
.A2(n_554),
.B1(n_503),
.B2(n_517),
.C1(n_522),
.C2(n_527),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_710),
.A2(n_600),
.B(n_596),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_646),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_682),
.Y(n_787)
);

INVx5_ASAP7_75t_L g788 ( 
.A(n_711),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_714),
.A2(n_723),
.B(n_717),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_708),
.Y(n_790)
);

BUFx12f_ASAP7_75t_L g791 ( 
.A(n_628),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_695),
.B(n_485),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_699),
.A2(n_600),
.B(n_571),
.C(n_517),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_623),
.A2(n_632),
.B(n_700),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_623),
.Y(n_795)
);

A2O1A1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_706),
.A2(n_522),
.B(n_492),
.C(n_503),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_607),
.Y(n_797)
);

AO21x2_ASAP7_75t_L g798 ( 
.A1(n_685),
.A2(n_567),
.B(n_527),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_685),
.A2(n_574),
.B1(n_567),
.B2(n_546),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_726),
.B(n_593),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_619),
.A2(n_549),
.B(n_604),
.C(n_603),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_708),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_708),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_715),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_SL g805 ( 
.A(n_615),
.B(n_598),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_619),
.A2(n_606),
.B(n_574),
.C(n_591),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_632),
.A2(n_599),
.B(n_537),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_708),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_628),
.B(n_17),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_709),
.A2(n_537),
.B(n_390),
.C(n_372),
.Y(n_810)
);

AND2x2_ASAP7_75t_SL g811 ( 
.A(n_615),
.B(n_18),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_656),
.A2(n_537),
.B1(n_390),
.B2(n_372),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_655),
.B(n_20),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_667),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_661),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_700),
.A2(n_605),
.B(n_565),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_704),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_653),
.Y(n_818)
);

BUFx12f_ASAP7_75t_L g819 ( 
.A(n_655),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_SL g820 ( 
.A(n_704),
.B(n_650),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_660),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_721),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_635),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_677),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_702),
.A2(n_605),
.B(n_565),
.Y(n_825)
);

AOI21xp33_ASAP7_75t_L g826 ( 
.A1(n_640),
.A2(n_372),
.B(n_390),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_688),
.B(n_23),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_688),
.A2(n_372),
.B1(n_390),
.B2(n_397),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_658),
.B(n_681),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_661),
.Y(n_830)
);

CKINVDCx8_ASAP7_75t_R g831 ( 
.A(n_676),
.Y(n_831)
);

O2A1O1Ixp5_ASAP7_75t_L g832 ( 
.A1(n_665),
.A2(n_605),
.B(n_565),
.C(n_526),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_661),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_712),
.B(n_24),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_683),
.B(n_25),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_667),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_673),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_673),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_678),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_661),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_650),
.B(n_26),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_707),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_658),
.B(n_27),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_656),
.B(n_27),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_678),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_751),
.A2(n_693),
.B(n_636),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_731),
.Y(n_847)
);

AO31x2_ASAP7_75t_L g848 ( 
.A1(n_796),
.A2(n_718),
.A3(n_705),
.B(n_702),
.Y(n_848)
);

AOI211x1_ASAP7_75t_L g849 ( 
.A1(n_729),
.A2(n_636),
.B(n_720),
.C(n_691),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_728),
.A2(n_654),
.B1(n_705),
.B2(n_639),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_834),
.Y(n_851)
);

OA21x2_ASAP7_75t_L g852 ( 
.A1(n_816),
.A2(n_609),
.B(n_633),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_834),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_SL g854 ( 
.A1(n_831),
.A2(n_823),
.B1(n_811),
.B2(n_731),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_732),
.B(n_616),
.Y(n_855)
);

AO21x2_ASAP7_75t_L g856 ( 
.A1(n_825),
.A2(n_622),
.B(n_617),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_734),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_742),
.A2(n_684),
.B(n_620),
.Y(n_858)
);

NAND2x1p5_ASAP7_75t_L g859 ( 
.A(n_783),
.B(n_614),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_835),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_732),
.A2(n_749),
.B1(n_737),
.B2(n_752),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_835),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_818),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_773),
.B(n_616),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_740),
.A2(n_727),
.B1(n_629),
.B2(n_621),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_730),
.Y(n_866)
);

AOI21xp33_ASAP7_75t_L g867 ( 
.A1(n_775),
.A2(n_668),
.B(n_644),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_821),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_L g869 ( 
.A1(n_737),
.A2(n_668),
.B1(n_690),
.B2(n_627),
.Y(n_869)
);

AO31x2_ASAP7_75t_L g870 ( 
.A1(n_799),
.A2(n_696),
.A3(n_669),
.B(n_689),
.Y(n_870)
);

OAI21x1_ASAP7_75t_L g871 ( 
.A1(n_756),
.A2(n_789),
.B(n_832),
.Y(n_871)
);

OAI21x1_ASAP7_75t_L g872 ( 
.A1(n_785),
.A2(n_625),
.B(n_686),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_749),
.B(n_670),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_824),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_781),
.Y(n_875)
);

OA21x2_ASAP7_75t_L g876 ( 
.A1(n_810),
.A2(n_703),
.B(n_697),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_781),
.B(n_641),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_804),
.Y(n_878)
);

OAI21x1_ASAP7_75t_L g879 ( 
.A1(n_807),
.A2(n_638),
.B(n_126),
.Y(n_879)
);

AO21x2_ASAP7_75t_L g880 ( 
.A1(n_826),
.A2(n_397),
.B(n_404),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_794),
.A2(n_526),
.B(n_511),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_783),
.B(n_28),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_752),
.A2(n_397),
.B1(n_404),
.B2(n_410),
.Y(n_883)
);

OAI21x1_ASAP7_75t_L g884 ( 
.A1(n_755),
.A2(n_124),
.B(n_168),
.Y(n_884)
);

AOI221xp5_ASAP7_75t_L g885 ( 
.A1(n_733),
.A2(n_397),
.B1(n_404),
.B2(n_410),
.C(n_412),
.Y(n_885)
);

OAI21x1_ASAP7_75t_L g886 ( 
.A1(n_757),
.A2(n_120),
.B(n_165),
.Y(n_886)
);

OAI21x1_ASAP7_75t_L g887 ( 
.A1(n_739),
.A2(n_117),
.B(n_164),
.Y(n_887)
);

INVxp67_ASAP7_75t_SL g888 ( 
.A(n_827),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_729),
.A2(n_404),
.B1(n_410),
.B2(n_412),
.Y(n_889)
);

OAI21xp33_ASAP7_75t_SL g890 ( 
.A1(n_766),
.A2(n_28),
.B(n_29),
.Y(n_890)
);

AOI32xp33_ASAP7_75t_L g891 ( 
.A1(n_827),
.A2(n_809),
.A3(n_829),
.B1(n_813),
.B2(n_800),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_784),
.A2(n_410),
.B1(n_412),
.B2(n_502),
.Y(n_892)
);

OR2x6_ASAP7_75t_L g893 ( 
.A(n_745),
.B(n_29),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_770),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_762),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_750),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_806),
.A2(n_412),
.B(n_31),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_SL g898 ( 
.A1(n_745),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_743),
.A2(n_132),
.B(n_200),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_795),
.B(n_30),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_763),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_747),
.B(n_34),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_777),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_793),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_904)
);

OAI21x1_ASAP7_75t_SL g905 ( 
.A1(n_766),
.A2(n_35),
.B(n_36),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_744),
.A2(n_799),
.B(n_746),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_762),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_778),
.Y(n_908)
);

CKINVDCx16_ASAP7_75t_R g909 ( 
.A(n_779),
.Y(n_909)
);

AO21x1_ASAP7_75t_L g910 ( 
.A1(n_844),
.A2(n_54),
.B(n_55),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_844),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_760),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_SL g913 ( 
.A1(n_747),
.A2(n_750),
.B(n_809),
.Y(n_913)
);

NOR2x1_ASAP7_75t_SL g914 ( 
.A(n_747),
.B(n_776),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_SL g915 ( 
.A1(n_774),
.A2(n_58),
.B(n_61),
.C(n_70),
.Y(n_915)
);

CKINVDCx16_ASAP7_75t_R g916 ( 
.A(n_791),
.Y(n_916)
);

CKINVDCx6p67_ASAP7_75t_R g917 ( 
.A(n_822),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_798),
.B(n_75),
.Y(n_918)
);

AO21x2_ASAP7_75t_L g919 ( 
.A1(n_826),
.A2(n_526),
.B(n_511),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_843),
.Y(n_920)
);

OAI21x1_ASAP7_75t_SL g921 ( 
.A1(n_774),
.A2(n_77),
.B(n_85),
.Y(n_921)
);

OAI21x1_ASAP7_75t_L g922 ( 
.A1(n_812),
.A2(n_86),
.B(n_90),
.Y(n_922)
);

OA21x2_ASAP7_75t_L g923 ( 
.A1(n_775),
.A2(n_511),
.B(n_502),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_784),
.B(n_93),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_736),
.B(n_96),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_736),
.B(n_105),
.Y(n_926)
);

OA21x2_ASAP7_75t_L g927 ( 
.A1(n_744),
.A2(n_501),
.B(n_500),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_769),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_802),
.B(n_111),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_802),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_765),
.B(n_152),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_815),
.A2(n_157),
.B(n_159),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_815),
.A2(n_160),
.B(n_162),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_819),
.A2(n_772),
.B1(n_800),
.B2(n_735),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_792),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_788),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_792),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_758),
.A2(n_501),
.B1(n_500),
.B2(n_476),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_788),
.B(n_500),
.Y(n_939)
);

AO21x2_ASAP7_75t_L g940 ( 
.A1(n_746),
.A2(n_476),
.B(n_174),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_750),
.Y(n_941)
);

OAI21x1_ASAP7_75t_L g942 ( 
.A1(n_833),
.A2(n_840),
.B(n_782),
.Y(n_942)
);

BUFx10_ASAP7_75t_L g943 ( 
.A(n_841),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_768),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_758),
.Y(n_945)
);

AOI221xp5_ASAP7_75t_L g946 ( 
.A1(n_748),
.A2(n_476),
.B1(n_175),
.B2(n_184),
.C(n_186),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_SL g947 ( 
.A1(n_745),
.A2(n_166),
.B1(n_767),
.B2(n_841),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_767),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_767),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_764),
.Y(n_950)
);

INVxp67_ASAP7_75t_SL g951 ( 
.A(n_754),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_788),
.Y(n_952)
);

OA21x2_ASAP7_75t_L g953 ( 
.A1(n_753),
.A2(n_828),
.B(n_797),
.Y(n_953)
);

INVx6_ASAP7_75t_L g954 ( 
.A(n_776),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_790),
.Y(n_955)
);

OA21x2_ASAP7_75t_L g956 ( 
.A1(n_814),
.A2(n_836),
.B(n_837),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_790),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_842),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_738),
.A2(n_786),
.B(n_782),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_780),
.B(n_787),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_842),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_790),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_801),
.A2(n_798),
.B1(n_838),
.B2(n_845),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_759),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_741),
.A2(n_839),
.B(n_820),
.C(n_805),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_817),
.B(n_830),
.Y(n_966)
);

OA21x2_ASAP7_75t_L g967 ( 
.A1(n_820),
.A2(n_805),
.B(n_842),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_786),
.A2(n_803),
.B1(n_808),
.B2(n_761),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_803),
.A2(n_808),
.B(n_776),
.Y(n_969)
);

O2A1O1Ixp5_ASAP7_75t_L g970 ( 
.A1(n_761),
.A2(n_771),
.B(n_808),
.C(n_803),
.Y(n_970)
);

INVx4_ASAP7_75t_L g971 ( 
.A(n_771),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_874),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_935),
.B(n_937),
.Y(n_973)
);

AND2x6_ASAP7_75t_SL g974 ( 
.A(n_893),
.B(n_901),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_861),
.A2(n_924),
.B1(n_945),
.B2(n_854),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_854),
.B(n_888),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_895),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_SL g978 ( 
.A1(n_948),
.A2(n_949),
.B1(n_893),
.B2(n_947),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_857),
.B(n_861),
.Y(n_979)
);

INVx6_ASAP7_75t_L g980 ( 
.A(n_916),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_902),
.A2(n_906),
.B1(n_947),
.B2(n_869),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_917),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_902),
.A2(n_906),
.B1(n_860),
.B2(n_862),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_SL g984 ( 
.A1(n_893),
.A2(n_882),
.B1(n_857),
.B2(n_943),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_891),
.A2(n_873),
.B1(n_851),
.B2(n_853),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_863),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_868),
.Y(n_987)
);

AO21x2_ASAP7_75t_L g988 ( 
.A1(n_897),
.A2(n_918),
.B(n_889),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_928),
.Y(n_989)
);

AOI211xp5_ASAP7_75t_L g990 ( 
.A1(n_890),
.A2(n_904),
.B(n_882),
.C(n_847),
.Y(n_990)
);

AOI221xp5_ASAP7_75t_L g991 ( 
.A1(n_875),
.A2(n_920),
.B1(n_850),
.B2(n_903),
.C(n_894),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_873),
.Y(n_992)
);

OAI221xp5_ASAP7_75t_L g993 ( 
.A1(n_934),
.A2(n_892),
.B1(n_865),
.B2(n_846),
.C(n_877),
.Y(n_993)
);

OR2x6_ASAP7_75t_L g994 ( 
.A(n_913),
.B(n_907),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_900),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_900),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_847),
.Y(n_997)
);

OA21x2_ASAP7_75t_L g998 ( 
.A1(n_871),
.A2(n_897),
.B(n_918),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_864),
.A2(n_911),
.B1(n_944),
.B2(n_926),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_878),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_925),
.A2(n_926),
.B1(n_855),
.B2(n_846),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_912),
.Y(n_1002)
);

OAI221xp5_ASAP7_75t_L g1003 ( 
.A1(n_898),
.A2(n_858),
.B1(n_855),
.B2(n_885),
.C(n_964),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_950),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_SL g1005 ( 
.A1(n_943),
.A2(n_925),
.B1(n_905),
.B2(n_914),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_SL g1006 ( 
.A1(n_929),
.A2(n_951),
.B1(n_931),
.B2(n_909),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_881),
.A2(n_858),
.B(n_965),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_964),
.A2(n_866),
.B1(n_936),
.B2(n_960),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_898),
.A2(n_849),
.B1(n_885),
.B2(n_929),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_952),
.Y(n_1010)
);

AOI222xp33_ASAP7_75t_L g1011 ( 
.A1(n_960),
.A2(n_963),
.B1(n_966),
.B2(n_908),
.C1(n_946),
.C2(n_936),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_952),
.Y(n_1012)
);

AO21x2_ASAP7_75t_L g1013 ( 
.A1(n_880),
.A2(n_940),
.B(n_919),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_930),
.B(n_952),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_963),
.A2(n_946),
.B1(n_904),
.B2(n_938),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_956),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_955),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_956),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_SL g1019 ( 
.A(n_971),
.B(n_941),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_848),
.B(n_859),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_867),
.A2(n_953),
.B1(n_930),
.B2(n_971),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_859),
.B(n_954),
.Y(n_1022)
);

OR2x6_ASAP7_75t_L g1023 ( 
.A(n_954),
.B(n_969),
.Y(n_1023)
);

AOI221xp5_ASAP7_75t_L g1024 ( 
.A1(n_867),
.A2(n_883),
.B1(n_938),
.B2(n_921),
.C(n_915),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_953),
.A2(n_968),
.B1(n_957),
.B2(n_962),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_957),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_852),
.A2(n_856),
.B1(n_957),
.B2(n_962),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_848),
.B(n_870),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_852),
.A2(n_856),
.B1(n_962),
.B2(n_961),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_872),
.A2(n_919),
.B(n_923),
.Y(n_1030)
);

AO31x2_ASAP7_75t_L g1031 ( 
.A1(n_910),
.A2(n_883),
.A3(n_870),
.B(n_923),
.Y(n_1031)
);

OA21x2_ASAP7_75t_L g1032 ( 
.A1(n_922),
.A2(n_899),
.B(n_887),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_958),
.A2(n_940),
.B1(n_959),
.B2(n_876),
.Y(n_1033)
);

AOI221xp5_ASAP7_75t_L g1034 ( 
.A1(n_970),
.A2(n_939),
.B1(n_848),
.B2(n_896),
.C(n_941),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_967),
.A2(n_941),
.B1(n_896),
.B2(n_927),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_870),
.B(n_942),
.Y(n_1036)
);

NOR2xp67_ASAP7_75t_L g1037 ( 
.A(n_970),
.B(n_879),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_884),
.A2(n_886),
.B1(n_932),
.B2(n_933),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_935),
.B(n_937),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_874),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_935),
.B(n_937),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_924),
.A2(n_634),
.B1(n_854),
.B2(n_861),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_924),
.A2(n_634),
.B1(n_854),
.B2(n_861),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_935),
.B(n_634),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_857),
.Y(n_1045)
);

AOI221xp5_ASAP7_75t_L g1046 ( 
.A1(n_861),
.A2(n_733),
.B1(n_619),
.B2(n_773),
.C(n_772),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_861),
.A2(n_935),
.B(n_945),
.C(n_937),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_861),
.A2(n_881),
.B(n_732),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_874),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_874),
.Y(n_1050)
);

AOI221xp5_ASAP7_75t_L g1051 ( 
.A1(n_861),
.A2(n_733),
.B1(n_619),
.B2(n_773),
.C(n_772),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_861),
.A2(n_906),
.B1(n_947),
.B2(n_937),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_SL g1053 ( 
.A1(n_854),
.A2(n_811),
.B1(n_745),
.B2(n_767),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_952),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_924),
.A2(n_634),
.B1(n_854),
.B2(n_861),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_917),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_874),
.Y(n_1057)
);

AND2x2_ASAP7_75t_SL g1058 ( 
.A(n_902),
.B(n_811),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_874),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_935),
.B(n_634),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_935),
.B(n_937),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_861),
.A2(n_906),
.B1(n_947),
.B2(n_937),
.Y(n_1062)
);

NAND2x1p5_ASAP7_75t_SL g1063 ( 
.A(n_1036),
.B(n_1012),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_992),
.B(n_1047),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_977),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_973),
.B(n_1044),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1060),
.B(n_979),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1016),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_975),
.B(n_972),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1018),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_1023),
.B(n_1048),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1050),
.B(n_1057),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1020),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_L g1075 ( 
.A(n_1062),
.B(n_1052),
.C(n_990),
.Y(n_1075)
);

INVx5_ASAP7_75t_SL g1076 ( 
.A(n_1022),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_1023),
.B(n_1037),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_SL g1078 ( 
.A1(n_1052),
.A2(n_1062),
.B(n_985),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_986),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1059),
.B(n_1039),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_1045),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_1010),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_987),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_1010),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_995),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1041),
.B(n_1061),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_996),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_985),
.B(n_997),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1000),
.B(n_1004),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_1058),
.B(n_978),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1002),
.B(n_981),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1046),
.B(n_1051),
.Y(n_1092)
);

AND2x4_ASAP7_75t_SL g1093 ( 
.A(n_1022),
.B(n_1014),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_1042),
.B(n_1043),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_1034),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_1054),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_1055),
.B(n_983),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1001),
.B(n_999),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_991),
.B(n_990),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1028),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1014),
.B(n_1006),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1025),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1053),
.B(n_984),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_1022),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_1054),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_1017),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1011),
.B(n_1009),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_976),
.B(n_1008),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1086),
.B(n_993),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1100),
.Y(n_1110)
);

OAI33xp33_ASAP7_75t_L g1111 ( 
.A1(n_1081),
.A2(n_1009),
.A3(n_1015),
.B1(n_989),
.B2(n_1035),
.B3(n_974),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_1063),
.Y(n_1112)
);

INVxp67_ASAP7_75t_SL g1113 ( 
.A(n_1068),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1086),
.B(n_994),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_L g1115 ( 
.A(n_1075),
.B(n_1011),
.C(n_1007),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1066),
.B(n_994),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1067),
.B(n_1029),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1070),
.Y(n_1118)
);

OAI211xp5_ASAP7_75t_L g1119 ( 
.A1(n_1090),
.A2(n_1103),
.B(n_1078),
.C(n_1092),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1075),
.A2(n_1003),
.B1(n_1005),
.B2(n_1015),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_1066),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1100),
.Y(n_1122)
);

AOI221xp5_ASAP7_75t_L g1123 ( 
.A1(n_1078),
.A2(n_1021),
.B1(n_982),
.B2(n_1056),
.C(n_1027),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1098),
.A2(n_994),
.B1(n_980),
.B2(n_1024),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_1063),
.Y(n_1125)
);

NAND4xp25_ASAP7_75t_L g1126 ( 
.A(n_1103),
.B(n_1033),
.C(n_1038),
.D(n_1030),
.Y(n_1126)
);

OAI33xp33_ASAP7_75t_L g1127 ( 
.A1(n_1079),
.A2(n_980),
.A3(n_1031),
.B1(n_988),
.B2(n_1019),
.B3(n_998),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1080),
.B(n_1071),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1080),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1070),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1071),
.B(n_1026),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1077),
.B(n_1013),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1073),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1073),
.B(n_1019),
.Y(n_1134)
);

INVx5_ASAP7_75t_L g1135 ( 
.A(n_1084),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1089),
.B(n_988),
.Y(n_1136)
);

INVxp67_ASAP7_75t_SL g1137 ( 
.A(n_1074),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1106),
.B(n_1032),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1121),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_1129),
.B(n_1067),
.Y(n_1140)
);

INVxp67_ASAP7_75t_SL g1141 ( 
.A(n_1113),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1133),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1130),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_1135),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1130),
.Y(n_1145)
);

OA21x2_ASAP7_75t_SL g1146 ( 
.A1(n_1128),
.A2(n_1107),
.B(n_1099),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1110),
.B(n_1088),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1137),
.B(n_1077),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1110),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1122),
.Y(n_1150)
);

OR2x6_ASAP7_75t_L g1151 ( 
.A(n_1112),
.B(n_1088),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1119),
.B(n_1108),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1122),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1116),
.B(n_1069),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_1135),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1118),
.Y(n_1156)
);

OAI221xp5_ASAP7_75t_L g1157 ( 
.A1(n_1120),
.A2(n_1107),
.B1(n_1099),
.B2(n_1094),
.C(n_1097),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1154),
.B(n_1117),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1143),
.B(n_1117),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1142),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1156),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1139),
.B(n_1069),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1140),
.B(n_1109),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1147),
.B(n_1091),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1147),
.B(n_1118),
.Y(n_1165)
);

NAND2x1_ASAP7_75t_L g1166 ( 
.A(n_1144),
.B(n_1112),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1148),
.B(n_1114),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1149),
.B(n_1091),
.Y(n_1168)
);

NOR2x1_ASAP7_75t_L g1169 ( 
.A(n_1144),
.B(n_1125),
.Y(n_1169)
);

NOR2xp67_ASAP7_75t_L g1170 ( 
.A(n_1155),
.B(n_1135),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1141),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1159),
.B(n_1151),
.Y(n_1172)
);

AOI211xp5_ASAP7_75t_L g1173 ( 
.A1(n_1170),
.A2(n_1157),
.B(n_1152),
.C(n_1120),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1164),
.A2(n_1152),
.B1(n_1157),
.B2(n_1111),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1161),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_R g1176 ( 
.A(n_1171),
.B(n_1125),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1169),
.A2(n_1115),
.B(n_1124),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_SL g1178 ( 
.A1(n_1171),
.A2(n_1146),
.B1(n_1148),
.B2(n_1101),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1167),
.A2(n_1123),
.B(n_1115),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_1165),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1161),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1160),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1166),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1159),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_1180),
.Y(n_1185)
);

INVxp67_ASAP7_75t_L g1186 ( 
.A(n_1182),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1174),
.B(n_1158),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1184),
.B(n_1158),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1178),
.B(n_1163),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1175),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1179),
.B(n_1162),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1173),
.A2(n_1151),
.B1(n_1101),
.B2(n_1168),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1183),
.A2(n_1093),
.B(n_1138),
.C(n_1141),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1172),
.B(n_1095),
.Y(n_1194)
);

XNOR2xp5_ASAP7_75t_L g1195 ( 
.A(n_1172),
.B(n_1065),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1186),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1193),
.A2(n_1183),
.B(n_1177),
.Y(n_1197)
);

AOI221x1_ASAP7_75t_L g1198 ( 
.A1(n_1191),
.A2(n_1183),
.B1(n_1126),
.B2(n_1079),
.C(n_1083),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1192),
.A2(n_1183),
.B(n_1093),
.C(n_1108),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1188),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1187),
.A2(n_1094),
.B(n_1097),
.C(n_1098),
.Y(n_1201)
);

OAI32xp33_ASAP7_75t_L g1202 ( 
.A1(n_1189),
.A2(n_1176),
.A3(n_1181),
.B1(n_1175),
.B2(n_1134),
.Y(n_1202)
);

OAI211xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1197),
.A2(n_1194),
.B(n_1185),
.C(n_1190),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1196),
.Y(n_1204)
);

AOI22x1_ASAP7_75t_SL g1205 ( 
.A1(n_1200),
.A2(n_1195),
.B1(n_1083),
.B2(n_1126),
.Y(n_1205)
);

AOI221xp5_ASAP7_75t_L g1206 ( 
.A1(n_1201),
.A2(n_1176),
.B1(n_1181),
.B2(n_1127),
.C(n_1153),
.Y(n_1206)
);

AOI221xp5_ASAP7_75t_L g1207 ( 
.A1(n_1202),
.A2(n_1150),
.B1(n_1095),
.B2(n_1145),
.C(n_1085),
.Y(n_1207)
);

AOI31xp33_ASAP7_75t_L g1208 ( 
.A1(n_1199),
.A2(n_1104),
.A3(n_1087),
.B(n_1131),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1204),
.Y(n_1209)
);

AOI221x1_ASAP7_75t_SL g1210 ( 
.A1(n_1203),
.A2(n_1198),
.B1(n_1199),
.B2(n_1087),
.C(n_1072),
.Y(n_1210)
);

NOR3xp33_ASAP7_75t_L g1211 ( 
.A(n_1208),
.B(n_1207),
.C(n_1206),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1205),
.Y(n_1212)
);

NAND5xp2_ASAP7_75t_L g1213 ( 
.A(n_1212),
.B(n_1064),
.C(n_1136),
.D(n_1102),
.E(n_1076),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_L g1214 ( 
.A(n_1211),
.B(n_1082),
.C(n_1084),
.Y(n_1214)
);

OR4x2_ASAP7_75t_L g1215 ( 
.A(n_1210),
.B(n_1151),
.C(n_1076),
.D(n_1063),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1214),
.A2(n_1209),
.B1(n_1076),
.B2(n_1132),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1215),
.B(n_1132),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1213),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1216),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1219),
.A2(n_1218),
.B(n_1217),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1220),
.A2(n_1076),
.B1(n_1093),
.B2(n_1132),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1221),
.Y(n_1222)
);

AOI222xp33_ASAP7_75t_L g1223 ( 
.A1(n_1222),
.A2(n_1076),
.B1(n_1082),
.B2(n_1096),
.C1(n_1105),
.C2(n_1135),
.Y(n_1223)
);


endmodule