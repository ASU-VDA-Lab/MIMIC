module fake_netlist_5_2448_n_1619 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1619);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1619;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_150;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_149;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_148;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_68),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_39),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_56),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_100),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_106),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_37),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_0),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_129),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_61),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_1),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_24),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_62),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_87),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_85),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_41),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_102),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_51),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_64),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_5),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_50),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_135),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_94),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_3),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_121),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_76),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_65),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_46),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_40),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_98),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_113),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_37),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_7),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_84),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_48),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_58),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_116),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_57),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_24),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_67),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_13),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_32),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_80),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_66),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_29),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_25),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_7),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_47),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_3),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_93),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_39),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_144),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_19),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_140),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_111),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_134),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_51),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_52),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_40),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_147),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_11),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_36),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_1),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_146),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_25),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_14),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_11),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_59),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_55),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_96),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_63),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_88),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_33),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_27),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_101),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_91),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_23),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_128),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_43),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_130),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_44),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_53),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_79),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_127),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_74),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_6),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_28),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_124),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_33),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_38),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_50),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_114),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_32),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_4),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_136),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_42),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_28),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_115),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_23),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_2),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_104),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_0),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_72),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_19),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_45),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_90),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_89),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_125),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_18),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_36),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_42),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_4),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_17),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_31),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_49),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_60),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_141),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_30),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_10),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_14),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_41),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_16),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_131),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_35),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_95),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_132),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_21),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_35),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_9),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_38),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_49),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_82),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_12),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_92),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g297 ( 
.A(n_249),
.B(n_2),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_155),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_282),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_155),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

INVxp33_ASAP7_75t_SL g303 ( 
.A(n_228),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_148),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_243),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_284),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_159),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_243),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_230),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_153),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_159),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_154),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_170),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_170),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_180),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_177),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_156),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_237),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_177),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_178),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_178),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_192),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_192),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_160),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_165),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_149),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_230),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_191),
.B(n_5),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_230),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_193),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_250),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_161),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_166),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_193),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_195),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_167),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_195),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_174),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_203),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_168),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_203),
.B(n_6),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_207),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_207),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_229),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_171),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_229),
.B(n_8),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_235),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_247),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_287),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_235),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_191),
.B(n_8),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_173),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_236),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_236),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_179),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_181),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_152),
.B(n_9),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_252),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_215),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_252),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_247),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_182),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_253),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_253),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_183),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_255),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_190),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_255),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_311),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_311),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_313),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_313),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_313),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_304),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_314),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_315),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_232),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_319),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_331),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_306),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_335),
.Y(n_386)
);

NOR2xp67_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_150),
.Y(n_387)
);

XNOR2x2_ASAP7_75t_L g388 ( 
.A(n_329),
.B(n_225),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_353),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_315),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_352),
.Y(n_391)
);

CKINVDCx11_ASAP7_75t_R g392 ( 
.A(n_312),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_317),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_363),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_329),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_352),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_318),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_321),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_328),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_318),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_336),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_365),
.B(n_246),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_299),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_337),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_365),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_330),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_299),
.B(n_258),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_298),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_360),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_333),
.B(n_296),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_298),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_322),
.A2(n_151),
.B(n_150),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_300),
.B(n_247),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_340),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_312),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_301),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_323),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_301),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_344),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_305),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_349),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_356),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_359),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_332),
.B(n_197),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_366),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_300),
.B(n_262),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_305),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_355),
.B(n_198),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_307),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_324),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_324),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_369),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_307),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_300),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_371),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_325),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_302),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_342),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_303),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_325),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_395),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_438),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_375),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_414),
.B(n_157),
.Y(n_448)
);

INVx5_ASAP7_75t_L g449 ( 
.A(n_391),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_444),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_327),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_176),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_430),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_441),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_438),
.B(n_308),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_444),
.A2(n_361),
.B1(n_341),
.B2(n_334),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_430),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_320),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_391),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_391),
.Y(n_461)
);

CKINVDCx8_ASAP7_75t_R g462 ( 
.A(n_378),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_419),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_428),
.B(n_320),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_391),
.Y(n_465)
);

INVx5_ASAP7_75t_L g466 ( 
.A(n_391),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_432),
.B(n_297),
.C(n_334),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_391),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_432),
.B(n_205),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_373),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_384),
.A2(n_341),
.B1(n_345),
.B2(n_350),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_417),
.B(n_345),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_373),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_374),
.Y(n_474)
);

BUFx10_ASAP7_75t_L g475 ( 
.A(n_442),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_384),
.A2(n_350),
.B1(n_297),
.B2(n_256),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_411),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_385),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_382),
.B(n_308),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_374),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_397),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_417),
.B(n_151),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_384),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_382),
.B(n_338),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_375),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_381),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_152),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_411),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_443),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

AO22x2_ASAP7_75t_L g491 ( 
.A1(n_388),
.A2(n_256),
.B1(n_275),
.B2(n_277),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_405),
.B(n_338),
.Y(n_492)
);

OR2x6_ASAP7_75t_L g493 ( 
.A(n_385),
.B(n_362),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_381),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_390),
.A2(n_277),
.B1(n_275),
.B2(n_291),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_397),
.Y(n_496)
);

BUFx10_ASAP7_75t_L g497 ( 
.A(n_379),
.Y(n_497)
);

BUFx4f_ASAP7_75t_L g498 ( 
.A(n_413),
.Y(n_498)
);

OR2x6_ASAP7_75t_L g499 ( 
.A(n_439),
.B(n_362),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_390),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_416),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_405),
.B(n_326),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_439),
.B(n_326),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_397),
.B(n_211),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_410),
.B(n_339),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_402),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_413),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_402),
.B(n_213),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_400),
.B(n_265),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_402),
.B(n_216),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_402),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

INVx4_ASAP7_75t_SL g515 ( 
.A(n_409),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_401),
.B(n_265),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_409),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_393),
.A2(n_291),
.B1(n_283),
.B2(n_164),
.Y(n_518)
);

AND2x2_ASAP7_75t_SL g519 ( 
.A(n_429),
.B(n_158),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_409),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_439),
.B(n_339),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_376),
.B(n_158),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_409),
.Y(n_523)
);

INVxp33_ASAP7_75t_SL g524 ( 
.A(n_404),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_408),
.B(n_343),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_418),
.B(n_343),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_423),
.B(n_162),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_398),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_416),
.B(n_346),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_398),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_376),
.B(n_162),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_425),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_399),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_377),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_409),
.B(n_217),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_392),
.B(n_283),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_L g537 ( 
.A(n_409),
.B(n_164),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_403),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_403),
.Y(n_539)
);

AND3x1_ASAP7_75t_L g540 ( 
.A(n_388),
.B(n_372),
.C(n_347),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_377),
.B(n_221),
.Y(n_541)
);

NOR2x1p5_ASAP7_75t_L g542 ( 
.A(n_426),
.B(n_188),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_431),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_431),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_406),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_406),
.Y(n_546)
);

AND2x2_ASAP7_75t_SL g547 ( 
.A(n_421),
.B(n_169),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_380),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_421),
.B(n_226),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_383),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_434),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_427),
.B(n_169),
.Y(n_552)
);

OR2x6_ASAP7_75t_L g553 ( 
.A(n_434),
.B(n_172),
.Y(n_553)
);

AND2x6_ASAP7_75t_L g554 ( 
.A(n_435),
.B(n_172),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_387),
.Y(n_555)
);

INVx8_ASAP7_75t_L g556 ( 
.A(n_436),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_386),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_435),
.B(n_440),
.Y(n_558)
);

CKINVDCx14_ASAP7_75t_R g559 ( 
.A(n_407),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_389),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_431),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_440),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_396),
.B(n_175),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_431),
.Y(n_564)
);

BUFx10_ASAP7_75t_L g565 ( 
.A(n_396),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_431),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_433),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_433),
.B(n_387),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_433),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_433),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_396),
.B(n_175),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_433),
.Y(n_572)
);

AND2x2_ASAP7_75t_SL g573 ( 
.A(n_412),
.B(n_184),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_412),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_433),
.Y(n_575)
);

INVx4_ASAP7_75t_SL g576 ( 
.A(n_412),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_415),
.B(n_346),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_415),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_420),
.B(n_184),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_420),
.B(n_347),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_422),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_422),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_538),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_464),
.B(n_185),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_464),
.B(n_185),
.Y(n_585)
);

NOR3xp33_ASAP7_75t_L g586 ( 
.A(n_445),
.B(n_199),
.C(n_189),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_451),
.B(n_186),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_451),
.B(n_186),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_503),
.B(n_187),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_519),
.B(n_231),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_538),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_525),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_545),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_503),
.B(n_187),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_L g595 ( 
.A(n_487),
.B(n_234),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_452),
.B(n_194),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_519),
.B(n_240),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_484),
.B(n_194),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_547),
.B(n_242),
.Y(n_599)
);

AOI221xp5_ASAP7_75t_L g600 ( 
.A1(n_491),
.A2(n_163),
.B1(n_267),
.B2(n_293),
.C(n_227),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_492),
.B(n_196),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_453),
.B(n_202),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_502),
.B(n_529),
.Y(n_603)
);

O2A1O1Ixp5_ASAP7_75t_L g604 ( 
.A1(n_482),
.A2(n_200),
.B(n_201),
.C(n_204),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_547),
.B(n_244),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_545),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_447),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_492),
.B(n_200),
.Y(n_608)
);

BUFx12f_ASAP7_75t_L g609 ( 
.A(n_557),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_459),
.B(n_257),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_446),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_448),
.B(n_206),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_447),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_485),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_483),
.B(n_201),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_483),
.B(n_479),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_467),
.A2(n_457),
.B1(n_553),
.B2(n_488),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_479),
.B(n_204),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_450),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_487),
.B(n_263),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_504),
.B(n_529),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_553),
.A2(n_233),
.B1(n_238),
.B2(n_245),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_469),
.B(n_233),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_525),
.Y(n_624)
);

A2O1A1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_495),
.A2(n_476),
.B(n_518),
.C(n_521),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_567),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_458),
.Y(n_627)
);

NAND2x1p5_ASAP7_75t_L g628 ( 
.A(n_502),
.B(n_238),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_472),
.B(n_245),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_470),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_485),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_540),
.A2(n_394),
.B1(n_222),
.B2(n_219),
.Y(n_632)
);

INVx8_ASAP7_75t_L g633 ( 
.A(n_556),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_526),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_472),
.B(n_254),
.Y(n_635)
);

OAI22xp33_ASAP7_75t_L g636 ( 
.A1(n_553),
.A2(n_477),
.B1(n_499),
.B2(n_558),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_493),
.B(n_348),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_555),
.B(n_254),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_555),
.B(n_260),
.Y(n_639)
);

BUFx5_ASAP7_75t_L g640 ( 
.A(n_487),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_521),
.B(n_260),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_473),
.B(n_268),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_556),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_476),
.A2(n_471),
.B1(n_456),
.B2(n_563),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_474),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_480),
.B(n_268),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_486),
.Y(n_647)
);

NAND3xp33_ASAP7_75t_SL g648 ( 
.A(n_563),
.B(n_571),
.C(n_552),
.Y(n_648)
);

NOR3xp33_ASAP7_75t_L g649 ( 
.A(n_508),
.B(n_218),
.C(n_214),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_494),
.B(n_269),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_500),
.Y(n_651)
);

BUFx6f_ASAP7_75t_SL g652 ( 
.A(n_497),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_501),
.B(n_269),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_528),
.B(n_424),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_530),
.B(n_424),
.Y(n_655)
);

NOR2xp67_ASAP7_75t_L g656 ( 
.A(n_526),
.B(n_270),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_504),
.B(n_573),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_487),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_455),
.B(n_259),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_527),
.B(n_208),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_573),
.B(n_278),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_524),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_533),
.B(n_424),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_527),
.B(n_209),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_491),
.A2(n_259),
.B1(n_264),
.B2(n_370),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_471),
.B(n_279),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_552),
.B(n_210),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_493),
.B(n_348),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_539),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_546),
.B(n_437),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_534),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_551),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_498),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_L g674 ( 
.A(n_487),
.B(n_285),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_510),
.B(n_212),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_454),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_562),
.B(n_437),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_577),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_574),
.B(n_288),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_579),
.B(n_351),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_478),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_582),
.B(n_294),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_582),
.B(n_351),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_549),
.B(n_354),
.Y(n_684)
);

AND2x2_ASAP7_75t_SL g685 ( 
.A(n_518),
.B(n_354),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_493),
.B(n_478),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_456),
.A2(n_280),
.B1(n_223),
.B2(n_224),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_541),
.B(n_357),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_506),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_578),
.B(n_498),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_506),
.B(n_259),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_463),
.B(n_281),
.C(n_239),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_499),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_499),
.A2(n_482),
.B1(n_579),
.B2(n_510),
.Y(n_694)
);

O2A1O1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_516),
.A2(n_372),
.B(n_370),
.C(n_368),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_578),
.B(n_505),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_489),
.B(n_259),
.Y(n_697)
);

OR2x6_ASAP7_75t_L g698 ( 
.A(n_556),
.B(n_358),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_578),
.B(n_358),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_578),
.B(n_364),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_509),
.B(n_364),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_516),
.B(n_220),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_542),
.Y(n_703)
);

A2O1A1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_495),
.A2(n_368),
.B(n_367),
.C(n_310),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_548),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_512),
.B(n_367),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_579),
.B(n_274),
.C(n_248),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_535),
.A2(n_276),
.B1(n_251),
.B2(n_295),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_462),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_567),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_465),
.B(n_286),
.Y(n_711)
);

NOR3xp33_ASAP7_75t_L g712 ( 
.A(n_559),
.B(n_273),
.C(n_266),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_581),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_490),
.B(n_496),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_507),
.A2(n_310),
.B(n_309),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_565),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_475),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_511),
.B(n_289),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_580),
.Y(n_719)
);

OR2x2_ASAP7_75t_SL g720 ( 
.A(n_491),
.B(n_264),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_554),
.B(n_290),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_554),
.B(n_272),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_513),
.B(n_271),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_554),
.B(n_292),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_566),
.B(n_241),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_576),
.B(n_569),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_576),
.B(n_264),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_554),
.B(n_309),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_567),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_576),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_592),
.B(n_550),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_624),
.B(n_497),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_696),
.A2(n_460),
.B(n_468),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_634),
.B(n_532),
.Y(n_734)
);

AOI21x1_ASAP7_75t_L g735 ( 
.A1(n_714),
.A2(n_568),
.B(n_570),
.Y(n_735)
);

O2A1O1Ixp5_ASAP7_75t_L g736 ( 
.A1(n_584),
.A2(n_514),
.B(n_517),
.C(n_575),
.Y(n_736)
);

CKINVDCx10_ASAP7_75t_R g737 ( 
.A(n_652),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_686),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_637),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_660),
.A2(n_537),
.B(n_517),
.C(n_514),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_656),
.B(n_532),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_644),
.A2(n_559),
.B1(n_536),
.B2(n_560),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_730),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_607),
.Y(n_744)
);

OA22x2_ASAP7_75t_L g745 ( 
.A1(n_689),
.A2(n_536),
.B1(n_475),
.B2(n_15),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_681),
.B(n_536),
.Y(n_746)
);

AOI21x1_ASAP7_75t_L g747 ( 
.A1(n_714),
.A2(n_515),
.B(n_520),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_630),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_612),
.B(n_460),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_657),
.A2(n_554),
.B1(n_537),
.B2(n_531),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_625),
.A2(n_481),
.B1(n_564),
.B2(n_449),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_645),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_633),
.Y(n_753)
);

NOR3xp33_ASAP7_75t_L g754 ( 
.A(n_660),
.B(n_564),
.C(n_522),
.Y(n_754)
);

NOR2x1_ASAP7_75t_L g755 ( 
.A(n_643),
.B(n_515),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_616),
.A2(n_523),
.B(n_461),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_647),
.Y(n_757)
);

O2A1O1Ixp5_ASAP7_75t_L g758 ( 
.A1(n_589),
.A2(n_522),
.B(n_531),
.C(n_515),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_657),
.A2(n_523),
.B(n_461),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_719),
.B(n_522),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_651),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_701),
.A2(n_706),
.B(n_626),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_626),
.A2(n_523),
.B(n_461),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_710),
.A2(n_523),
.B(n_461),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_611),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_625),
.A2(n_522),
.B(n_531),
.C(n_15),
.Y(n_766)
);

AO21x1_ASAP7_75t_L g767 ( 
.A1(n_628),
.A2(n_522),
.B(n_531),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_659),
.B(n_10),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_694),
.B(n_617),
.Y(n_769)
);

BUFx12f_ASAP7_75t_L g770 ( 
.A(n_609),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_617),
.B(n_572),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_668),
.B(n_13),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_587),
.B(n_531),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_729),
.A2(n_682),
.B(n_688),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_612),
.B(n_648),
.Y(n_775)
);

OAI321xp33_ASAP7_75t_L g776 ( 
.A1(n_664),
.A2(n_16),
.A3(n_17),
.B1(n_18),
.B2(n_20),
.C(n_21),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_588),
.B(n_466),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_730),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_676),
.B(n_22),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_603),
.B(n_466),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_669),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_L g782 ( 
.A(n_603),
.B(n_640),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_598),
.A2(n_572),
.B1(n_561),
.B2(n_544),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_611),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_664),
.B(n_22),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_684),
.A2(n_683),
.B(n_679),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_691),
.B(n_26),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_603),
.B(n_572),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_709),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_629),
.A2(n_561),
.B(n_544),
.Y(n_790)
);

AO21x1_ASAP7_75t_L g791 ( 
.A1(n_628),
.A2(n_34),
.B(n_43),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_693),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_599),
.A2(n_544),
.B1(n_543),
.B2(n_86),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_667),
.A2(n_544),
.B(n_543),
.C(n_47),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_635),
.A2(n_690),
.B(n_610),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_690),
.A2(n_543),
.B(n_81),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_603),
.B(n_543),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_603),
.B(n_78),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_672),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_619),
.Y(n_800)
);

NAND2x1_ASAP7_75t_L g801 ( 
.A(n_613),
.B(n_99),
.Y(n_801)
);

INVx8_ASAP7_75t_L g802 ( 
.A(n_633),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_601),
.B(n_103),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_608),
.B(n_75),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_673),
.B(n_107),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_667),
.A2(n_46),
.B(n_48),
.C(n_52),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_697),
.B(n_54),
.Y(n_807)
);

NOR2x1p5_ASAP7_75t_L g808 ( 
.A(n_643),
.B(n_69),
.Y(n_808)
);

OAI321xp33_ASAP7_75t_L g809 ( 
.A1(n_622),
.A2(n_70),
.A3(n_71),
.B1(n_108),
.B2(n_109),
.C(n_110),
.Y(n_809)
);

AOI21xp33_ASAP7_75t_L g810 ( 
.A1(n_618),
.A2(n_112),
.B(n_118),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_623),
.B(n_139),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_627),
.Y(n_812)
);

AO21x1_ASAP7_75t_L g813 ( 
.A1(n_594),
.A2(n_137),
.B(n_138),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_633),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_685),
.B(n_596),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_654),
.A2(n_655),
.B(n_677),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_666),
.A2(n_605),
.B(n_599),
.C(n_661),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_678),
.B(n_602),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_602),
.B(n_590),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_666),
.A2(n_661),
.B(n_631),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_590),
.B(n_597),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_663),
.A2(n_670),
.B(n_620),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_605),
.A2(n_597),
.B1(n_702),
.B2(n_675),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_675),
.A2(n_702),
.B1(n_636),
.B2(n_606),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_636),
.A2(n_583),
.B1(n_593),
.B2(n_591),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_685),
.B(n_680),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_725),
.A2(n_641),
.B(n_639),
.C(n_638),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_614),
.B(n_631),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_595),
.A2(n_674),
.B(n_715),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_720),
.B(n_687),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_709),
.Y(n_831)
);

O2A1O1Ixp5_ASAP7_75t_L g832 ( 
.A1(n_711),
.A2(n_723),
.B(n_718),
.C(n_722),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_658),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_699),
.A2(n_700),
.B(n_728),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_713),
.B(n_671),
.Y(n_835)
);

AO21x1_ASAP7_75t_L g836 ( 
.A1(n_622),
.A2(n_718),
.B(n_711),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_L g837 ( 
.A(n_600),
.B(n_665),
.C(n_586),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_725),
.B(n_646),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_723),
.A2(n_726),
.B(n_721),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_724),
.A2(n_705),
.B(n_642),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_703),
.A2(n_649),
.B1(n_692),
.B2(n_632),
.Y(n_841)
);

AO32x1_ASAP7_75t_L g842 ( 
.A1(n_708),
.A2(n_604),
.A3(n_716),
.B1(n_650),
.B2(n_653),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_727),
.B(n_704),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_658),
.A2(n_727),
.B(n_640),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_707),
.A2(n_695),
.B(n_704),
.C(n_658),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_658),
.A2(n_640),
.B(n_698),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_662),
.B(n_717),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_698),
.B(n_712),
.Y(n_848)
);

OR2x6_ASAP7_75t_L g849 ( 
.A(n_652),
.B(n_640),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_640),
.B(n_616),
.Y(n_850)
);

AOI21x1_ASAP7_75t_L g851 ( 
.A1(n_714),
.A2(n_726),
.B(n_615),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_696),
.A2(n_621),
.B(n_555),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_696),
.A2(n_621),
.B(n_555),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_592),
.B(n_457),
.Y(n_854)
);

AO21x1_ASAP7_75t_L g855 ( 
.A1(n_644),
.A2(n_585),
.B(n_584),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_660),
.A2(n_464),
.B(n_667),
.C(n_664),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_616),
.B(n_719),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_696),
.A2(n_621),
.B(n_555),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_660),
.A2(n_464),
.B(n_667),
.C(n_664),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_592),
.B(n_624),
.Y(n_860)
);

OA22x2_ASAP7_75t_L g861 ( 
.A1(n_644),
.A2(n_592),
.B1(n_634),
.B2(n_624),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_719),
.B(n_464),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_719),
.B(n_464),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_633),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_592),
.B(n_624),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_630),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_592),
.B(n_395),
.Y(n_867)
);

AOI21x1_ASAP7_75t_L g868 ( 
.A1(n_714),
.A2(n_726),
.B(n_615),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_697),
.Y(n_869)
);

INVx4_ASAP7_75t_L g870 ( 
.A(n_633),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_SL g871 ( 
.A1(n_720),
.A2(n_335),
.B1(n_353),
.B2(n_319),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_696),
.A2(n_621),
.B(n_555),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_607),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_696),
.A2(n_621),
.B(n_555),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_616),
.A2(n_621),
.B(n_657),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_696),
.A2(n_621),
.B(n_555),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_719),
.B(n_464),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_644),
.A2(n_621),
.B1(n_657),
.B2(n_464),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_696),
.A2(n_621),
.B(n_555),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_630),
.Y(n_880)
);

OAI21x1_ASAP7_75t_L g881 ( 
.A1(n_696),
.A2(n_714),
.B(n_730),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_719),
.B(n_464),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_616),
.A2(n_621),
.B(n_657),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_719),
.B(n_464),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_607),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_696),
.A2(n_621),
.B(n_555),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_696),
.A2(n_621),
.B(n_555),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_644),
.A2(n_464),
.B1(n_547),
.B2(n_519),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_681),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_856),
.A2(n_859),
.B(n_888),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_878),
.A2(n_815),
.B(n_861),
.Y(n_891)
);

AND2x6_ASAP7_75t_L g892 ( 
.A(n_833),
.B(n_823),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_862),
.B(n_863),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_829),
.A2(n_782),
.B(n_774),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_881),
.A2(n_747),
.B(n_735),
.Y(n_895)
);

AOI21x1_ASAP7_75t_L g896 ( 
.A1(n_850),
.A2(n_804),
.B(n_803),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_862),
.B(n_863),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_753),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_733),
.A2(n_868),
.B(n_851),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_835),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_877),
.B(n_882),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_819),
.B(n_775),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_884),
.B(n_857),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_789),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_835),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_786),
.A2(n_834),
.B(n_822),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_852),
.A2(n_858),
.B(n_853),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_748),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_840),
.A2(n_736),
.B(n_839),
.Y(n_909)
);

OA21x2_ASAP7_75t_L g910 ( 
.A1(n_820),
.A2(n_883),
.B(n_875),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_884),
.B(n_815),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_861),
.A2(n_817),
.B(n_769),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_753),
.Y(n_913)
);

OAI21x1_ASAP7_75t_L g914 ( 
.A1(n_872),
.A2(n_876),
.B(n_874),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_785),
.A2(n_758),
.B(n_843),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_753),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_821),
.B(n_838),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_818),
.B(n_860),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_879),
.A2(n_887),
.B(n_886),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_814),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_865),
.A2(n_806),
.B(n_869),
.C(n_830),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_867),
.B(n_749),
.Y(n_922)
);

AO31x2_ASAP7_75t_L g923 ( 
.A1(n_855),
.A2(n_836),
.A3(n_767),
.B(n_751),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_762),
.A2(n_816),
.B(n_795),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_833),
.Y(n_925)
);

OAI21x1_ASAP7_75t_L g926 ( 
.A1(n_844),
.A2(n_759),
.B(n_828),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_787),
.B(n_824),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_807),
.B(n_752),
.Y(n_928)
);

OAI21x1_ASAP7_75t_SL g929 ( 
.A1(n_846),
.A2(n_813),
.B(n_791),
.Y(n_929)
);

AND2x6_ASAP7_75t_L g930 ( 
.A(n_833),
.B(n_750),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_757),
.B(n_761),
.Y(n_931)
);

AOI221xp5_ASAP7_75t_L g932 ( 
.A1(n_837),
.A2(n_776),
.B1(n_871),
.B2(n_742),
.C(n_731),
.Y(n_932)
);

AOI21x1_ASAP7_75t_L g933 ( 
.A1(n_803),
.A2(n_804),
.B(n_751),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_870),
.B(n_814),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_781),
.B(n_799),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_827),
.B(n_826),
.Y(n_936)
);

AO31x2_ASAP7_75t_L g937 ( 
.A1(n_794),
.A2(n_740),
.A3(n_845),
.B(n_773),
.Y(n_937)
);

AOI21x1_ASAP7_75t_L g938 ( 
.A1(n_777),
.A2(n_773),
.B(n_756),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_784),
.B(n_814),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_854),
.B(n_889),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_738),
.Y(n_941)
);

OAI21x1_ASAP7_75t_L g942 ( 
.A1(n_780),
.A2(n_788),
.B(n_797),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_777),
.A2(n_780),
.B(n_788),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_797),
.A2(n_760),
.B(n_798),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_832),
.A2(n_825),
.B(n_766),
.C(n_768),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_831),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_798),
.A2(n_811),
.B(n_754),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_811),
.A2(n_793),
.B(n_885),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_792),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_734),
.B(n_739),
.Y(n_950)
);

NAND3xp33_ASAP7_75t_L g951 ( 
.A(n_841),
.B(n_880),
.C(n_866),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_771),
.A2(n_783),
.B(n_790),
.Y(n_952)
);

O2A1O1Ixp5_ASAP7_75t_L g953 ( 
.A1(n_805),
.A2(n_783),
.B(n_796),
.C(n_810),
.Y(n_953)
);

OAI21x1_ASAP7_75t_L g954 ( 
.A1(n_763),
.A2(n_764),
.B(n_873),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_800),
.B(n_812),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_SL g956 ( 
.A1(n_870),
.A2(n_849),
.B(n_864),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_743),
.A2(n_778),
.B(n_801),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_772),
.B(n_765),
.Y(n_958)
);

AO31x2_ASAP7_75t_L g959 ( 
.A1(n_842),
.A2(n_746),
.A3(n_809),
.B(n_810),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_778),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_849),
.A2(n_745),
.B1(n_808),
.B2(n_732),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_741),
.B(n_848),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_755),
.B(n_849),
.Y(n_963)
);

INVx5_ASAP7_75t_L g964 ( 
.A(n_864),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_779),
.A2(n_842),
.B(n_847),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_864),
.A2(n_802),
.B1(n_842),
.B2(n_770),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_802),
.B(n_737),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_856),
.A2(n_859),
.B(n_775),
.C(n_819),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_829),
.A2(n_782),
.B(n_696),
.Y(n_969)
);

NAND2x1_ASAP7_75t_L g970 ( 
.A(n_833),
.B(n_603),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_833),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_753),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_867),
.B(n_395),
.Y(n_973)
);

O2A1O1Ixp5_ASAP7_75t_L g974 ( 
.A1(n_856),
.A2(n_859),
.B(n_819),
.C(n_785),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_738),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_829),
.A2(n_782),
.B(n_696),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_835),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_881),
.A2(n_747),
.B(n_735),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_829),
.A2(n_782),
.B(n_696),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_881),
.A2(n_747),
.B(n_735),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_829),
.A2(n_782),
.B(n_696),
.Y(n_981)
);

AOI21xp33_ASAP7_75t_L g982 ( 
.A1(n_888),
.A2(n_859),
.B(n_856),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_770),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_738),
.Y(n_984)
);

AOI21x1_ASAP7_75t_L g985 ( 
.A1(n_850),
.A2(n_747),
.B(n_829),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_888),
.A2(n_859),
.B1(n_856),
.B2(n_644),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_856),
.A2(n_859),
.B(n_888),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_829),
.A2(n_782),
.B(n_696),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_856),
.A2(n_859),
.B(n_888),
.Y(n_989)
);

OAI22xp33_ASAP7_75t_L g990 ( 
.A1(n_823),
.A2(n_830),
.B1(n_624),
.B2(n_634),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_854),
.B(n_457),
.Y(n_991)
);

CKINVDCx16_ASAP7_75t_R g992 ( 
.A(n_770),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_784),
.B(n_753),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_829),
.A2(n_782),
.B(n_696),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_856),
.B(n_859),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_862),
.B(n_863),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_829),
.A2(n_782),
.B(n_696),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_835),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_867),
.B(n_395),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_856),
.A2(n_859),
.B(n_775),
.C(n_819),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_862),
.B(n_863),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_819),
.A2(n_775),
.B1(n_823),
.B2(n_856),
.Y(n_1002)
);

NOR2xp67_ASAP7_75t_SL g1003 ( 
.A(n_809),
.B(n_643),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_829),
.A2(n_782),
.B(n_696),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_744),
.Y(n_1005)
);

NAND2x1_ASAP7_75t_L g1006 ( 
.A(n_833),
.B(n_603),
.Y(n_1006)
);

AOI221xp5_ASAP7_75t_L g1007 ( 
.A1(n_837),
.A2(n_600),
.B1(n_540),
.B2(n_687),
.C(n_856),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_867),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_856),
.B(n_859),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_888),
.A2(n_859),
.B1(n_856),
.B2(n_644),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_862),
.B(n_863),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_829),
.A2(n_782),
.B(n_696),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_784),
.B(n_753),
.Y(n_1013)
);

OA21x2_ASAP7_75t_L g1014 ( 
.A1(n_820),
.A2(n_883),
.B(n_875),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_835),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_829),
.A2(n_782),
.B(n_696),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_SL g1017 ( 
.A1(n_767),
.A2(n_846),
.B(n_813),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_973),
.B(n_999),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_955),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_894),
.A2(n_906),
.B(n_924),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_970),
.Y(n_1021)
);

CKINVDCx16_ASAP7_75t_R g1022 ( 
.A(n_992),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_913),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_939),
.B(n_993),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_911),
.B(n_893),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_969),
.A2(n_979),
.B(n_976),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_983),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_904),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_1007),
.A2(n_1002),
.B1(n_932),
.B2(n_902),
.Y(n_1029)
);

AOI21xp33_ASAP7_75t_SL g1030 ( 
.A1(n_962),
.A2(n_991),
.B(n_961),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_931),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_922),
.B(n_918),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_941),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_964),
.B(n_1006),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_935),
.Y(n_1035)
);

OAI21xp33_ASAP7_75t_L g1036 ( 
.A1(n_940),
.A2(n_917),
.B(n_903),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_1008),
.B(n_917),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_974),
.A2(n_890),
.B(n_989),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_949),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_946),
.B(n_958),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_1005),
.Y(n_1041)
);

AND2x6_ASAP7_75t_L g1042 ( 
.A(n_936),
.B(n_900),
.Y(n_1042)
);

CKINVDCx8_ASAP7_75t_R g1043 ( 
.A(n_964),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_990),
.B(n_903),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_SL g1045 ( 
.A1(n_890),
.A2(n_987),
.B1(n_989),
.B2(n_1010),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_987),
.A2(n_986),
.B1(n_1010),
.B2(n_982),
.Y(n_1046)
);

NAND2x1p5_ASAP7_75t_L g1047 ( 
.A(n_964),
.B(n_898),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_981),
.A2(n_994),
.B(n_1016),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_911),
.B(n_893),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_975),
.B(n_928),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_905),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_913),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_897),
.B(n_901),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_939),
.B(n_993),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_925),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1001),
.B(n_1011),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_897),
.B(n_901),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_977),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_927),
.B(n_996),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_996),
.B(n_950),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_998),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_L g1062 ( 
.A(n_961),
.B(n_921),
.C(n_951),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_951),
.B(n_1015),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_960),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_967),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_968),
.B(n_1000),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_986),
.A2(n_982),
.B1(n_995),
.B2(n_1009),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1013),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_936),
.B(n_912),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_891),
.B(n_912),
.Y(n_1070)
);

AND2x6_ASAP7_75t_L g1071 ( 
.A(n_925),
.B(n_971),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_913),
.B(n_916),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_945),
.A2(n_891),
.B(n_915),
.C(n_953),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_971),
.Y(n_1074)
);

AO21x2_ASAP7_75t_L g1075 ( 
.A1(n_933),
.A2(n_947),
.B(n_929),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_988),
.A2(n_997),
.B(n_1004),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_916),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_965),
.B(n_963),
.Y(n_1078)
);

NAND2x1p5_ASAP7_75t_L g1079 ( 
.A(n_920),
.B(n_972),
.Y(n_1079)
);

AND2x6_ASAP7_75t_L g1080 ( 
.A(n_920),
.B(n_972),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_892),
.B(n_930),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_967),
.B(n_934),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_934),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_967),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_892),
.B(n_930),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_892),
.A2(n_1003),
.B1(n_930),
.B2(n_915),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_892),
.A2(n_930),
.B1(n_966),
.B2(n_1014),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_966),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_910),
.B(n_1014),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_910),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_937),
.B(n_923),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1012),
.A2(n_919),
.B(n_907),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_942),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_923),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_948),
.A2(n_914),
.B(n_944),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_948),
.A2(n_943),
.B(n_909),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_956),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_952),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_1017),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_926),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_957),
.A2(n_899),
.B(n_978),
.C(n_895),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_896),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_980),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_985),
.A2(n_938),
.B1(n_959),
.B2(n_954),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_959),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_959),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_984),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_908),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_973),
.B(n_999),
.Y(n_1109)
);

INVx1_ASAP7_75t_SL g1110 ( 
.A(n_946),
.Y(n_1110)
);

INVxp67_ASAP7_75t_L g1111 ( 
.A(n_940),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_939),
.B(n_993),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_908),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_968),
.A2(n_859),
.B(n_856),
.C(n_1000),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_913),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_973),
.B(n_999),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_939),
.B(n_993),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_939),
.B(n_993),
.Y(n_1118)
);

NOR2x1p5_ASAP7_75t_L g1119 ( 
.A(n_927),
.B(n_643),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_941),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_939),
.B(n_993),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_941),
.Y(n_1122)
);

INVxp67_ASAP7_75t_L g1123 ( 
.A(n_940),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_911),
.B(n_893),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_973),
.B(n_999),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_941),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_939),
.B(n_993),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_939),
.B(n_993),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1002),
.A2(n_888),
.B1(n_859),
.B2(n_856),
.Y(n_1129)
);

BUFx12f_ASAP7_75t_L g1130 ( 
.A(n_983),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_911),
.B(n_893),
.Y(n_1131)
);

NAND2x1p5_ASAP7_75t_L g1132 ( 
.A(n_964),
.B(n_970),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_911),
.B(n_893),
.Y(n_1133)
);

OA21x2_ASAP7_75t_L g1134 ( 
.A1(n_912),
.A2(n_909),
.B(n_890),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_904),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_908),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_908),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_973),
.B(n_999),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_968),
.A2(n_859),
.B(n_856),
.C(n_1000),
.Y(n_1139)
);

OAI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1029),
.A2(n_1129),
.B1(n_1059),
.B2(n_1057),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_1028),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_SL g1142 ( 
.A1(n_1081),
.A2(n_1085),
.B(n_1030),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1044),
.B(n_1138),
.Y(n_1143)
);

NAND3xp33_ASAP7_75t_L g1144 ( 
.A(n_1062),
.B(n_1129),
.C(n_1114),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1108),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_1135),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1066),
.A2(n_1139),
.B(n_1114),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_1080),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1043),
.Y(n_1149)
);

INVx6_ASAP7_75t_L g1150 ( 
.A(n_1083),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1113),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1137),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1051),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1071),
.Y(n_1154)
);

CKINVDCx6p67_ASAP7_75t_R g1155 ( 
.A(n_1130),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_1023),
.Y(n_1156)
);

AO21x1_ASAP7_75t_SL g1157 ( 
.A1(n_1086),
.A2(n_1087),
.B(n_1085),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1058),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1032),
.B(n_1056),
.Y(n_1159)
);

CKINVDCx6p67_ASAP7_75t_R g1160 ( 
.A(n_1022),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1061),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1096),
.A2(n_1095),
.B(n_1076),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1045),
.A2(n_1046),
.B1(n_1067),
.B2(n_1038),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1018),
.A2(n_1116),
.B1(n_1109),
.B2(n_1125),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1040),
.B(n_1050),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1036),
.B(n_1111),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1136),
.Y(n_1167)
);

NOR2x1_ASAP7_75t_L g1168 ( 
.A(n_1053),
.B(n_1057),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_1107),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1019),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1094),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_1033),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1097),
.B(n_1021),
.Y(n_1173)
);

BUFx4f_ASAP7_75t_SL g1174 ( 
.A(n_1084),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1090),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1025),
.B(n_1049),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_SL g1177 ( 
.A1(n_1067),
.A2(n_1038),
.B1(n_1081),
.B2(n_1102),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1039),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1045),
.A2(n_1063),
.B1(n_1069),
.B2(n_1070),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1023),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1070),
.A2(n_1035),
.B1(n_1031),
.B2(n_1060),
.Y(n_1181)
);

BUFx8_ASAP7_75t_L g1182 ( 
.A(n_1120),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_SL g1183 ( 
.A1(n_1042),
.A2(n_1088),
.B1(n_1065),
.B2(n_1099),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1111),
.B(n_1123),
.Y(n_1184)
);

BUFx2_ASAP7_75t_R g1185 ( 
.A(n_1027),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1064),
.Y(n_1186)
);

INVx4_ASAP7_75t_SL g1187 ( 
.A(n_1071),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1041),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1037),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1110),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_SL g1191 ( 
.A1(n_1042),
.A2(n_1088),
.B1(n_1124),
.B2(n_1131),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1134),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1098),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1134),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1123),
.B(n_1122),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1049),
.A2(n_1133),
.B1(n_1131),
.B2(n_1124),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1089),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_1126),
.Y(n_1198)
);

BUFx5_ASAP7_75t_L g1199 ( 
.A(n_1042),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_SL g1200 ( 
.A1(n_1042),
.A2(n_1133),
.B1(n_1105),
.B2(n_1097),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1074),
.Y(n_1201)
);

BUFx4f_ASAP7_75t_L g1202 ( 
.A(n_1080),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1068),
.Y(n_1203)
);

NAND2x1p5_ASAP7_75t_L g1204 ( 
.A(n_1082),
.B(n_1021),
.Y(n_1204)
);

AOI222xp33_ASAP7_75t_L g1205 ( 
.A1(n_1073),
.A2(n_1119),
.B1(n_1121),
.B2(n_1024),
.C1(n_1118),
.C2(n_1128),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1024),
.A2(n_1121),
.B1(n_1127),
.B2(n_1054),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_1054),
.Y(n_1207)
);

BUFx12f_ASAP7_75t_L g1208 ( 
.A(n_1112),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1042),
.A2(n_1078),
.B1(n_1098),
.B2(n_1075),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_SL g1210 ( 
.A1(n_1112),
.A2(n_1118),
.B1(n_1117),
.B2(n_1127),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1055),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1055),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1117),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1139),
.B(n_1128),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1091),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1106),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1072),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1075),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1079),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1023),
.B(n_1077),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_1052),
.Y(n_1221)
);

CKINVDCx11_ASAP7_75t_R g1222 ( 
.A(n_1052),
.Y(n_1222)
);

INVxp67_ASAP7_75t_SL g1223 ( 
.A(n_1020),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_1077),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1047),
.Y(n_1225)
);

BUFx8_ASAP7_75t_L g1226 ( 
.A(n_1080),
.Y(n_1226)
);

AO21x1_ASAP7_75t_L g1227 ( 
.A1(n_1104),
.A2(n_1095),
.B(n_1026),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_SL g1228 ( 
.A1(n_1047),
.A2(n_1132),
.B1(n_1034),
.B2(n_1115),
.Y(n_1228)
);

OAI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1115),
.A2(n_1132),
.B1(n_1034),
.B2(n_1103),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1100),
.B(n_1103),
.Y(n_1230)
);

AO21x2_ASAP7_75t_L g1231 ( 
.A1(n_1026),
.A2(n_1048),
.B(n_1076),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1048),
.A2(n_1101),
.B1(n_1092),
.B2(n_1093),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1092),
.A2(n_888),
.B1(n_859),
.B2(n_856),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1028),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1108),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1033),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1032),
.B(n_1056),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1108),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1028),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1022),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1192),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1143),
.B(n_1159),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1216),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1173),
.B(n_1197),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1196),
.B(n_1140),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1227),
.A2(n_1233),
.A3(n_1232),
.B(n_1194),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1143),
.B(n_1237),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1193),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1226),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1153),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1215),
.B(n_1147),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1226),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1190),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1196),
.B(n_1140),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1189),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1168),
.B(n_1176),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1230),
.B(n_1144),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1163),
.B(n_1175),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1163),
.B(n_1175),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1193),
.Y(n_1260)
);

INVxp67_ASAP7_75t_SL g1261 ( 
.A(n_1170),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1203),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1181),
.B(n_1179),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1171),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1171),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1170),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1179),
.B(n_1158),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1181),
.B(n_1218),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1177),
.A2(n_1166),
.B(n_1191),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1218),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1161),
.B(n_1157),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1166),
.A2(n_1214),
.B(n_1223),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1165),
.B(n_1214),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1200),
.B(n_1152),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1231),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1199),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1162),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1195),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1142),
.A2(n_1229),
.B(n_1186),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_1240),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1162),
.A2(n_1209),
.B(n_1154),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1162),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1183),
.B(n_1173),
.Y(n_1283)
);

AO21x2_ASAP7_75t_L g1284 ( 
.A1(n_1229),
.A2(n_1167),
.B(n_1201),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1199),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1169),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1199),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1209),
.B(n_1145),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1184),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1226),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1151),
.Y(n_1291)
);

AO21x1_ASAP7_75t_L g1292 ( 
.A1(n_1148),
.A2(n_1238),
.B(n_1235),
.Y(n_1292)
);

INVxp33_ASAP7_75t_L g1293 ( 
.A(n_1172),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1188),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1202),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1211),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1150),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1228),
.A2(n_1205),
.B(n_1204),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1204),
.B(n_1212),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1164),
.B(n_1213),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1187),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_SL g1302 ( 
.A1(n_1269),
.A2(n_1210),
.B(n_1206),
.Y(n_1302)
);

NAND2x1p5_ASAP7_75t_L g1303 ( 
.A(n_1276),
.B(n_1202),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1243),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1268),
.B(n_1236),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1241),
.B(n_1220),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1244),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1243),
.Y(n_1308)
);

OAI221xp5_ASAP7_75t_L g1309 ( 
.A1(n_1269),
.A2(n_1198),
.B1(n_1207),
.B2(n_1213),
.C(n_1178),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1244),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1244),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1251),
.B(n_1248),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1268),
.B(n_1246),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1251),
.B(n_1149),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1246),
.B(n_1160),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1246),
.B(n_1219),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1248),
.B(n_1260),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1246),
.B(n_1156),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1277),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1287),
.B(n_1225),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1260),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1282),
.A2(n_1221),
.B(n_1217),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1246),
.B(n_1180),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1284),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1244),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1270),
.B(n_1149),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1281),
.B(n_1156),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1270),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1242),
.B(n_1247),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1309),
.A2(n_1272),
.B1(n_1245),
.B2(n_1254),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1312),
.B(n_1272),
.Y(n_1331)
);

OAI21xp33_ASAP7_75t_L g1332 ( 
.A1(n_1329),
.A2(n_1263),
.B(n_1254),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1312),
.B(n_1278),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1324),
.A2(n_1275),
.B(n_1292),
.Y(n_1334)
);

AOI21xp33_ASAP7_75t_L g1335 ( 
.A1(n_1315),
.A2(n_1309),
.B(n_1329),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1319),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1305),
.B(n_1255),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1314),
.B(n_1298),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1304),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1302),
.A2(n_1298),
.B(n_1245),
.Y(n_1340)
);

NAND3xp33_ASAP7_75t_L g1341 ( 
.A(n_1315),
.B(n_1257),
.C(n_1263),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1305),
.B(n_1257),
.Y(n_1342)
);

NAND3xp33_ASAP7_75t_L g1343 ( 
.A(n_1315),
.B(n_1271),
.C(n_1256),
.Y(n_1343)
);

NOR3xp33_ASAP7_75t_SL g1344 ( 
.A(n_1302),
.B(n_1256),
.C(n_1299),
.Y(n_1344)
);

NAND2xp33_ASAP7_75t_R g1345 ( 
.A(n_1326),
.B(n_1273),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_SL g1346 ( 
.A1(n_1303),
.A2(n_1283),
.B(n_1271),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1307),
.B(n_1288),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1317),
.B(n_1273),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1303),
.A2(n_1283),
.B(n_1295),
.Y(n_1349)
);

OAI221xp5_ASAP7_75t_L g1350 ( 
.A1(n_1313),
.A2(n_1286),
.B1(n_1262),
.B2(n_1253),
.C(n_1141),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1303),
.B(n_1295),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1304),
.Y(n_1352)
);

NAND3xp33_ASAP7_75t_L g1353 ( 
.A(n_1324),
.B(n_1288),
.C(n_1274),
.Y(n_1353)
);

NAND3xp33_ASAP7_75t_L g1354 ( 
.A(n_1316),
.B(n_1274),
.C(n_1299),
.Y(n_1354)
);

OAI21xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1318),
.A2(n_1261),
.B(n_1250),
.Y(n_1355)
);

NAND3xp33_ASAP7_75t_L g1356 ( 
.A(n_1313),
.B(n_1316),
.C(n_1291),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1317),
.B(n_1289),
.Y(n_1357)
);

OAI221xp5_ASAP7_75t_L g1358 ( 
.A1(n_1313),
.A2(n_1300),
.B1(n_1293),
.B2(n_1234),
.C(n_1239),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1303),
.A2(n_1300),
.B1(n_1267),
.B2(n_1290),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1326),
.B(n_1280),
.Y(n_1360)
);

NAND3xp33_ASAP7_75t_L g1361 ( 
.A(n_1316),
.B(n_1291),
.C(n_1294),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1321),
.B(n_1267),
.Y(n_1362)
);

OAI221xp5_ASAP7_75t_L g1363 ( 
.A1(n_1326),
.A2(n_1146),
.B1(n_1239),
.B2(n_1234),
.C(n_1295),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1320),
.B(n_1249),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1310),
.B(n_1285),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1321),
.B(n_1258),
.Y(n_1366)
);

AOI221x1_ASAP7_75t_SL g1367 ( 
.A1(n_1308),
.A2(n_1265),
.B1(n_1264),
.B2(n_1294),
.C(n_1296),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1306),
.B(n_1258),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1311),
.B(n_1284),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1306),
.B(n_1259),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1311),
.A2(n_1259),
.B1(n_1174),
.B2(n_1208),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1306),
.B(n_1266),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_SL g1373 ( 
.A1(n_1318),
.A2(n_1149),
.B(n_1301),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1336),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1339),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1339),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1352),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1369),
.B(n_1318),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1342),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1369),
.B(n_1323),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1336),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1352),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1332),
.B(n_1340),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1347),
.B(n_1323),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1361),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1356),
.B(n_1322),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1347),
.B(n_1323),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1331),
.B(n_1328),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1361),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1365),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1356),
.B(n_1322),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1332),
.A2(n_1240),
.B1(n_1279),
.B2(n_1284),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1337),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1353),
.A2(n_1279),
.B1(n_1284),
.B2(n_1252),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1366),
.B(n_1322),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1362),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1372),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1334),
.B(n_1327),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1334),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1334),
.B(n_1327),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1333),
.B(n_1328),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1334),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1355),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1368),
.B(n_1327),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1370),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1377),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1377),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1377),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1378),
.B(n_1364),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1382),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1395),
.B(n_1354),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1403),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1383),
.B(n_1360),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1403),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1383),
.B(n_1394),
.C(n_1392),
.Y(n_1415)
);

NOR2x1p5_ASAP7_75t_L g1416 ( 
.A(n_1390),
.B(n_1155),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1382),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1395),
.B(n_1341),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1382),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1378),
.B(n_1373),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1375),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1378),
.B(n_1348),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1393),
.B(n_1335),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1401),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1375),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1374),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1376),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1392),
.A2(n_1338),
.B1(n_1344),
.B2(n_1330),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1374),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1380),
.B(n_1311),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1390),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1380),
.B(n_1325),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1395),
.B(n_1357),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1374),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1393),
.B(n_1367),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1379),
.B(n_1174),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1389),
.B(n_1343),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1379),
.B(n_1350),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1376),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1374),
.Y(n_1440)
);

NOR2x1_ASAP7_75t_SL g1441 ( 
.A(n_1386),
.B(n_1349),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1403),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1381),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1394),
.A2(n_1346),
.B1(n_1358),
.B2(n_1345),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1441),
.B(n_1420),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1421),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_1437),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1435),
.B(n_1404),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1441),
.B(n_1380),
.Y(n_1449)
);

NAND2x1_ASAP7_75t_L g1450 ( 
.A(n_1412),
.B(n_1390),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1438),
.B(n_1404),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1423),
.B(n_1404),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1421),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1412),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1426),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1425),
.Y(n_1456)
);

OR2x6_ASAP7_75t_L g1457 ( 
.A(n_1415),
.B(n_1249),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1420),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1413),
.B(n_1388),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1428),
.B(n_1388),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1409),
.B(n_1384),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1425),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1416),
.B(n_1389),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1409),
.B(n_1384),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1427),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1436),
.B(n_1396),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1424),
.B(n_1405),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1433),
.B(n_1405),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1427),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1444),
.A2(n_1386),
.B1(n_1391),
.B2(n_1385),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1439),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1437),
.B(n_1385),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1422),
.B(n_1405),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_1411),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1439),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1433),
.B(n_1405),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1411),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1418),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1422),
.B(n_1396),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1406),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1406),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1407),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1414),
.A2(n_1359),
.B1(n_1363),
.B2(n_1385),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1407),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1426),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1442),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_SL g1487 ( 
.A1(n_1418),
.A2(n_1371),
.B(n_1386),
.Y(n_1487)
);

OAI222xp33_ASAP7_75t_L g1488 ( 
.A1(n_1457),
.A2(n_1391),
.B1(n_1399),
.B2(n_1398),
.C1(n_1400),
.C2(n_1431),
.Y(n_1488)
);

CKINVDCx16_ASAP7_75t_R g1489 ( 
.A(n_1457),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1454),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1445),
.B(n_1430),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1486),
.B(n_1431),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1457),
.A2(n_1391),
.B1(n_1399),
.B2(n_1400),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1480),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1481),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1445),
.B(n_1430),
.Y(n_1496)
);

NOR2x1_ASAP7_75t_L g1497 ( 
.A(n_1450),
.B(n_1472),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1449),
.B(n_1432),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1449),
.B(n_1432),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1460),
.A2(n_1397),
.B1(n_1351),
.B2(n_1400),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1458),
.B(n_1384),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1447),
.B(n_1408),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1454),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1478),
.Y(n_1504)
);

AO22x1_ASAP7_75t_L g1505 ( 
.A1(n_1459),
.A2(n_1252),
.B1(n_1249),
.B2(n_1290),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_1486),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1448),
.B(n_1408),
.Y(n_1507)
);

NAND3xp33_ASAP7_75t_L g1508 ( 
.A(n_1472),
.B(n_1487),
.C(n_1459),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1474),
.B(n_1410),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1463),
.Y(n_1510)
);

CKINVDCx16_ASAP7_75t_R g1511 ( 
.A(n_1463),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1482),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1484),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1477),
.B(n_1410),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1446),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1461),
.B(n_1464),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1461),
.B(n_1387),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1452),
.B(n_1451),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1453),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1485),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1485),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1485),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1455),
.A2(n_1402),
.B(n_1440),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1504),
.B(n_1479),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_1504),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1518),
.B(n_1473),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1490),
.Y(n_1527)
);

AOI21xp33_ASAP7_75t_L g1528 ( 
.A1(n_1508),
.A2(n_1470),
.B(n_1466),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1490),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1508),
.B(n_1466),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1510),
.B(n_1463),
.Y(n_1531)
);

OAI32xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1488),
.A2(n_1483),
.A3(n_1467),
.B1(n_1462),
.B2(n_1465),
.Y(n_1532)
);

INVxp67_ASAP7_75t_L g1533 ( 
.A(n_1510),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1494),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1511),
.B(n_1464),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1494),
.Y(n_1536)
);

NOR3xp33_ASAP7_75t_L g1537 ( 
.A(n_1489),
.B(n_1469),
.C(n_1456),
.Y(n_1537)
);

AOI31xp33_ASAP7_75t_L g1538 ( 
.A1(n_1506),
.A2(n_1185),
.A3(n_1468),
.B(n_1476),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1518),
.B(n_1471),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1511),
.B(n_1506),
.Y(n_1540)
);

AOI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1488),
.A2(n_1475),
.B1(n_1398),
.B2(n_1402),
.C(n_1455),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1489),
.A2(n_1493),
.B1(n_1500),
.B2(n_1510),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1503),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_SL g1544 ( 
.A(n_1493),
.B(n_1402),
.C(n_1398),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1495),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1501),
.A2(n_1397),
.B1(n_1355),
.B2(n_1401),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1495),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1507),
.B(n_1146),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1525),
.B(n_1501),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1525),
.B(n_1503),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1530),
.B(n_1507),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1529),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1531),
.B(n_1491),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1543),
.B(n_1516),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1533),
.B(n_1516),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1524),
.B(n_1502),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1527),
.B(n_1491),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1540),
.B(n_1496),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1534),
.Y(n_1559)
);

AOI21xp33_ASAP7_75t_L g1560 ( 
.A1(n_1528),
.A2(n_1514),
.B(n_1497),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1536),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1531),
.B(n_1496),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1535),
.B(n_1514),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1539),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1545),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1526),
.B(n_1502),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1547),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1550),
.Y(n_1568)
);

NAND4xp25_ASAP7_75t_L g1569 ( 
.A(n_1551),
.B(n_1537),
.C(n_1542),
.D(n_1541),
.Y(n_1569)
);

AND2x2_ASAP7_75t_SL g1570 ( 
.A(n_1551),
.B(n_1548),
.Y(n_1570)
);

NOR2x1_ASAP7_75t_L g1571 ( 
.A(n_1552),
.B(n_1549),
.Y(n_1571)
);

AND4x1_ASAP7_75t_L g1572 ( 
.A(n_1563),
.B(n_1497),
.C(n_1532),
.D(n_1546),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_L g1573 ( 
.A1(n_1560),
.A2(n_1544),
.B1(n_1563),
.B2(n_1564),
.C(n_1554),
.Y(n_1573)
);

AOI21xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1556),
.A2(n_1538),
.B(n_1505),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1558),
.A2(n_1505),
.B(n_1509),
.Y(n_1575)
);

NAND3xp33_ASAP7_75t_SL g1576 ( 
.A(n_1555),
.B(n_1509),
.C(n_1515),
.Y(n_1576)
);

OAI211xp5_ASAP7_75t_SL g1577 ( 
.A1(n_1557),
.A2(n_1515),
.B(n_1519),
.C(n_1513),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1559),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1568),
.Y(n_1579)
);

AO22x1_ASAP7_75t_L g1580 ( 
.A1(n_1571),
.A2(n_1562),
.B1(n_1553),
.B2(n_1567),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1578),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1576),
.Y(n_1582)
);

AOI211xp5_ASAP7_75t_L g1583 ( 
.A1(n_1569),
.A2(n_1562),
.B(n_1566),
.C(n_1565),
.Y(n_1583)
);

NOR2x1_ASAP7_75t_L g1584 ( 
.A(n_1577),
.B(n_1561),
.Y(n_1584)
);

NOR2x1_ASAP7_75t_L g1585 ( 
.A(n_1575),
.B(n_1519),
.Y(n_1585)
);

NOR3x1_ASAP7_75t_L g1586 ( 
.A(n_1572),
.B(n_1513),
.C(n_1512),
.Y(n_1586)
);

OAI211xp5_ASAP7_75t_SL g1587 ( 
.A1(n_1573),
.A2(n_1512),
.B(n_1520),
.C(n_1521),
.Y(n_1587)
);

NOR2xp67_ASAP7_75t_L g1588 ( 
.A(n_1574),
.B(n_1522),
.Y(n_1588)
);

NAND4xp25_ASAP7_75t_L g1589 ( 
.A(n_1583),
.B(n_1570),
.C(n_1498),
.D(n_1499),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1580),
.B(n_1498),
.Y(n_1590)
);

AND3x1_ASAP7_75t_L g1591 ( 
.A(n_1582),
.B(n_1499),
.C(n_1520),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1588),
.Y(n_1592)
);

NOR3xp33_ASAP7_75t_SL g1593 ( 
.A(n_1587),
.B(n_1579),
.C(n_1581),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1592),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1591),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1590),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1593),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1589),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1589),
.A2(n_1584),
.B1(n_1585),
.B2(n_1492),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1599),
.B(n_1492),
.Y(n_1600)
);

NAND4xp25_ASAP7_75t_L g1601 ( 
.A(n_1598),
.B(n_1586),
.C(n_1521),
.D(n_1520),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1595),
.Y(n_1602)
);

AOI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1597),
.A2(n_1521),
.B1(n_1522),
.B2(n_1492),
.C(n_1517),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1594),
.B(n_1492),
.Y(n_1604)
);

AOI211x1_ASAP7_75t_L g1605 ( 
.A1(n_1600),
.A2(n_1601),
.B(n_1604),
.C(n_1596),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1602),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1603),
.B(n_1594),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1607),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1608),
.A2(n_1606),
.B1(n_1605),
.B2(n_1522),
.Y(n_1609)
);

OAI22x1_ASAP7_75t_L g1610 ( 
.A1(n_1609),
.A2(n_1522),
.B1(n_1182),
.B2(n_1517),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1609),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1610),
.A2(n_1523),
.B(n_1434),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1611),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1613),
.Y(n_1614)
);

OR3x1_ASAP7_75t_L g1615 ( 
.A(n_1612),
.B(n_1182),
.C(n_1222),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1614),
.B(n_1523),
.Y(n_1616)
);

AOI322xp5_ASAP7_75t_L g1617 ( 
.A1(n_1616),
.A2(n_1615),
.A3(n_1224),
.B1(n_1419),
.B2(n_1417),
.C1(n_1440),
.C2(n_1443),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1617),
.A2(n_1417),
.B1(n_1419),
.B2(n_1434),
.C(n_1429),
.Y(n_1618)
);

AOI211xp5_ASAP7_75t_L g1619 ( 
.A1(n_1618),
.A2(n_1290),
.B(n_1252),
.C(n_1297),
.Y(n_1619)
);


endmodule