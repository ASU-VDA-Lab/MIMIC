module fake_jpeg_13796_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_46),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_50),
.Y(n_100)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_6),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_49),
.B(n_54),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_15),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_6),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_78),
.Y(n_106)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_14),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_70),
.Y(n_113)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_14),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_43),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_76),
.Y(n_96)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_17),
.A2(n_5),
.B(n_7),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_80),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_82),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_28),
.B(n_5),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_90),
.Y(n_120)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_84),
.Y(n_124)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_86),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_87),
.B(n_89),
.Y(n_129)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_38),
.Y(n_137)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_28),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_36),
.B1(n_44),
.B2(n_41),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_92),
.A2(n_111),
.B1(n_115),
.B2(n_117),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_56),
.A2(n_44),
.B1(n_26),
.B2(n_34),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_97),
.A2(n_127),
.B1(n_91),
.B2(n_45),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_26),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_23),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_46),
.A2(n_55),
.B1(n_69),
.B2(n_86),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_58),
.A2(n_45),
.B1(n_44),
.B2(n_27),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_137),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_59),
.A2(n_87),
.B1(n_75),
.B2(n_68),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_49),
.B(n_22),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_134),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_54),
.B(n_34),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_28),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_61),
.Y(n_139)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_141),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_41),
.B(n_31),
.C(n_29),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_142),
.B(n_150),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_96),
.A2(n_62),
.B1(n_31),
.B2(n_29),
.Y(n_143)
);

OAI22x1_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_156),
.B1(n_163),
.B2(n_170),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_24),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_147),
.Y(n_183)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_107),
.A2(n_23),
.B(n_17),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_157),
.C(n_160),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_113),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_27),
.B1(n_24),
.B2(n_21),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_SL g184 ( 
.A1(n_153),
.A2(n_154),
.B(n_158),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_96),
.A2(n_61),
.B(n_21),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_121),
.A2(n_40),
.B1(n_45),
.B2(n_71),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_1),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_92),
.A2(n_76),
.B1(n_80),
.B2(n_40),
.Y(n_158)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_80),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_110),
.B1(n_133),
.B2(n_136),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_121),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_92),
.A2(n_1),
.B1(n_3),
.B2(n_7),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_110),
.B1(n_129),
.B2(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_1),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_166),
.C(n_168),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_7),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_12),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_105),
.A2(n_12),
.B1(n_14),
.B2(n_92),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_105),
.A2(n_12),
.B1(n_125),
.B2(n_128),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_171),
.A2(n_125),
.B1(n_126),
.B2(n_122),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_173),
.B1(n_160),
.B2(n_138),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_141),
.A2(n_132),
.B1(n_114),
.B2(n_120),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_150),
.B(n_130),
.CI(n_124),
.CON(n_177),
.SN(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_L g220 ( 
.A1(n_177),
.A2(n_174),
.B(n_175),
.C(n_180),
.D(n_172),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_192),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_155),
.B(n_151),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_148),
.B1(n_102),
.B2(n_159),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_165),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_SL g204 ( 
.A1(n_193),
.A2(n_160),
.B(n_169),
.C(n_167),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_128),
.B1(n_103),
.B2(n_95),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_197),
.B1(n_199),
.B2(n_126),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_95),
.B1(n_103),
.B2(n_99),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_162),
.A2(n_99),
.B1(n_102),
.B2(n_122),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_200),
.A2(n_221),
.B1(n_173),
.B2(n_184),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_186),
.A2(n_166),
.B1(n_147),
.B2(n_142),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_205),
.Y(n_233)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_220),
.B(n_176),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_194),
.A2(n_132),
.B1(n_149),
.B2(n_152),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_194),
.B(n_140),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_210),
.C(n_212),
.Y(n_226)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_152),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_191),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_183),
.B(n_140),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_179),
.B(n_152),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_168),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_213),
.B(n_215),
.Y(n_225)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_168),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_216),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_176),
.B(n_178),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_145),
.B1(n_146),
.B2(n_161),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

INVx6_ASAP7_75t_SL g223 ( 
.A(n_217),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_223),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_231),
.B(n_204),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_175),
.C(n_176),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_205),
.C(n_220),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_201),
.B1(n_221),
.B2(n_204),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_240),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_237),
.B(n_191),
.Y(n_245)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_245),
.C(n_256),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_242),
.A2(n_246),
.B1(n_251),
.B2(n_239),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_203),
.B1(n_214),
.B2(n_211),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_223),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_250),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_208),
.B1(n_204),
.B2(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_240),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_224),
.A2(n_221),
.B1(n_204),
.B2(n_207),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

AO22x1_ASAP7_75t_L g267 ( 
.A1(n_253),
.A2(n_237),
.B1(n_222),
.B2(n_233),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_188),
.B1(n_190),
.B2(n_187),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_236),
.B1(n_235),
.B2(n_229),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_178),
.C(n_187),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_253),
.A2(n_228),
.B(n_231),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_268),
.B1(n_243),
.B2(n_247),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_230),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_269),
.C(n_245),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_233),
.B(n_226),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_265),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_254),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_258),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_237),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_279),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_275),
.B1(n_278),
.B2(n_268),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_243),
.B1(n_254),
.B2(n_250),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_242),
.C(n_244),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_280),
.C(n_264),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_255),
.B1(n_252),
.B2(n_225),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_246),
.C(n_251),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_289),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_288),
.B1(n_238),
.B2(n_235),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_267),
.B(n_259),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_SL g291 ( 
.A1(n_285),
.A2(n_287),
.B(n_284),
.C(n_286),
.Y(n_291)
);

O2A1O1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_272),
.B(n_267),
.C(n_276),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_226),
.B1(n_266),
.B2(n_261),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_273),
.B(n_259),
.CI(n_225),
.CON(n_289),
.SN(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_284),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_292),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_291),
.A2(n_287),
.B(n_285),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_286),
.A2(n_271),
.B1(n_249),
.B2(n_229),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_293),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_283),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_295),
.B(n_283),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_296),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_289),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_291),
.A3(n_289),
.B1(n_238),
.B2(n_236),
.C1(n_190),
.C2(n_112),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_303),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_299),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_303),
.Y(n_306)
);

AOI321xp33_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_304),
.A3(n_236),
.B1(n_185),
.B2(n_181),
.C(n_182),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_307),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_185),
.B(n_189),
.C(n_112),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_189),
.Y(n_310)
);


endmodule