module fake_jpeg_4093_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_17),
.B(n_8),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.C(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_41),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_18),
.B(n_0),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_31),
.C(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_57),
.Y(n_81)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_37),
.Y(n_56)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_56),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_20),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_32),
.B1(n_16),
.B2(n_28),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_61),
.B1(n_16),
.B2(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_32),
.B1(n_16),
.B2(n_28),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_36),
.B(n_33),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_20),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_29),
.B(n_41),
.C(n_22),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_39),
.A2(n_32),
.B1(n_28),
.B2(n_31),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_68),
.B1(n_17),
.B2(n_22),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_32),
.B1(n_31),
.B2(n_20),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_29),
.Y(n_93)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_73),
.A2(n_62),
.B1(n_59),
.B2(n_16),
.Y(n_116)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_78),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_45),
.C(n_24),
.Y(n_114)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_89),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_60),
.B1(n_66),
.B2(n_64),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_66),
.B1(n_57),
.B2(n_55),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_53),
.B(n_47),
.Y(n_109)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_29),
.B(n_17),
.C(n_24),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_51),
.B(n_52),
.C(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_21),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_76),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_99),
.B(n_111),
.Y(n_137)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_106),
.Y(n_141)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_47),
.B1(n_66),
.B2(n_58),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_81),
.B1(n_75),
.B2(n_87),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_112),
.B(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_23),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_96),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_116),
.A2(n_120),
.B1(n_123),
.B2(n_61),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_59),
.B1(n_56),
.B2(n_62),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_89),
.B1(n_62),
.B2(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_45),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_72),
.Y(n_148)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_78),
.A2(n_59),
.B1(n_40),
.B2(n_69),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_136),
.Y(n_170)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_134),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_102),
.B1(n_105),
.B2(n_103),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_135),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_87),
.B1(n_67),
.B2(n_79),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_140),
.B1(n_144),
.B2(n_106),
.Y(n_169)
);

BUFx4f_ASAP7_75t_SL g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_97),
.A2(n_91),
.B1(n_79),
.B2(n_70),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

OA21x2_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_91),
.B(n_48),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_142),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_69),
.B1(n_78),
.B2(n_48),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_145),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_72),
.B1(n_77),
.B2(n_41),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_23),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_109),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_21),
.Y(n_174)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_152),
.B(n_154),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_150),
.B(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_155),
.B(n_156),
.Y(n_202)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_165),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_112),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_160),
.A2(n_161),
.B(n_166),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_147),
.A2(n_98),
.B(n_103),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_133),
.B1(n_139),
.B2(n_131),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_105),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_174),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_57),
.Y(n_166)
);

NOR2x1p5_ASAP7_75t_SL g167 ( 
.A(n_151),
.B(n_57),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_169),
.B1(n_129),
.B2(n_26),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_134),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_114),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_178),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_134),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_130),
.A2(n_104),
.B(n_119),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_167),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_190),
.Y(n_219)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_139),
.B1(n_128),
.B2(n_125),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_193),
.B1(n_195),
.B2(n_176),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_128),
.C(n_86),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_199),
.C(n_200),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_159),
.A2(n_77),
.B1(n_113),
.B2(n_125),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_159),
.A2(n_113),
.B1(n_122),
.B2(n_83),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_178),
.B(n_173),
.Y(n_218)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_165),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_126),
.B1(n_127),
.B2(n_86),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_198),
.A2(n_204),
.B1(n_206),
.B2(n_196),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_37),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_126),
.C(n_42),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_42),
.C(n_127),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_168),
.C(n_152),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_21),
.Y(n_203)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_162),
.B1(n_175),
.B2(n_164),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_21),
.Y(n_205)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_160),
.A2(n_49),
.B1(n_24),
.B2(n_22),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_153),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_226),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_171),
.Y(n_210)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_167),
.B(n_177),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_183),
.B(n_204),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_212),
.A2(n_194),
.B1(n_186),
.B2(n_203),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_216),
.B(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_224),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_231),
.B(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_223),
.C(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_172),
.C(n_171),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_181),
.B(n_157),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_166),
.B1(n_49),
.B2(n_26),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_225),
.A2(n_83),
.B1(n_27),
.B2(n_30),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_166),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_181),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_187),
.B(n_71),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_229),
.Y(n_239)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_42),
.C(n_71),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_49),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_42),
.C(n_71),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_193),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_235),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_201),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_206),
.B1(n_194),
.B2(n_188),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_236),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_214),
.C(n_223),
.Y(n_259)
);

XNOR2x1_ASAP7_75t_SL g240 ( 
.A(n_211),
.B(n_180),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_21),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_208),
.A2(n_222),
.B1(n_207),
.B2(n_215),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_243),
.B1(n_245),
.B2(n_253),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_207),
.A2(n_191),
.B1(n_197),
.B2(n_190),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_180),
.B1(n_195),
.B2(n_183),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_254),
.B1(n_234),
.B2(n_240),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_248),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_210),
.Y(n_257)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_218),
.B1(n_214),
.B2(n_212),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_225),
.A2(n_1),
.B(n_2),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_258),
.A2(n_260),
.B(n_2),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_264),
.C(n_18),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_232),
.B(n_226),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_83),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_27),
.B1(n_65),
.B2(n_21),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_27),
.C(n_21),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_1),
.Y(n_265)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_27),
.B1(n_30),
.B2(n_25),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_266),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_272),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_1),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_2),
.B(n_3),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_27),
.B1(n_30),
.B2(n_25),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_235),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_237),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_253),
.A2(n_30),
.B1(n_3),
.B2(n_4),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_268),
.A2(n_242),
.B1(n_238),
.B2(n_254),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_274),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_249),
.B(n_250),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_275),
.A2(n_276),
.B(n_283),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_260),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_237),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_280),
.A2(n_286),
.B(n_12),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_255),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_264),
.C(n_261),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_273),
.A2(n_3),
.B(n_4),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_3),
.B(n_5),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_265),
.B(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_259),
.C(n_255),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_295),
.C(n_296),
.Y(n_304)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_300),
.B(n_301),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_261),
.C(n_256),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_272),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_297),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_263),
.C(n_7),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_276),
.C(n_286),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_5),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_299),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_18),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_303),
.B1(n_285),
.B2(n_289),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_10),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_5),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_SL g307 ( 
.A(n_290),
.B(n_282),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_14),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_311),
.B(n_14),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_292),
.A2(n_291),
.B(n_303),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_288),
.B1(n_10),
.B2(n_11),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_321),
.C(n_306),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_316),
.A2(n_317),
.B(n_318),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g317 ( 
.A1(n_309),
.A2(n_11),
.B(n_13),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_13),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_319),
.B(n_320),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_13),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_326),
.B(n_15),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_304),
.C(n_312),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_323),
.A2(n_313),
.B(n_15),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_313),
.B(n_307),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_328),
.C(n_325),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_329),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_324),
.Y(n_331)
);


endmodule