module fake_netlist_5_1537_n_776 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_776);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_776;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_607;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_344;
wire n_287;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_289;
wire n_174;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_12),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_35),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_120),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_31),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_63),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_38),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_53),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_9),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_55),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_17),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_0),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_117),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_48),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_75),
.Y(n_173)
);

BUFx2_ASAP7_75t_SL g174 ( 
.A(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_50),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_81),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_143),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_124),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_78),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_17),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_60),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_77),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_86),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_93),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_72),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_90),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_24),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_83),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_98),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_4),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_13),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_36),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_26),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_144),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_4),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_67),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_68),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_12),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_22),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_97),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_201),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_0),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_165),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_156),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_201),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_159),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_157),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_1),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_166),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_171),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_172),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_179),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_159),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_180),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_173),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_182),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_173),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_1),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_160),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_181),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

NOR2xp67_ASAP7_75t_L g236 ( 
.A(n_170),
.B(n_2),
.Y(n_236)
);

BUFx2_ASAP7_75t_SL g237 ( 
.A(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_162),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_163),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_167),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_197),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_154),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_175),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_184),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_186),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_176),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

CKINVDCx8_ASAP7_75t_R g253 ( 
.A(n_210),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_208),
.A2(n_191),
.B1(n_204),
.B2(n_205),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_170),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_177),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_155),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_216),
.B(n_155),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_188),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_219),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_221),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_223),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_236),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_231),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_226),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_190),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_227),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_242),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_241),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_214),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_222),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_225),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_227),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_233),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_234),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_234),
.B(n_183),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_207),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_207),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_213),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_213),
.Y(n_293)
);

AOI22x1_ASAP7_75t_L g294 ( 
.A1(n_255),
.A2(n_203),
.B1(n_192),
.B2(n_200),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_247),
.B(n_196),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_250),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_251),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

AO21x2_ASAP7_75t_L g302 ( 
.A1(n_256),
.A2(n_198),
.B(n_195),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_264),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_258),
.B(n_195),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_258),
.B(n_158),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_265),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_268),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_265),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_266),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_266),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_278),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_263),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_158),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_266),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_247),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_247),
.B(n_187),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_261),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_266),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_249),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_247),
.B(n_189),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_247),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_249),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_272),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_270),
.B(n_199),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_269),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_267),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_260),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_267),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_276),
.B(n_199),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_289),
.Y(n_336)
);

OR2x6_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_174),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_260),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_255),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_273),
.B(n_193),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_257),
.B(n_202),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_277),
.Y(n_342)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_276),
.B(n_23),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_277),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_269),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_269),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_269),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_275),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_278),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_272),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_248),
.B(n_202),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_254),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_280),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_253),
.B(n_25),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_280),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_253),
.B(n_2),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_344),
.B(n_279),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_320),
.B(n_27),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_312),
.A2(n_282),
.B1(n_284),
.B2(n_293),
.Y(n_360)
);

OAI22xp33_ASAP7_75t_L g361 ( 
.A1(n_353),
.A2(n_279),
.B1(n_293),
.B2(n_281),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_311),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

NAND2xp33_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_279),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

AO22x2_ASAP7_75t_L g366 ( 
.A1(n_355),
.A2(n_285),
.B1(n_288),
.B2(n_292),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_312),
.B(n_327),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_303),
.Y(n_368)
);

BUFx8_ASAP7_75t_L g369 ( 
.A(n_316),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_297),
.Y(n_370)
);

AO22x2_ASAP7_75t_L g371 ( 
.A1(n_355),
.A2(n_285),
.B1(n_288),
.B2(n_292),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_304),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_318),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_R g374 ( 
.A(n_329),
.B(n_279),
.Y(n_374)
);

AO22x2_ASAP7_75t_L g375 ( 
.A1(n_354),
.A2(n_286),
.B1(n_291),
.B2(n_283),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_306),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_327),
.B(n_28),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_297),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_351),
.B(n_279),
.Y(n_379)
);

BUFx6f_ASAP7_75t_SL g380 ( 
.A(n_317),
.Y(n_380)
);

NAND2x1p5_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_298),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_342),
.A2(n_283),
.B1(n_287),
.B2(n_290),
.Y(n_382)
);

BUFx8_ASAP7_75t_L g383 ( 
.A(n_350),
.Y(n_383)
);

AO22x2_ASAP7_75t_L g384 ( 
.A1(n_356),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_309),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_299),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_351),
.Y(n_387)
);

AO22x2_ASAP7_75t_L g388 ( 
.A1(n_345),
.A2(n_342),
.B1(n_349),
.B2(n_339),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_328),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_300),
.Y(n_391)
);

NAND3xp33_ASAP7_75t_SL g392 ( 
.A(n_357),
.B(n_271),
.C(n_5),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_305),
.B(n_336),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_327),
.B(n_29),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_330),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_327),
.B(n_30),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_301),
.Y(n_397)
);

NOR4xp25_ASAP7_75t_SL g398 ( 
.A(n_347),
.B(n_271),
.C(n_6),
.D(n_7),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_337),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_305),
.B(n_3),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_338),
.B(n_32),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_338),
.B(n_330),
.Y(n_402)
);

AO22x2_ASAP7_75t_L g403 ( 
.A1(n_308),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_344),
.A2(n_85),
.B1(n_151),
.B2(n_149),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_344),
.B(n_8),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_299),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_307),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

AO22x2_ASAP7_75t_L g409 ( 
.A1(n_295),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_409)
);

OAI221xp5_ASAP7_75t_L g410 ( 
.A1(n_294),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.C(n_15),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_307),
.Y(n_411)
);

A2O1A1Ixp33_ASAP7_75t_L g412 ( 
.A1(n_310),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_336),
.B(n_16),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_335),
.Y(n_414)
);

AO22x2_ASAP7_75t_L g415 ( 
.A1(n_295),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_344),
.A2(n_89),
.B1(n_148),
.B2(n_145),
.Y(n_416)
);

NAND2xp33_ASAP7_75t_L g417 ( 
.A(n_348),
.B(n_33),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_322),
.B(n_34),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

AO22x2_ASAP7_75t_L g420 ( 
.A1(n_340),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_326),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_326),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_310),
.B(n_21),
.Y(n_423)
);

NAND2x1_ASAP7_75t_L g424 ( 
.A(n_298),
.B(n_37),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_363),
.B(n_348),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_373),
.B(n_331),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_395),
.B(n_335),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_414),
.B(n_387),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_393),
.B(n_331),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_379),
.B(n_346),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_379),
.B(n_346),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_374),
.B(n_341),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_400),
.B(n_352),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_337),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_423),
.B(n_321),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_367),
.B(n_402),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_413),
.B(n_325),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_397),
.B(n_340),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_SL g439 ( 
.A(n_380),
.B(n_302),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_361),
.B(n_357),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_360),
.B(n_302),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_SL g442 ( 
.A(n_398),
.B(n_333),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_401),
.B(n_333),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_401),
.B(n_332),
.Y(n_444)
);

NAND2xp33_ASAP7_75t_SL g445 ( 
.A(n_408),
.B(n_334),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_358),
.B(n_296),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_362),
.B(n_365),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_368),
.B(n_296),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_372),
.B(n_314),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_376),
.B(n_385),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_389),
.B(n_296),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_390),
.B(n_296),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_381),
.B(n_315),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_SL g454 ( 
.A(n_405),
.B(n_319),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_375),
.B(n_323),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_388),
.B(n_343),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_418),
.B(n_343),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_SL g458 ( 
.A(n_424),
.B(n_343),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_418),
.B(n_343),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_382),
.B(n_343),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_370),
.B(n_39),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_SL g462 ( 
.A(n_377),
.B(n_21),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_388),
.B(n_22),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_378),
.B(n_40),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_386),
.B(n_41),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_411),
.B(n_42),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_406),
.B(n_43),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_407),
.B(n_44),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_419),
.B(n_45),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_394),
.B(n_46),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_359),
.B(n_47),
.Y(n_471)
);

XNOR2x2_ASAP7_75t_L g472 ( 
.A(n_403),
.B(n_49),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_392),
.B(n_51),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_421),
.B(n_52),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_422),
.B(n_54),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_396),
.B(n_56),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_404),
.B(n_57),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_SL g478 ( 
.A(n_366),
.B(n_58),
.Y(n_478)
);

NAND2xp33_ASAP7_75t_SL g479 ( 
.A(n_366),
.B(n_371),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_416),
.B(n_59),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_364),
.B(n_61),
.Y(n_481)
);

AOI221x1_ASAP7_75t_L g482 ( 
.A1(n_479),
.A2(n_371),
.B1(n_415),
.B2(n_409),
.C(n_375),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_440),
.A2(n_433),
.B1(n_434),
.B2(n_438),
.Y(n_483)
);

AOI211x1_ASAP7_75t_L g484 ( 
.A1(n_463),
.A2(n_410),
.B(n_409),
.C(n_415),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_436),
.B(n_412),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_457),
.A2(n_417),
.B(n_399),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_459),
.A2(n_62),
.B(n_64),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_449),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_427),
.B(n_403),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_447),
.Y(n_490)
);

NAND3xp33_ASAP7_75t_SL g491 ( 
.A(n_473),
.B(n_420),
.C(n_369),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_455),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_450),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_435),
.B(n_420),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_437),
.B(n_384),
.Y(n_495)
);

AO21x2_ASAP7_75t_L g496 ( 
.A1(n_456),
.A2(n_384),
.B(n_66),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_430),
.A2(n_431),
.B(n_443),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_434),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_473),
.A2(n_369),
.B(n_383),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_475),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_444),
.A2(n_65),
.B(n_69),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_481),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_441),
.B(n_70),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_432),
.B(n_71),
.Y(n_505)
);

A2O1A1Ixp33_ASAP7_75t_L g506 ( 
.A1(n_442),
.A2(n_73),
.B(n_76),
.C(n_79),
.Y(n_506)
);

OAI22xp33_ASAP7_75t_L g507 ( 
.A1(n_428),
.A2(n_460),
.B1(n_472),
.B2(n_480),
.Y(n_507)
);

AO31x2_ASAP7_75t_L g508 ( 
.A1(n_478),
.A2(n_80),
.A3(n_82),
.B(n_84),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_425),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_426),
.B(n_87),
.Y(n_510)
);

OA21x2_ASAP7_75t_L g511 ( 
.A1(n_471),
.A2(n_88),
.B(n_91),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_429),
.B(n_92),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_448),
.Y(n_513)
);

OAI21x1_ASAP7_75t_SL g514 ( 
.A1(n_458),
.A2(n_94),
.B(n_95),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_451),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_452),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_477),
.B(n_96),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g518 ( 
.A(n_474),
.B(n_99),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_446),
.B(n_100),
.Y(n_519)
);

A2O1A1Ixp33_ASAP7_75t_L g520 ( 
.A1(n_439),
.A2(n_101),
.B(n_103),
.C(n_104),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_476),
.B(n_106),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_454),
.A2(n_108),
.B(n_109),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_453),
.B(n_110),
.Y(n_523)
);

O2A1O1Ixp33_ASAP7_75t_L g524 ( 
.A1(n_467),
.A2(n_111),
.B(n_112),
.C(n_113),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_R g525 ( 
.A(n_445),
.B(n_115),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_462),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_468),
.A2(n_116),
.B(n_118),
.Y(n_527)
);

NAND2x1p5_ASAP7_75t_L g528 ( 
.A(n_500),
.B(n_487),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_489),
.B(n_469),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_492),
.Y(n_530)
);

AOI221xp5_ASAP7_75t_L g531 ( 
.A1(n_507),
.A2(n_470),
.B1(n_466),
.B2(n_465),
.C(n_464),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_491),
.A2(n_461),
.B1(n_121),
.B2(n_122),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_488),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_485),
.Y(n_534)
);

NAND2x1p5_ASAP7_75t_L g535 ( 
.A(n_500),
.B(n_119),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_490),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_498),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_503),
.A2(n_123),
.B(n_125),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_511),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_502),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_485),
.A2(n_129),
.B(n_130),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_503),
.A2(n_131),
.B(n_133),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_526),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_489),
.B(n_134),
.Y(n_544)
);

OAI21x1_ASAP7_75t_SL g545 ( 
.A1(n_514),
.A2(n_136),
.B(n_137),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_483),
.B(n_140),
.Y(n_546)
);

AO21x2_ASAP7_75t_L g547 ( 
.A1(n_504),
.A2(n_141),
.B(n_142),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_527),
.A2(n_153),
.B(n_497),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_504),
.A2(n_517),
.B(n_505),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_494),
.A2(n_523),
.B1(n_493),
.B2(n_495),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_494),
.B(n_495),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_523),
.B(n_486),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_522),
.A2(n_505),
.B(n_512),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_522),
.A2(n_512),
.B(n_501),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_496),
.Y(n_555)
);

AOI21x1_ASAP7_75t_L g556 ( 
.A1(n_517),
.A2(n_513),
.B(n_516),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_509),
.A2(n_521),
.B1(n_510),
.B2(n_519),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_524),
.A2(n_511),
.B(n_515),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_509),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_509),
.B(n_518),
.Y(n_560)
);

BUFx2_ASAP7_75t_R g561 ( 
.A(n_496),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_484),
.B(n_482),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_520),
.B(n_506),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_508),
.Y(n_564)
);

OA21x2_ASAP7_75t_L g565 ( 
.A1(n_508),
.A2(n_499),
.B(n_525),
.Y(n_565)
);

OA21x2_ASAP7_75t_L g566 ( 
.A1(n_508),
.A2(n_485),
.B(n_482),
.Y(n_566)
);

NOR3xp33_ASAP7_75t_L g567 ( 
.A(n_491),
.B(n_281),
.C(n_290),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_492),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_534),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_566),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_551),
.B(n_534),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_566),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_566),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_549),
.A2(n_553),
.B(n_529),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_533),
.B(n_550),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_539),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_552),
.B(n_546),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_556),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_568),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_528),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_568),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_528),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_552),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_528),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_556),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_562),
.B(n_552),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_564),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_546),
.A2(n_563),
.B1(n_567),
.B2(n_544),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_536),
.Y(n_589)
);

BUFx4f_ASAP7_75t_SL g590 ( 
.A(n_543),
.Y(n_590)
);

INVxp67_ASAP7_75t_SL g591 ( 
.A(n_530),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_548),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_543),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_546),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_533),
.B(n_536),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_564),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_548),
.A2(n_554),
.B(n_553),
.Y(n_597)
);

HB1xp67_ASAP7_75t_SL g598 ( 
.A(n_537),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_560),
.B(n_563),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_554),
.A2(n_542),
.B(n_538),
.Y(n_601)
);

O2A1O1Ixp33_ASAP7_75t_L g602 ( 
.A1(n_563),
.A2(n_545),
.B(n_559),
.C(n_532),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_538),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_555),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_560),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_561),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_558),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_560),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_535),
.Y(n_609)
);

OAI21x1_ASAP7_75t_L g610 ( 
.A1(n_542),
.A2(n_558),
.B(n_545),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_557),
.B(n_565),
.Y(n_611)
);

AO21x1_ASAP7_75t_SL g612 ( 
.A1(n_565),
.A2(n_547),
.B(n_531),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_535),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_593),
.B(n_535),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_605),
.B(n_541),
.Y(n_615)
);

OR2x6_ASAP7_75t_L g616 ( 
.A(n_594),
.B(n_565),
.Y(n_616)
);

NAND2xp33_ASAP7_75t_R g617 ( 
.A(n_600),
.B(n_547),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_R g618 ( 
.A(n_600),
.B(n_547),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_608),
.B(n_540),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_569),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_590),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_569),
.Y(n_622)
);

INVx8_ASAP7_75t_L g623 ( 
.A(n_595),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_594),
.B(n_605),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_598),
.B(n_600),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_569),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_589),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_600),
.B(n_606),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_579),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_577),
.B(n_581),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_589),
.Y(n_631)
);

CKINVDCx14_ASAP7_75t_R g632 ( 
.A(n_581),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_577),
.B(n_594),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_586),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g635 ( 
.A(n_588),
.B(n_606),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_586),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_591),
.B(n_594),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_595),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_594),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_571),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_SL g641 ( 
.A(n_594),
.B(n_571),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_575),
.Y(n_642)
);

NAND2xp33_ASAP7_75t_R g643 ( 
.A(n_611),
.B(n_583),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_577),
.B(n_602),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_577),
.B(n_609),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_583),
.B(n_611),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_609),
.B(n_613),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_576),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_574),
.B(n_604),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_599),
.B(n_604),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_640),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_620),
.Y(n_652)
);

AND2x4_ASAP7_75t_SL g653 ( 
.A(n_625),
.B(n_599),
.Y(n_653)
);

INVxp67_ASAP7_75t_SL g654 ( 
.A(n_649),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_633),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_646),
.B(n_634),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_622),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_629),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_626),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_650),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_636),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_633),
.B(n_587),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_648),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_627),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_631),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_616),
.B(n_587),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_647),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_647),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_616),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_638),
.B(n_596),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_623),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_645),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_630),
.B(n_596),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_642),
.B(n_578),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_637),
.B(n_578),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_635),
.A2(n_613),
.B1(n_584),
.B2(n_580),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_645),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_656),
.B(n_630),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_676),
.B(n_644),
.C(n_628),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_656),
.B(n_570),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_666),
.B(n_570),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g682 ( 
.A(n_654),
.B(n_617),
.C(n_618),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_658),
.A2(n_632),
.B1(n_614),
.B2(n_653),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_651),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_661),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_671),
.Y(n_686)
);

NAND2x1p5_ASAP7_75t_L g687 ( 
.A(n_674),
.B(n_580),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_666),
.B(n_572),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_661),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_669),
.B(n_572),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_655),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_671),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_684),
.B(n_675),
.Y(n_693)
);

NOR2x1_ASAP7_75t_L g694 ( 
.A(n_682),
.B(n_674),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_685),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_691),
.B(n_669),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_678),
.B(n_681),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_686),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_689),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_690),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_679),
.B(n_667),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_680),
.B(n_688),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_690),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_678),
.B(n_688),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_701),
.B(n_681),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_SL g706 ( 
.A(n_693),
.B(n_686),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_701),
.A2(n_641),
.B1(n_683),
.B2(n_643),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_695),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_698),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_708),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_705),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_709),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_707),
.Y(n_713)
);

NOR2x1_ASAP7_75t_L g714 ( 
.A(n_706),
.B(n_694),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_705),
.B(n_702),
.Y(n_715)
);

OAI22xp33_ASAP7_75t_L g716 ( 
.A1(n_714),
.A2(n_692),
.B1(n_697),
.B2(n_704),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_712),
.B(n_702),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_713),
.A2(n_667),
.B(n_668),
.C(n_699),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_717),
.B(n_712),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_715),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_718),
.B(n_711),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_719),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_721),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_720),
.Y(n_724)
);

INVxp33_ASAP7_75t_SL g725 ( 
.A(n_719),
.Y(n_725)
);

NAND4xp25_ASAP7_75t_L g726 ( 
.A(n_724),
.B(n_672),
.C(n_677),
.D(n_668),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_725),
.B(n_621),
.Y(n_727)
);

NOR2x1_ASAP7_75t_L g728 ( 
.A(n_723),
.B(n_692),
.Y(n_728)
);

NAND5xp2_ASAP7_75t_L g729 ( 
.A(n_725),
.B(n_619),
.C(n_672),
.D(n_677),
.E(n_696),
.Y(n_729)
);

NOR2x1_ASAP7_75t_L g730 ( 
.A(n_722),
.B(n_692),
.Y(n_730)
);

NAND3xp33_ASAP7_75t_SL g731 ( 
.A(n_724),
.B(n_710),
.C(n_696),
.Y(n_731)
);

NAND4xp75_ASAP7_75t_L g732 ( 
.A(n_723),
.B(n_710),
.C(n_703),
.D(n_700),
.Y(n_732)
);

OAI221xp5_ASAP7_75t_SL g733 ( 
.A1(n_726),
.A2(n_624),
.B1(n_670),
.B2(n_655),
.C(n_660),
.Y(n_733)
);

NAND4xp25_ASAP7_75t_SL g734 ( 
.A(n_728),
.B(n_680),
.C(n_692),
.D(n_660),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_730),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_727),
.Y(n_736)
);

OAI221xp5_ASAP7_75t_L g737 ( 
.A1(n_731),
.A2(n_732),
.B1(n_729),
.B2(n_692),
.C(n_687),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_727),
.A2(n_653),
.B1(n_687),
.B2(n_655),
.Y(n_738)
);

AOI221xp5_ASAP7_75t_L g739 ( 
.A1(n_731),
.A2(n_664),
.B1(n_652),
.B2(n_657),
.C(n_659),
.Y(n_739)
);

AOI211xp5_ASAP7_75t_L g740 ( 
.A1(n_731),
.A2(n_615),
.B(n_639),
.C(n_664),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_735),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_736),
.B(n_673),
.Y(n_742)
);

NAND4xp75_ASAP7_75t_L g743 ( 
.A(n_739),
.B(n_662),
.C(n_652),
.D(n_657),
.Y(n_743)
);

XOR2xp5_ASAP7_75t_L g744 ( 
.A(n_738),
.B(n_639),
.Y(n_744)
);

XOR2x2_ASAP7_75t_L g745 ( 
.A(n_737),
.B(n_662),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_734),
.B(n_673),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_740),
.B(n_659),
.C(n_670),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_733),
.Y(n_748)
);

NOR2x1_ASAP7_75t_L g749 ( 
.A(n_735),
.B(n_624),
.Y(n_749)
);

NOR3xp33_ASAP7_75t_SL g750 ( 
.A(n_741),
.B(n_585),
.C(n_573),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_742),
.B(n_665),
.Y(n_751)
);

XNOR2x1_ASAP7_75t_L g752 ( 
.A(n_748),
.B(n_610),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_749),
.B(n_665),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_SL g754 ( 
.A(n_744),
.B(n_663),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_SL g755 ( 
.A(n_745),
.B(n_743),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_746),
.B(n_623),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_R g757 ( 
.A(n_747),
.B(n_603),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_L g758 ( 
.A(n_741),
.B(n_663),
.C(n_585),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_752),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_753),
.A2(n_603),
.B(n_580),
.C(n_582),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_751),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_756),
.A2(n_580),
.B1(n_582),
.B2(n_584),
.Y(n_762)
);

INVx5_ASAP7_75t_L g763 ( 
.A(n_755),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_763),
.Y(n_764)
);

OAI21x1_ASAP7_75t_L g765 ( 
.A1(n_759),
.A2(n_758),
.B(n_757),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_761),
.B(n_750),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_762),
.Y(n_767)
);

AOI21xp33_ASAP7_75t_L g768 ( 
.A1(n_764),
.A2(n_760),
.B(n_754),
.Y(n_768)
);

AO22x2_ASAP7_75t_L g769 ( 
.A1(n_767),
.A2(n_603),
.B1(n_582),
.B2(n_584),
.Y(n_769)
);

XNOR2xp5_ASAP7_75t_L g770 ( 
.A(n_765),
.B(n_610),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_768),
.A2(n_766),
.B1(n_612),
.B2(n_582),
.Y(n_771)
);

XOR2xp5_ASAP7_75t_L g772 ( 
.A(n_771),
.B(n_770),
.Y(n_772)
);

OA21x2_ASAP7_75t_L g773 ( 
.A1(n_772),
.A2(n_769),
.B(n_601),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_773),
.Y(n_774)
);

OAI221xp5_ASAP7_75t_L g775 ( 
.A1(n_774),
.A2(n_603),
.B1(n_592),
.B2(n_584),
.C(n_607),
.Y(n_775)
);

AOI211xp5_ASAP7_75t_L g776 ( 
.A1(n_775),
.A2(n_601),
.B(n_607),
.C(n_597),
.Y(n_776)
);


endmodule