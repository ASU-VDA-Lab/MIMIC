module fake_jpeg_32069_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx6_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_1),
.B(n_2),
.Y(n_11)
);

AOI21xp5_ASAP7_75t_L g12 ( 
.A1(n_0),
.A2(n_2),
.B(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_20),
.Y(n_25)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_23),
.Y(n_27)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_4),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_4),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_9),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_33),
.Y(n_45)
);

NOR2x1_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_23),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_17),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_16),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_22),
.B(n_19),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_19),
.C(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_40),
.B1(n_35),
.B2(n_38),
.Y(n_41)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_8),
.B1(n_10),
.B2(n_17),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_10),
.B(n_8),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_36),
.C(n_33),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_16),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

HAxp5_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_34),
.CON(n_51),
.SN(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_42),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_52),
.C(n_51),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_58),
.B(n_52),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_57),
.C(n_39),
.Y(n_60)
);

AOI221xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_5),
.B1(n_14),
.B2(n_40),
.C(n_54),
.Y(n_61)
);


endmodule