module real_aes_7971_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_314;
wire n_252;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
INVx1_ASAP7_75t_L g475 ( .A(n_1), .Y(n_475) );
INVx1_ASAP7_75t_L g188 ( .A(n_2), .Y(n_188) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_3), .A2(n_101), .B1(n_728), .B2(n_737), .C1(n_747), .C2(n_753), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_3), .A2(n_77), .B1(n_741), .B2(n_742), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_3), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_4), .A2(n_38), .B1(n_144), .B2(n_491), .Y(n_501) );
AOI21xp33_ASAP7_75t_L g168 ( .A1(n_5), .A2(n_125), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_6), .B(n_118), .Y(n_466) );
AND2x6_ASAP7_75t_L g130 ( .A(n_7), .B(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_8), .A2(n_227), .B(n_228), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_9), .B(n_39), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_10), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g175 ( .A(n_11), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_12), .B(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g123 ( .A(n_13), .Y(n_123) );
INVx1_ASAP7_75t_L g470 ( .A(n_14), .Y(n_470) );
INVx1_ASAP7_75t_L g233 ( .A(n_15), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_16), .B(n_156), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_17), .B(n_119), .Y(n_447) );
AO32x2_ASAP7_75t_L g499 ( .A1(n_18), .A2(n_118), .A3(n_153), .B1(n_453), .B2(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_19), .B(n_144), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_20), .B(n_139), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_21), .B(n_119), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_22), .A2(n_50), .B1(n_144), .B2(n_491), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_23), .B(n_125), .Y(n_199) );
AOI22xp33_ASAP7_75t_SL g497 ( .A1(n_24), .A2(n_74), .B1(n_144), .B2(n_156), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_25), .B(n_144), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_26), .B(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_27), .A2(n_231), .B(n_232), .C(n_234), .Y(n_230) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_28), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_29), .B(n_177), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_30), .B(n_173), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_31), .A2(n_42), .B1(n_718), .B2(n_719), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_31), .Y(n_718) );
INVx1_ASAP7_75t_L g162 ( .A(n_32), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_33), .B(n_177), .Y(n_514) );
INVx2_ASAP7_75t_L g128 ( .A(n_34), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_35), .B(n_144), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_36), .B(n_177), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_37), .A2(n_130), .B(n_134), .C(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g160 ( .A(n_40), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_41), .B(n_173), .Y(n_243) );
CKINVDCx14_ASAP7_75t_R g719 ( .A(n_42), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_43), .B(n_144), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_44), .A2(n_85), .B1(n_206), .B2(n_491), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_45), .B(n_144), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_46), .B(n_144), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g163 ( .A(n_47), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_48), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_49), .B(n_125), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_51), .A2(n_60), .B1(n_144), .B2(n_156), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g155 ( .A1(n_52), .A2(n_134), .B1(n_156), .B2(n_158), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_53), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_54), .B(n_144), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_55), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_56), .B(n_144), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_57), .A2(n_143), .B(n_172), .C(n_174), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_58), .Y(n_247) );
INVx1_ASAP7_75t_L g170 ( .A(n_59), .Y(n_170) );
INVx1_ASAP7_75t_L g131 ( .A(n_61), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_62), .B(n_144), .Y(n_476) );
INVx1_ASAP7_75t_L g122 ( .A(n_63), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_64), .Y(n_733) );
AO32x2_ASAP7_75t_L g494 ( .A1(n_65), .A2(n_118), .A3(n_213), .B1(n_453), .B2(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g533 ( .A(n_66), .Y(n_533) );
INVx1_ASAP7_75t_L g509 ( .A(n_67), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_SL g138 ( .A1(n_68), .A2(n_139), .B(n_140), .C(n_143), .Y(n_138) );
INVxp67_ASAP7_75t_L g141 ( .A(n_69), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_70), .B(n_156), .Y(n_510) );
INVx1_ASAP7_75t_L g732 ( .A(n_71), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_72), .Y(n_166) );
INVx1_ASAP7_75t_L g240 ( .A(n_73), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_75), .A2(n_130), .B(n_134), .C(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_76), .B(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_77), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_78), .B(n_156), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_79), .B(n_189), .Y(n_202) );
INVx2_ASAP7_75t_L g120 ( .A(n_80), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_81), .B(n_139), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_82), .B(n_156), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_83), .A2(n_130), .B(n_134), .C(n_187), .Y(n_186) );
OR2x2_ASAP7_75t_L g106 ( .A(n_84), .B(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g438 ( .A(n_84), .Y(n_438) );
OR2x2_ASAP7_75t_L g736 ( .A(n_84), .B(n_727), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_86), .A2(n_99), .B1(n_156), .B2(n_157), .Y(n_450) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_87), .A2(n_103), .B1(n_717), .B2(n_720), .C1(n_723), .C2(n_724), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_88), .B(n_177), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_89), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_90), .A2(n_130), .B(n_134), .C(n_216), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_91), .Y(n_223) );
INVx1_ASAP7_75t_L g137 ( .A(n_92), .Y(n_137) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_93), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_94), .B(n_189), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_95), .B(n_156), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_96), .B(n_118), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_97), .A2(n_125), .B(n_132), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_98), .B(n_732), .Y(n_731) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_110), .B1(n_435), .B2(n_439), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g722 ( .A(n_105), .Y(n_722) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g437 ( .A(n_107), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g727 ( .A(n_107), .Y(n_727) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g721 ( .A(n_110), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_110), .A2(n_721), .B1(n_739), .B2(n_740), .Y(n_738) );
AND2x2_ASAP7_75t_SL g110 ( .A(n_111), .B(n_372), .Y(n_110) );
NOR4xp25_ASAP7_75t_L g111 ( .A(n_112), .B(n_302), .C(n_333), .D(n_352), .Y(n_111) );
NAND4xp25_ASAP7_75t_L g112 ( .A(n_113), .B(n_260), .C(n_275), .D(n_293), .Y(n_112) );
AOI222xp33_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_195), .B1(n_236), .B2(n_248), .C1(n_253), .C2(n_255), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_178), .Y(n_114) );
INVx1_ASAP7_75t_L g316 ( .A(n_115), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_149), .Y(n_115) );
AND2x2_ASAP7_75t_L g179 ( .A(n_116), .B(n_167), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_116), .B(n_182), .Y(n_345) );
INVx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g252 ( .A(n_117), .B(n_151), .Y(n_252) );
AND2x2_ASAP7_75t_L g261 ( .A(n_117), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g287 ( .A(n_117), .Y(n_287) );
AND2x2_ASAP7_75t_L g308 ( .A(n_117), .B(n_151), .Y(n_308) );
BUFx2_ASAP7_75t_L g331 ( .A(n_117), .Y(n_331) );
AND2x2_ASAP7_75t_L g355 ( .A(n_117), .B(n_152), .Y(n_355) );
AND2x2_ASAP7_75t_L g419 ( .A(n_117), .B(n_167), .Y(n_419) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_124), .B(n_146), .Y(n_117) );
INVx4_ASAP7_75t_L g148 ( .A(n_118), .Y(n_148) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_118), .A2(n_458), .B(n_466), .Y(n_457) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g153 ( .A(n_119), .Y(n_153) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_120), .B(n_121), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
BUFx2_ASAP7_75t_L g227 ( .A(n_125), .Y(n_227) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_130), .Y(n_125) );
NAND2x1p5_ASAP7_75t_L g164 ( .A(n_126), .B(n_130), .Y(n_164) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVx1_ASAP7_75t_L g465 ( .A(n_127), .Y(n_465) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g135 ( .A(n_128), .Y(n_135) );
INVx1_ASAP7_75t_L g157 ( .A(n_128), .Y(n_157) );
INVx1_ASAP7_75t_L g136 ( .A(n_129), .Y(n_136) );
INVx1_ASAP7_75t_L g139 ( .A(n_129), .Y(n_139) );
INVx3_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_129), .Y(n_159) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_129), .Y(n_173) );
INVx4_ASAP7_75t_SL g145 ( .A(n_130), .Y(n_145) );
BUFx3_ASAP7_75t_L g453 ( .A(n_130), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_130), .A2(n_459), .B(n_462), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_130), .A2(n_469), .B(n_473), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_130), .A2(n_484), .B(n_488), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_130), .A2(n_508), .B(n_511), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_137), .B(n_138), .C(n_145), .Y(n_132) );
O2A1O1Ixp33_ASAP7_75t_L g169 ( .A1(n_133), .A2(n_145), .B(n_170), .C(n_171), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_133), .A2(n_145), .B(n_229), .C(n_230), .Y(n_228) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_135), .Y(n_144) );
BUFx3_ASAP7_75t_L g206 ( .A(n_135), .Y(n_206) );
INVx1_ASAP7_75t_L g491 ( .A(n_135), .Y(n_491) );
INVx1_ASAP7_75t_L g487 ( .A(n_139), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_142), .B(n_175), .Y(n_174) );
INVx5_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g495 ( .A1(n_142), .A2(n_173), .B1(n_496), .B2(n_497), .Y(n_495) );
O2A1O1Ixp5_ASAP7_75t_SL g508 ( .A1(n_143), .A2(n_189), .B(n_509), .C(n_510), .Y(n_508) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_144), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g154 ( .A1(n_145), .A2(n_155), .B1(n_163), .B2(n_164), .Y(n_154) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_147), .A2(n_168), .B(n_176), .Y(n_167) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_SL g208 ( .A(n_148), .B(n_209), .Y(n_208) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_148), .B(n_449), .C(n_453), .Y(n_448) );
AO21x1_ASAP7_75t_L g541 ( .A1(n_148), .A2(n_449), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g320 ( .A(n_149), .B(n_251), .Y(n_320) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_150), .B(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_167), .Y(n_150) );
OR2x2_ASAP7_75t_L g280 ( .A(n_151), .B(n_183), .Y(n_280) );
AND2x2_ASAP7_75t_L g292 ( .A(n_151), .B(n_251), .Y(n_292) );
BUFx2_ASAP7_75t_L g424 ( .A(n_151), .Y(n_424) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OR2x2_ASAP7_75t_L g181 ( .A(n_152), .B(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g274 ( .A(n_152), .B(n_183), .Y(n_274) );
AND2x2_ASAP7_75t_L g327 ( .A(n_152), .B(n_167), .Y(n_327) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_152), .Y(n_363) );
AO21x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_165), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_153), .B(n_166), .Y(n_165) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_153), .A2(n_184), .B(n_192), .Y(n_183) );
INVx2_ASAP7_75t_L g207 ( .A(n_153), .Y(n_207) );
INVx2_ASAP7_75t_L g191 ( .A(n_156), .Y(n_191) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g158 ( .A1(n_159), .A2(n_160), .B1(n_161), .B2(n_162), .Y(n_158) );
INVx2_ASAP7_75t_L g161 ( .A(n_159), .Y(n_161) );
INVx4_ASAP7_75t_L g231 ( .A(n_159), .Y(n_231) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_164), .A2(n_185), .B(n_186), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_164), .A2(n_240), .B(n_241), .Y(n_239) );
AND2x2_ASAP7_75t_L g250 ( .A(n_167), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_SL g262 ( .A(n_167), .Y(n_262) );
INVx2_ASAP7_75t_L g273 ( .A(n_167), .Y(n_273) );
BUFx2_ASAP7_75t_L g297 ( .A(n_167), .Y(n_297) );
AND2x2_ASAP7_75t_SL g354 ( .A(n_167), .B(n_355), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_172), .A2(n_489), .B(n_490), .Y(n_488) );
O2A1O1Ixp5_ASAP7_75t_L g532 ( .A1(n_172), .A2(n_474), .B(n_533), .C(n_534), .Y(n_532) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx4_ASAP7_75t_L g219 ( .A(n_173), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_173), .A2(n_450), .B1(n_451), .B2(n_452), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_173), .A2(n_451), .B1(n_501), .B2(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g194 ( .A(n_177), .Y(n_194) );
INVx2_ASAP7_75t_L g213 ( .A(n_177), .Y(n_213) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_177), .A2(n_226), .B(n_235), .Y(n_225) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_177), .A2(n_483), .B(n_492), .Y(n_482) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_177), .A2(n_507), .B(n_514), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
AOI332xp33_ASAP7_75t_L g275 ( .A1(n_179), .A2(n_276), .A3(n_280), .B1(n_281), .B2(n_285), .B3(n_288), .C1(n_289), .C2(n_291), .Y(n_275) );
NAND2x1_ASAP7_75t_L g360 ( .A(n_179), .B(n_251), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_179), .B(n_265), .Y(n_411) );
A2O1A1Ixp33_ASAP7_75t_SL g293 ( .A1(n_180), .A2(n_294), .B(n_297), .C(n_298), .Y(n_293) );
AND2x2_ASAP7_75t_L g432 ( .A(n_180), .B(n_273), .Y(n_432) );
INVx3_ASAP7_75t_SL g180 ( .A(n_181), .Y(n_180) );
OR2x2_ASAP7_75t_L g329 ( .A(n_181), .B(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g334 ( .A(n_181), .B(n_331), .Y(n_334) );
INVx1_ASAP7_75t_L g265 ( .A(n_182), .Y(n_265) );
AND2x2_ASAP7_75t_L g368 ( .A(n_182), .B(n_327), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_182), .B(n_308), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_182), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_182), .B(n_286), .Y(n_394) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx3_ASAP7_75t_L g251 ( .A(n_183), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .C(n_191), .Y(n_187) );
INVx2_ASAP7_75t_L g451 ( .A(n_189), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_189), .A2(n_460), .B(n_461), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_189), .A2(n_530), .B(n_531), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_191), .A2(n_470), .B(n_471), .C(n_472), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_194), .B(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_194), .B(n_247), .Y(n_246) );
OAI31xp33_ASAP7_75t_L g433 ( .A1(n_195), .A2(n_354), .A3(n_361), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_210), .Y(n_195) );
AND2x2_ASAP7_75t_L g236 ( .A(n_196), .B(n_237), .Y(n_236) );
NAND2x1_ASAP7_75t_SL g256 ( .A(n_196), .B(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_196), .Y(n_343) );
AND2x2_ASAP7_75t_L g348 ( .A(n_196), .B(n_259), .Y(n_348) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_197), .A2(n_261), .B(n_263), .C(n_266), .Y(n_260) );
OR2x2_ASAP7_75t_L g277 ( .A(n_197), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g290 ( .A(n_197), .Y(n_290) );
AND2x2_ASAP7_75t_L g296 ( .A(n_197), .B(n_238), .Y(n_296) );
INVx2_ASAP7_75t_L g314 ( .A(n_197), .Y(n_314) );
AND2x2_ASAP7_75t_L g325 ( .A(n_197), .B(n_279), .Y(n_325) );
AND2x2_ASAP7_75t_L g357 ( .A(n_197), .B(n_315), .Y(n_357) );
AND2x2_ASAP7_75t_L g361 ( .A(n_197), .B(n_284), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_197), .B(n_210), .Y(n_366) );
AND2x2_ASAP7_75t_L g400 ( .A(n_197), .B(n_401), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_197), .B(n_303), .Y(n_434) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_208), .Y(n_197) );
AOI21xp5_ASAP7_75t_SL g198 ( .A1(n_199), .A2(n_200), .B(n_207), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_204), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_204), .A2(n_243), .B(n_244), .Y(n_242) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g234 ( .A(n_206), .Y(n_234) );
INVx1_ASAP7_75t_L g245 ( .A(n_207), .Y(n_245) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_207), .A2(n_468), .B(n_477), .Y(n_467) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_207), .A2(n_528), .B(n_535), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_210), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g342 ( .A(n_210), .Y(n_342) );
AND2x2_ASAP7_75t_L g404 ( .A(n_210), .B(n_325), .Y(n_404) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_224), .Y(n_210) );
OR2x2_ASAP7_75t_L g258 ( .A(n_211), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g268 ( .A(n_211), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_211), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g376 ( .A(n_211), .Y(n_376) );
AND2x2_ASAP7_75t_L g393 ( .A(n_211), .B(n_238), .Y(n_393) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g284 ( .A(n_212), .B(n_224), .Y(n_284) );
AND2x2_ASAP7_75t_L g313 ( .A(n_212), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g324 ( .A(n_212), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_212), .B(n_279), .Y(n_415) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_222), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_221), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_220), .Y(n_216) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g237 ( .A(n_225), .B(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g259 ( .A(n_225), .Y(n_259) );
AND2x2_ASAP7_75t_L g315 ( .A(n_225), .B(n_279), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_231), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g472 ( .A(n_231), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_231), .A2(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g417 ( .A(n_236), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_237), .Y(n_421) );
INVx2_ASAP7_75t_L g279 ( .A(n_238), .Y(n_279) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_245), .B(n_246), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_249), .B(n_252), .Y(n_248) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_250), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_250), .B(n_355), .Y(n_413) );
OR2x2_ASAP7_75t_L g254 ( .A(n_251), .B(n_252), .Y(n_254) );
INVx1_ASAP7_75t_SL g306 ( .A(n_251), .Y(n_306) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AOI221xp5_ASAP7_75t_L g309 ( .A1(n_257), .A2(n_310), .B1(n_312), .B2(n_316), .C(n_317), .Y(n_309) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g337 ( .A(n_258), .B(n_301), .Y(n_337) );
INVx2_ASAP7_75t_L g269 ( .A(n_259), .Y(n_269) );
INVx1_ASAP7_75t_L g295 ( .A(n_259), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_259), .B(n_279), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_259), .B(n_282), .Y(n_389) );
INVx1_ASAP7_75t_L g397 ( .A(n_259), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_261), .B(n_265), .Y(n_311) );
AND2x4_ASAP7_75t_L g286 ( .A(n_262), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g399 ( .A(n_265), .B(n_355), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_267), .B(n_270), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_268), .B(n_300), .Y(n_299) );
INVxp67_ASAP7_75t_L g407 ( .A(n_269), .Y(n_407) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g307 ( .A(n_273), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g379 ( .A(n_273), .B(n_355), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_273), .B(n_292), .Y(n_385) );
AOI322xp5_ASAP7_75t_L g339 ( .A1(n_274), .A2(n_308), .A3(n_315), .B1(n_340), .B2(n_343), .C1(n_344), .C2(n_346), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_274), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g405 ( .A(n_277), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g351 ( .A(n_278), .Y(n_351) );
INVx2_ASAP7_75t_L g282 ( .A(n_279), .Y(n_282) );
INVx1_ASAP7_75t_L g341 ( .A(n_279), .Y(n_341) );
CKINVDCx16_ASAP7_75t_R g288 ( .A(n_280), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g377 ( .A(n_282), .B(n_290), .Y(n_377) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g289 ( .A(n_284), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g332 ( .A(n_284), .B(n_325), .Y(n_332) );
AND2x2_ASAP7_75t_L g336 ( .A(n_284), .B(n_296), .Y(n_336) );
OAI21xp33_ASAP7_75t_SL g346 ( .A1(n_285), .A2(n_347), .B(n_349), .Y(n_346) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_285), .A2(n_417), .B1(n_418), .B2(n_420), .Y(n_416) );
INVx3_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g291 ( .A(n_286), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_286), .B(n_306), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_288), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g428 ( .A(n_295), .Y(n_428) );
INVx4_ASAP7_75t_L g301 ( .A(n_296), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_296), .B(n_323), .Y(n_371) );
INVx1_ASAP7_75t_SL g383 ( .A(n_297), .Y(n_383) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NOR2xp67_ASAP7_75t_L g396 ( .A(n_301), .B(n_397), .Y(n_396) );
OAI211xp5_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_304), .B(n_309), .C(n_326), .Y(n_302) );
OAI221xp5_ASAP7_75t_SL g422 ( .A1(n_304), .A2(n_342), .B1(n_421), .B2(n_423), .C(n_425), .Y(n_422) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_306), .B(n_419), .Y(n_418) );
OAI31xp33_ASAP7_75t_L g398 ( .A1(n_307), .A2(n_384), .A3(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g338 ( .A(n_308), .Y(n_338) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx1_ASAP7_75t_L g388 ( .A(n_313), .Y(n_388) );
AND2x2_ASAP7_75t_L g401 ( .A(n_315), .B(n_324), .Y(n_401) );
AOI21xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B(n_321), .Y(n_317) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVxp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_325), .B(n_428), .Y(n_427) );
OAI21xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_328), .B(n_332), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI221xp5_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_335), .B1(n_337), .B2(n_338), .C(n_339), .Y(n_333) );
A2O1A1Ixp33_ASAP7_75t_L g402 ( .A1(n_334), .A2(n_403), .B(n_405), .C(n_408), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_337), .B(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g364 ( .A(n_345), .Y(n_364) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g350 ( .A(n_348), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g392 ( .A(n_348), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OAI211xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_356), .B(n_358), .C(n_367), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_356), .A2(n_366), .B1(n_430), .B2(n_431), .C(n_433), .Y(n_429) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B1(n_362), .B2(n_365), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI21xp5_ASAP7_75t_SL g367 ( .A1(n_368), .A2(n_369), .B(n_370), .Y(n_367) );
INVx1_ASAP7_75t_SL g430 ( .A(n_369), .Y(n_430) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR4xp25_ASAP7_75t_L g372 ( .A(n_373), .B(n_402), .C(n_422), .D(n_429), .Y(n_372) );
OAI211xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_378), .B(n_380), .C(n_398), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_384), .B(n_386), .C(n_390), .Y(n_380) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g409 ( .A(n_387), .Y(n_409) );
OR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
OR2x2_ASAP7_75t_L g420 ( .A(n_388), .B(n_421), .Y(n_420) );
OAI21xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_394), .B(n_395), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_412), .B2(n_414), .C(n_416), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_419), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI22x1_ASAP7_75t_SL g720 ( .A1(n_437), .A2(n_440), .B1(n_721), .B2(n_722), .Y(n_720) );
NOR2x2_ASAP7_75t_L g726 ( .A(n_438), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_SL g441 ( .A(n_442), .B(n_651), .Y(n_441) );
NOR5xp2_ASAP7_75t_L g442 ( .A(n_443), .B(n_564), .C(n_610), .D(n_623), .E(n_635), .Y(n_442) );
OAI211xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_478), .B(n_518), .C(n_545), .Y(n_443) );
INVx1_ASAP7_75t_SL g646 ( .A(n_444), .Y(n_646) );
OR2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_454), .Y(n_444) );
AND2x2_ASAP7_75t_L g570 ( .A(n_445), .B(n_455), .Y(n_570) );
AND2x2_ASAP7_75t_L g598 ( .A(n_445), .B(n_544), .Y(n_598) );
AND2x2_ASAP7_75t_L g606 ( .A(n_445), .B(n_549), .Y(n_606) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g536 ( .A(n_446), .B(n_456), .Y(n_536) );
INVx2_ASAP7_75t_L g548 ( .A(n_446), .Y(n_548) );
AND2x2_ASAP7_75t_L g673 ( .A(n_446), .B(n_615), .Y(n_673) );
OR2x2_ASAP7_75t_L g675 ( .A(n_446), .B(n_676), .Y(n_675) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g542 ( .A(n_447), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_451), .A2(n_463), .B(n_464), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_451), .A2(n_474), .B(n_475), .C(n_476), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_453), .A2(n_529), .B(n_532), .Y(n_528) );
INVx2_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g586 ( .A(n_455), .B(n_558), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_455), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g700 ( .A(n_455), .B(n_540), .Y(n_700) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_467), .Y(n_455) );
AND2x2_ASAP7_75t_L g543 ( .A(n_456), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g590 ( .A(n_456), .Y(n_590) );
AND2x2_ASAP7_75t_L g615 ( .A(n_456), .B(n_527), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_456), .B(n_648), .Y(n_685) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g549 ( .A(n_457), .B(n_527), .Y(n_549) );
AND2x2_ASAP7_75t_L g563 ( .A(n_457), .B(n_526), .Y(n_563) );
AND2x2_ASAP7_75t_L g580 ( .A(n_457), .B(n_467), .Y(n_580) );
AND2x2_ASAP7_75t_L g637 ( .A(n_457), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_457), .B(n_544), .Y(n_650) );
AND2x2_ASAP7_75t_L g702 ( .A(n_457), .B(n_627), .Y(n_702) );
INVx2_ASAP7_75t_L g474 ( .A(n_465), .Y(n_474) );
AND2x2_ASAP7_75t_L g525 ( .A(n_467), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g544 ( .A(n_467), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_467), .B(n_527), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_503), .B(n_515), .Y(n_478) );
INVx1_ASAP7_75t_SL g634 ( .A(n_479), .Y(n_634) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_493), .Y(n_479) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_SL g522 ( .A(n_481), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g517 ( .A(n_482), .Y(n_517) );
INVx1_ASAP7_75t_L g554 ( .A(n_482), .Y(n_554) );
AND2x2_ASAP7_75t_L g575 ( .A(n_482), .B(n_498), .Y(n_575) );
AND2x2_ASAP7_75t_L g609 ( .A(n_482), .B(n_499), .Y(n_609) );
OR2x2_ASAP7_75t_L g628 ( .A(n_482), .B(n_505), .Y(n_628) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_482), .Y(n_642) );
AND2x2_ASAP7_75t_L g655 ( .A(n_482), .B(n_656), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_487), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_493), .A2(n_577), .B1(n_578), .B2(n_587), .Y(n_576) );
AND2x2_ASAP7_75t_L g660 ( .A(n_493), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_498), .Y(n_493) );
INVx1_ASAP7_75t_L g521 ( .A(n_494), .Y(n_521) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_494), .Y(n_558) );
INVx1_ASAP7_75t_L g569 ( .A(n_494), .Y(n_569) );
AND2x2_ASAP7_75t_L g584 ( .A(n_494), .B(n_499), .Y(n_584) );
OR2x2_ASAP7_75t_L g538 ( .A(n_498), .B(n_523), .Y(n_538) );
AND2x2_ASAP7_75t_L g568 ( .A(n_498), .B(n_569), .Y(n_568) );
NOR2xp67_ASAP7_75t_L g656 ( .A(n_498), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g516 ( .A(n_499), .B(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g625 ( .A(n_499), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_503), .B(n_641), .Y(n_640) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g603 ( .A(n_504), .B(n_569), .Y(n_603) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g515 ( .A(n_505), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g574 ( .A(n_505), .Y(n_574) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g523 ( .A(n_506), .Y(n_523) );
OR2x2_ASAP7_75t_L g553 ( .A(n_506), .B(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_506), .Y(n_608) );
AOI32xp33_ASAP7_75t_L g645 ( .A1(n_515), .A2(n_575), .A3(n_646), .B1(n_647), .B2(n_649), .Y(n_645) );
AND2x2_ASAP7_75t_L g571 ( .A(n_516), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_516), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_516), .B(n_603), .Y(n_689) );
INVx1_ASAP7_75t_L g694 ( .A(n_516), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_524), .B1(n_537), .B2(n_539), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .Y(n_519) );
AND2x2_ASAP7_75t_L g624 ( .A(n_520), .B(n_625), .Y(n_624) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_521), .B(n_523), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_522), .A2(n_546), .B1(n_550), .B2(n_560), .Y(n_545) );
AND2x2_ASAP7_75t_L g567 ( .A(n_522), .B(n_568), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g618 ( .A1(n_522), .A2(n_536), .B(n_584), .C(n_619), .Y(n_618) );
OAI332xp33_ASAP7_75t_L g623 ( .A1(n_522), .A2(n_624), .A3(n_626), .B1(n_628), .B2(n_629), .B3(n_631), .C1(n_632), .C2(n_634), .Y(n_623) );
INVx2_ASAP7_75t_L g664 ( .A(n_522), .Y(n_664) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_523), .Y(n_582) );
INVx1_ASAP7_75t_L g657 ( .A(n_523), .Y(n_657) );
AND2x2_ASAP7_75t_L g711 ( .A(n_523), .B(n_575), .Y(n_711) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_536), .Y(n_524) );
AND2x2_ASAP7_75t_L g591 ( .A(n_526), .B(n_541), .Y(n_591) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g540 ( .A(n_527), .B(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g639 ( .A(n_527), .B(n_541), .Y(n_639) );
INVx1_ASAP7_75t_L g648 ( .A(n_527), .Y(n_648) );
INVx1_ASAP7_75t_L g622 ( .A(n_536), .Y(n_622) );
INVxp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g706 ( .A(n_538), .B(n_558), .Y(n_706) );
INVx1_ASAP7_75t_SL g617 ( .A(n_539), .Y(n_617) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .Y(n_539) );
AND2x2_ASAP7_75t_L g644 ( .A(n_540), .B(n_602), .Y(n_644) );
INVx1_ASAP7_75t_L g663 ( .A(n_540), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_540), .B(n_630), .Y(n_665) );
INVx1_ASAP7_75t_L g562 ( .A(n_541), .Y(n_562) );
AND2x2_ASAP7_75t_L g566 ( .A(n_543), .B(n_547), .Y(n_566) );
AND2x2_ASAP7_75t_L g633 ( .A(n_543), .B(n_591), .Y(n_633) );
INVx2_ASAP7_75t_L g676 ( .A(n_543), .Y(n_676) );
INVx2_ASAP7_75t_L g559 ( .A(n_544), .Y(n_559) );
AND2x2_ASAP7_75t_L g561 ( .A(n_544), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
INVx1_ASAP7_75t_L g577 ( .A(n_547), .Y(n_577) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_548), .B(n_621), .Y(n_627) );
OR2x2_ASAP7_75t_L g691 ( .A(n_548), .B(n_650), .Y(n_691) );
INVx1_ASAP7_75t_L g715 ( .A(n_548), .Y(n_715) );
INVx1_ASAP7_75t_L g671 ( .A(n_549), .Y(n_671) );
AND2x2_ASAP7_75t_L g716 ( .A(n_549), .B(n_559), .Y(n_716) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_553), .A2(n_579), .B1(n_581), .B2(n_585), .Y(n_578) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI322xp33_ASAP7_75t_SL g662 ( .A1(n_556), .A2(n_663), .A3(n_664), .B1(n_665), .B2(n_666), .C1(n_669), .C2(n_671), .Y(n_662) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
AND2x2_ASAP7_75t_L g659 ( .A(n_557), .B(n_575), .Y(n_659) );
OR2x2_ASAP7_75t_L g693 ( .A(n_557), .B(n_694), .Y(n_693) );
OR2x2_ASAP7_75t_L g696 ( .A(n_557), .B(n_628), .Y(n_696) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g641 ( .A(n_558), .B(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g697 ( .A(n_558), .B(n_628), .Y(n_697) );
INVx3_ASAP7_75t_L g630 ( .A(n_559), .Y(n_630) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
INVx1_ASAP7_75t_L g686 ( .A(n_561), .Y(n_686) );
AOI222xp33_ASAP7_75t_L g565 ( .A1(n_563), .A2(n_566), .B1(n_567), .B2(n_570), .C1(n_571), .C2(n_573), .Y(n_565) );
INVx1_ASAP7_75t_L g596 ( .A(n_563), .Y(n_596) );
NAND3xp33_ASAP7_75t_SL g564 ( .A(n_565), .B(n_576), .C(n_593), .Y(n_564) );
AND2x2_ASAP7_75t_L g681 ( .A(n_568), .B(n_582), .Y(n_681) );
BUFx2_ASAP7_75t_L g572 ( .A(n_569), .Y(n_572) );
INVx1_ASAP7_75t_L g613 ( .A(n_569), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_570), .A2(n_606), .B1(n_659), .B2(n_660), .C(n_662), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_572), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_575), .Y(n_599) );
AND2x2_ASAP7_75t_L g612 ( .A(n_575), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_580), .B(n_591), .Y(n_592) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
OAI21xp33_ASAP7_75t_L g587 ( .A1(n_582), .A2(n_588), .B(n_592), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_582), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g679 ( .A(n_584), .B(n_661), .Y(n_679) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g602 ( .A(n_590), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_591), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g708 ( .A(n_591), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_599), .B1(n_600), .B2(n_603), .C(n_604), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_595), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g704 ( .A(n_603), .B(n_609), .Y(n_704) );
INVxp67_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
OAI31xp33_ASAP7_75t_SL g672 ( .A1(n_607), .A2(n_646), .A3(n_673), .B(n_674), .Y(n_672) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g661 ( .A(n_608), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_609), .B(n_613), .Y(n_712) );
OAI221xp5_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_614), .B1(n_616), .B2(n_617), .C(n_618), .Y(n_610) );
INVx1_ASAP7_75t_L g616 ( .A(n_612), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_615), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g631 ( .A(n_624), .Y(n_631) );
INVx2_ASAP7_75t_L g667 ( .A(n_625), .Y(n_667) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g653 ( .A(n_630), .B(n_639), .Y(n_653) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_630), .A2(n_647), .B(n_704), .C(n_705), .Y(n_703) );
OAI221xp5_ASAP7_75t_SL g635 ( .A1(n_631), .A2(n_636), .B1(n_640), .B2(n_643), .C(n_645), .Y(n_635) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_634), .A2(n_699), .B(n_701), .C(n_703), .Y(n_698) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_637), .A2(n_688), .B1(n_690), .B2(n_692), .C(n_695), .Y(n_687) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
NOR4xp25_ASAP7_75t_L g651 ( .A(n_652), .B(n_677), .C(n_698), .D(n_709), .Y(n_651) );
OAI211xp5_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B(n_658), .C(n_672), .Y(n_652) );
INVx1_ASAP7_75t_SL g707 ( .A(n_659), .Y(n_707) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_SL g670 ( .A(n_668), .Y(n_670) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_675), .A2(n_684), .B1(n_696), .B2(n_697), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B(n_682), .C(n_687), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AOI31xp33_ASAP7_75t_L g709 ( .A1(n_680), .A2(n_710), .A3(n_712), .B(n_713), .Y(n_709) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g723 ( .A(n_717), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_734), .Y(n_729) );
NOR2xp33_ASAP7_75t_SL g730 ( .A(n_731), .B(n_733), .Y(n_730) );
INVx1_ASAP7_75t_SL g752 ( .A(n_731), .Y(n_752) );
INVx1_ASAP7_75t_L g751 ( .A(n_733), .Y(n_751) );
OA21x2_ASAP7_75t_L g754 ( .A1(n_733), .A2(n_752), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g743 ( .A(n_734), .Y(n_743) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_736), .Y(n_746) );
BUFx2_ASAP7_75t_L g755 ( .A(n_736), .Y(n_755) );
OAI21xp5_ASAP7_75t_SL g737 ( .A1(n_738), .A2(n_743), .B(n_744), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
endmodule