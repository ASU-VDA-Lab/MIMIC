module fake_jpeg_4143_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_17),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_32),
.B1(n_24),
.B2(n_21),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_62),
.B1(n_70),
.B2(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_66),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_57),
.B(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_59),
.B(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_24),
.B1(n_33),
.B2(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_26),
.B1(n_20),
.B2(n_22),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_32),
.B1(n_21),
.B2(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_71),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_39),
.A2(n_21),
.B1(n_33),
.B2(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_36),
.A2(n_21),
.B1(n_25),
.B2(n_23),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_23),
.B1(n_25),
.B2(n_19),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_75),
.A2(n_77),
.B1(n_80),
.B2(n_81),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_80),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_77),
.B(n_87),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_78),
.A2(n_88),
.B1(n_90),
.B2(n_51),
.Y(n_106)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_36),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_84),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_48),
.B1(n_46),
.B2(n_45),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_51),
.B1(n_69),
.B2(n_50),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_57),
.B1(n_52),
.B2(n_72),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_48),
.B1(n_46),
.B2(n_45),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_20),
.B1(n_29),
.B2(n_22),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_26),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_96),
.Y(n_128)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_27),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_27),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_42),
.Y(n_124)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_99),
.Y(n_126)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_103),
.B(n_108),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_104),
.A2(n_109),
.B1(n_113),
.B2(n_81),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_42),
.B(n_29),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_140)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_51),
.B1(n_69),
.B2(n_50),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_89),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_82),
.Y(n_134)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_71),
.C(n_67),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_18),
.Y(n_151)
);

AO22x1_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_41),
.B1(n_37),
.B2(n_30),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_125),
.A2(n_103),
.B1(n_106),
.B2(n_110),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_85),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_137),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_143),
.B1(n_151),
.B2(n_155),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_134),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_126),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_97),
.C(n_96),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_18),
.C(n_31),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_129),
.A2(n_120),
.B1(n_122),
.B2(n_108),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_82),
.B(n_19),
.Y(n_146)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_146),
.B(n_104),
.CI(n_109),
.CON(n_161),
.SN(n_161)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_114),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_86),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_152),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_90),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_153),
.B(n_117),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_27),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_18),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_113),
.A2(n_100),
.B1(n_99),
.B2(n_68),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_101),
.A2(n_102),
.B(n_111),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_130),
.B(n_27),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_102),
.A2(n_100),
.B1(n_99),
.B2(n_68),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_167),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_123),
.B1(n_115),
.B2(n_112),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_163),
.A2(n_176),
.B1(n_183),
.B2(n_145),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_171),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_170),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_158),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_173),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_146),
.B(n_118),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_135),
.A2(n_56),
.B1(n_127),
.B2(n_37),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_141),
.B(n_0),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_177),
.A2(n_147),
.B(n_137),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_178),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_180),
.A2(n_31),
.B(n_30),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_31),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_185),
.C(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_18),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_153),
.B(n_107),
.Y(n_210)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

INVxp33_ASAP7_75t_SL g231 ( 
.A(n_188),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_149),
.B1(n_132),
.B2(n_142),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_191),
.A2(n_211),
.B1(n_215),
.B2(n_167),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_144),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_197),
.C(n_201),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_143),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_199),
.B(n_206),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_149),
.Y(n_201)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_151),
.B(n_131),
.C(n_31),
.D(n_41),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_210),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_151),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_209),
.C(n_180),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_210),
.Y(n_224)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_183),
.A2(n_166),
.B(n_160),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_212),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_158),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_214),
.B1(n_170),
.B2(n_168),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_186),
.A2(n_145),
.B1(n_119),
.B2(n_136),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_136),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_186),
.A2(n_119),
.B1(n_30),
.B2(n_2),
.Y(n_215)
);

HB1xp67_ASAP7_75t_SL g216 ( 
.A(n_212),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_235),
.B(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_218),
.Y(n_250)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_198),
.A2(n_176),
.B1(n_160),
.B2(n_172),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_219),
.A2(n_221),
.B1(n_238),
.B2(n_239),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_184),
.B1(n_161),
.B2(n_174),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_223),
.A2(n_240),
.B1(n_189),
.B2(n_193),
.Y(n_257)
);

OAI211xp5_ASAP7_75t_L g256 ( 
.A1(n_224),
.A2(n_242),
.B(n_223),
.C(n_231),
.Y(n_256)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_192),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_165),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_196),
.Y(n_247)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_230),
.Y(n_255)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_194),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_236),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_209),
.C(n_204),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_213),
.A2(n_164),
.B1(n_162),
.B2(n_161),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_194),
.A2(n_173),
.B1(n_179),
.B2(n_161),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_191),
.A2(n_179),
.B1(n_177),
.B2(n_169),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_208),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_201),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_247),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_246),
.A2(n_1),
.B(n_2),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_252),
.C(n_258),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_223),
.A2(n_189),
.B(n_195),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_228),
.B(n_224),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_202),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_205),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_220),
.Y(n_268)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_264),
.B1(n_1),
.B2(n_2),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_206),
.C(n_203),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_203),
.C(n_119),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_265),
.C(n_263),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_218),
.A2(n_223),
.B1(n_225),
.B2(n_241),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_0),
.C(n_1),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_238),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_266),
.B(n_270),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_284),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_269),
.A2(n_274),
.B(n_277),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_258),
.B(n_240),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_259),
.A2(n_235),
.B1(n_219),
.B2(n_220),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_280),
.B1(n_251),
.B2(n_261),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_260),
.C(n_265),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_275),
.A2(n_276),
.B1(n_255),
.B2(n_262),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_245),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_250),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_250),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_283),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_259),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_3),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_246),
.Y(n_282)
);

INVxp33_ASAP7_75t_SL g294 ( 
.A(n_282),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_10),
.C(n_15),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_244),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_288),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_252),
.Y(n_288)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_248),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_292),
.C(n_298),
.Y(n_306)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_274),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_299),
.B1(n_300),
.B2(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_243),
.C(n_253),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_278),
.A2(n_243),
.B1(n_10),
.B2(n_11),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_301),
.B(n_303),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_294),
.B(n_271),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_314),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_273),
.B(n_267),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_309),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_290),
.B(n_275),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_300),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_284),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_310),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_276),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_281),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_10),
.B(n_15),
.Y(n_311)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_311),
.A2(n_12),
.B(n_15),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_5),
.C(n_6),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_7),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_285),
.B(n_288),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_319),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_318),
.B(n_323),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_305),
.A2(n_296),
.B1(n_293),
.B2(n_285),
.Y(n_319)
);

NAND2xp33_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_296),
.Y(n_320)
);

NOR2x1_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_16),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_306),
.A2(n_312),
.B1(n_314),
.B2(n_313),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_13),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_16),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_306),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_327),
.A2(n_329),
.B(n_330),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_313),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_316),
.A2(n_9),
.B(n_11),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_13),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_331),
.A2(n_7),
.B(n_8),
.Y(n_334)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_332),
.A2(n_7),
.B(n_8),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_333),
.B(n_334),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_315),
.Y(n_335)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_335),
.Y(n_339)
);

AOI21x1_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_321),
.B(n_337),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_340),
.B(n_325),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_325),
.B(n_338),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_336),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_8),
.Y(n_344)
);


endmodule