module real_jpeg_13689_n_17 (n_5, n_4, n_8, n_0, n_12, n_299, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_299;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_249;
wire n_288;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_184;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_65;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_240;
wire n_55;
wire n_185;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_202;
wire n_295;
wire n_167;
wire n_179;
wire n_133;
wire n_216;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_3),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_42),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_3),
.A2(n_42),
.B1(n_60),
.B2(n_62),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_59),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_59),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_8),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_8),
.A2(n_60),
.B1(n_62),
.B2(n_85),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_85),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_85),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_9),
.A2(n_60),
.B1(n_62),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_9),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_151),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_151),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_9),
.A2(n_39),
.B1(n_40),
.B2(n_151),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_10),
.A2(n_60),
.B1(n_62),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_10),
.B(n_29),
.C(n_65),
.Y(n_143)
);

NAND2x1_ASAP7_75t_SL g147 ( 
.A(n_10),
.B(n_83),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_10),
.A2(n_95),
.B(n_155),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_10),
.A2(n_44),
.B(n_82),
.C(n_182),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_139),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_10),
.B(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_10),
.B(n_39),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_11),
.A2(n_35),
.B1(n_60),
.B2(n_62),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_12),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g240 ( 
.A(n_12),
.B(n_45),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_13),
.A2(n_53),
.B1(n_60),
.B2(n_62),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_53),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_14),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_104),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_14),
.A2(n_60),
.B1(n_62),
.B2(n_104),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_104),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_15),
.A2(n_60),
.B1(n_62),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_15),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_70),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_70),
.Y(n_115)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_126),
.B1(n_296),
.B2(n_297),
.Y(n_18)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_19),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_124),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_107),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_21),
.B(n_107),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_73),
.C(n_89),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_22),
.A2(n_23),
.B1(n_73),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_55),
.B2(n_72),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_36),
.B1(n_37),
.B2(n_54),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_26),
.A2(n_37),
.B(n_72),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_26),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.Y(n_26)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_27),
.A2(n_32),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_27),
.B(n_156),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_27),
.A2(n_32),
.B1(n_94),
.B2(n_244),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_28),
.A2(n_29),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_28),
.B(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_32),
.B(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_34),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_92)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B(n_47),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_38),
.A2(n_43),
.B1(n_49),
.B2(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_40),
.A2(n_49),
.B(n_139),
.C(n_226),
.Y(n_225)
);

AOI32xp33_ASAP7_75t_L g239 ( 
.A1(n_40),
.A2(n_44),
.A3(n_46),
.B1(n_227),
.B2(n_240),
.Y(n_239)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_43),
.B(n_52),
.Y(n_106)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_43),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_43),
.A2(n_47),
.B(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_43),
.A2(n_49),
.B1(n_103),
.B2(n_254),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_44),
.A2(n_45),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_49),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_63),
.B1(n_68),
.B2(n_71),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_63),
.B1(n_71),
.B2(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_60),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

AO22x1_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_62),
.B1(n_81),
.B2(n_82),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_60),
.B(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_62),
.A2(n_81),
.B(n_139),
.Y(n_182)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_63),
.A2(n_71),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_63),
.B(n_141),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_63),
.A2(n_71),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_63),
.A2(n_71),
.B1(n_99),
.B2(n_233),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_69),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_67),
.A2(n_150),
.B(n_152),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_67),
.B(n_139),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_67),
.A2(n_152),
.B(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_71),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_73),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B(n_88),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_77),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_SL g137 ( 
.A1(n_75),
.A2(n_138),
.B(n_140),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_75),
.A2(n_140),
.B(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_84),
.B1(n_86),
.B2(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_78),
.A2(n_187),
.B(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_78),
.A2(n_86),
.B1(n_202),
.B2(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_78),
.A2(n_188),
.B(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_83),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_79),
.B(n_189),
.Y(n_203)
);

NOR2x1_ASAP7_75t_R g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_83),
.B(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_86),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_86),
.A2(n_101),
.B(n_203),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_89),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.C(n_102),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_90),
.A2(n_91),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_92),
.A2(n_97),
.B1(n_98),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_92),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_95),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_95),
.A2(n_96),
.B1(n_184),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_95),
.A2(n_96),
.B1(n_210),
.B2(n_243),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_96),
.A2(n_161),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_96),
.B(n_139),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_96),
.A2(n_169),
.B(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_100),
.B(n_102),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_106),
.B(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_110)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_126),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_290),
.B(n_295),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_278),
.B(n_289),
.Y(n_128)
);

OAI321xp33_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_246),
.A3(n_271),
.B1(n_276),
.B2(n_277),
.C(n_299),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_219),
.B(n_245),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_196),
.B(n_218),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_177),
.B(n_195),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_157),
.B(n_176),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_135),
.B(n_144),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_137),
.B1(n_142),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_142),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_149),
.C(n_153),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_154),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_165),
.B(n_175),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_163),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_170),
.B(n_174),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_167),
.B(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_178),
.B(n_179),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_185),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_190),
.C(n_194),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_183),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_185)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_192),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_197),
.B(n_198),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_211),
.B2(n_212),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_214),
.C(n_216),
.Y(n_220)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_205),
.C(n_209),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_220),
.B(n_221),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_235),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_236),
.C(n_237),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_228),
.B2(n_234),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_229),
.C(n_231),
.Y(n_260)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_242),
.Y(n_256)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_261),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_261),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_257),
.C(n_260),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_248),
.A2(n_249),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_256),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_255),
.C(n_256),
.Y(n_270)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_253),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_260),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_259),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_270),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_265),
.C(n_270),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_269),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_268),
.C(n_269),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_288),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_288),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_283),
.C(n_284),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);


endmodule