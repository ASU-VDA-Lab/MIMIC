module fake_jpeg_24353_n_35 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

MAJIxp5_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_2),
.C(n_4),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

NOR2x1_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_20),
.Y(n_24)
);

AOI32xp33_ASAP7_75t_L g15 ( 
.A1(n_10),
.A2(n_0),
.A3(n_1),
.B1(n_3),
.B2(n_6),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_15),
.A2(n_17),
.B1(n_18),
.B2(n_14),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_13),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_7),
.C(n_11),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_20),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_29),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_21),
.C(n_26),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_25),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_23),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_30),
.C(n_32),
.Y(n_35)
);


endmodule