module fake_jpeg_3100_n_99 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_99);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_99;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_24),
.B(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx2_ASAP7_75t_SL g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g28 ( 
.A1(n_15),
.A2(n_0),
.B(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_11),
.B1(n_20),
.B2(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_43),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_25),
.B1(n_26),
.B2(n_23),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_29),
.B1(n_34),
.B2(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_13),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_22),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_57),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_68)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_61),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_44),
.C(n_42),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_61),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_72),
.B1(n_61),
.B2(n_52),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_41),
.B(n_27),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_41),
.B1(n_47),
.B2(n_0),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_74),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_79),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_80),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_63),
.C(n_66),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_68),
.C(n_62),
.Y(n_89)
);

AOI22x1_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_69),
.B1(n_72),
.B2(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

A2O1A1O1Ixp25_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_50),
.B(n_65),
.C(n_71),
.D(n_53),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_88),
.B(n_89),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_51),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_93),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_83),
.C(n_84),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_86),
.C(n_64),
.Y(n_95)
);

AOI31xp67_ASAP7_75t_SL g96 ( 
.A1(n_95),
.A2(n_86),
.A3(n_73),
.B(n_94),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_96),
.B(n_73),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_8),
.C(n_9),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_0),
.Y(n_99)
);


endmodule