module real_jpeg_24452_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx6_ASAP7_75t_L g102 ( 
.A(n_0),
.Y(n_102)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_0),
.Y(n_132)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_0),
.Y(n_202)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_0),
.Y(n_285)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_2),
.A2(n_40),
.B1(n_64),
.B2(n_67),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_47),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_47),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_3),
.A2(n_47),
.B1(n_64),
.B2(n_67),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_7),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_7),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_88),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_88),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_7),
.A2(n_64),
.B1(n_67),
.B2(n_88),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_55),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_55),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_8),
.A2(n_55),
.B1(n_64),
.B2(n_67),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_11),
.A2(n_57),
.B1(n_87),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_11),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_117),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_117),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_11),
.A2(n_64),
.B1(n_67),
.B2(n_117),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_13),
.A2(n_46),
.B1(n_86),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_13),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_171),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_171),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_13),
.A2(n_64),
.B1(n_67),
.B2(n_171),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_14),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_142),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_142),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_14),
.A2(n_64),
.B1(n_67),
.B2(n_142),
.Y(n_282)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_15),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_15),
.B(n_53),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_15),
.B(n_28),
.C(n_30),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_195),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_15),
.B(n_37),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_195),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_15),
.B(n_64),
.C(n_66),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_15),
.A2(n_101),
.B(n_283),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_16),
.A2(n_45),
.B1(n_57),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_16),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_77),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_16),
.A2(n_27),
.B1(n_28),
.B2(n_77),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_16),
.A2(n_64),
.B1(n_67),
.B2(n_77),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_95),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_94),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_21),
.B(n_78),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_60),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_41),
.B1(n_58),
.B2(n_59),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_37),
.B(n_38),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_24),
.A2(n_37),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_24),
.B(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_24),
.A2(n_37),
.B1(n_189),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_25),
.A2(n_26),
.B1(n_39),
.B2(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_25),
.A2(n_26),
.B1(n_92),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_25),
.A2(n_26),
.B1(n_121),
.B2(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_25),
.A2(n_188),
.B(n_190),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_25),
.A2(n_190),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_26),
.A2(n_138),
.B(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_26),
.A2(n_174),
.B(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_27),
.A2(n_28),
.B1(n_65),
.B2(n_66),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_28),
.B(n_292),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_34),
.B1(n_50),
.B2(n_51),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_SL g196 ( 
.A(n_33),
.B(n_45),
.C(n_51),
.Y(n_196)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_34),
.A2(n_50),
.B(n_194),
.C(n_196),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_34),
.B(n_248),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_37),
.B(n_175),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_52),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_48),
.A2(n_53),
.B1(n_141),
.B2(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_48),
.A2(n_144),
.B(n_194),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_75),
.B1(n_76),
.B2(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_84),
.B(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_52),
.B(n_116),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_52),
.A2(n_114),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_72),
.C(n_74),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_72),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_83),
.C(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_61),
.A2(n_82),
.B1(n_90),
.B2(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_68),
.B(n_70),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_62),
.A2(n_68),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_62),
.A2(n_68),
.B1(n_108),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_62),
.A2(n_68),
.B1(n_255),
.B2(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_62),
.B(n_222),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_63),
.A2(n_71),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_63),
.A2(n_123),
.B1(n_136),
.B2(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_63),
.A2(n_181),
.B(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_63),
.A2(n_221),
.B(n_256),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_63),
.B(n_195),
.Y(n_304)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_63)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_67),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_68),
.B(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_75),
.A2(n_140),
.B(n_143),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.C(n_89),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_79),
.A2(n_83),
.B1(n_154),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_79),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_83),
.A2(n_151),
.B1(n_152),
.B2(n_154),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_83),
.Y(n_154)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

HAxp5_ASAP7_75t_SL g194 ( 
.A(n_87),
.B(n_195),
.CON(n_194),
.SN(n_194)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_89),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI31xp33_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_155),
.A3(n_161),
.B(n_345),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_145),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_97),
.B(n_145),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_118),
.C(n_126),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_98),
.A2(n_118),
.B1(n_119),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_98),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_110),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_99),
.A2(n_100),
.B(n_112),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_106),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_100),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_100),
.A2(n_106),
.B1(n_107),
.B2(n_111),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B(n_105),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_101),
.A2(n_105),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_101),
.A2(n_103),
.B1(n_131),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_101),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_101),
.A2(n_200),
.B1(n_202),
.B2(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_101),
.B(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_101),
.A2(n_282),
.B(n_283),
.Y(n_281)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_122),
.B(n_125),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_122),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_123),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_123),
.A2(n_271),
.B(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_126),
.A2(n_127),
.B1(n_340),
.B2(n_342),
.Y(n_339)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_137),
.C(n_139),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_128),
.A2(n_129),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_130),
.A2(n_133),
.B1(n_134),
.B2(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_130),
.Y(n_183)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_132),
.Y(n_298)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_137),
.B(n_139),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_148),
.C(n_150),
.Y(n_160)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_156),
.A2(n_346),
.B(n_347),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_157),
.B(n_160),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_338),
.B(n_344),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_210),
.B(n_337),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_203),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_164),
.B(n_203),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_182),
.C(n_184),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_165),
.A2(n_166),
.B1(n_182),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_176),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_172),
.B2(n_173),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_172),
.C(n_176),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_170),
.Y(n_186)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_177),
.B(n_180),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_197)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_182),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_184),
.B(n_334),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_191),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_185),
.B(n_187),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_191),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_193),
.B1(n_197),
.B2(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_195),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_198),
.A2(n_296),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_202),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_205),
.B(n_206),
.C(n_209),
.Y(n_343)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_240),
.B(n_331),
.C(n_336),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_234),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_234),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_224),
.C(n_227),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_213),
.A2(n_214),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_223),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_219),
.C(n_223),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_218),
.Y(n_229)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_227),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.C(n_232),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_265),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_235),
.B(n_238),
.C(n_239),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_324),
.B(n_330),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_272),
.B(n_323),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_261),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_245),
.B(n_261),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_254),
.C(n_258),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_246),
.B(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_249),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B(n_252),
.Y(n_249)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_252),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_253),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_254),
.A2(n_258),
.B1(n_259),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_254),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_257),
.Y(n_270)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_266),
.B2(n_267),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_262),
.B(n_268),
.C(n_269),
.Y(n_329)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_317),
.B(n_322),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_293),
.B(n_316),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_287),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_275),
.B(n_287),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_277),
.B(n_280),
.C(n_281),
.Y(n_321)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_285),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_302),
.B(n_315),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_300),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_300),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_308),
.B(n_314),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_305),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_313),
.Y(n_308)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_321),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_321),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_329),
.Y(n_330)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_333),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_339),
.B(n_343),
.Y(n_344)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_340),
.Y(n_342)
);


endmodule