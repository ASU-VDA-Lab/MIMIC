module fake_jpeg_24211_n_132 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_11),
.B(n_2),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_37),
.Y(n_46)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_39),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_38),
.B1(n_28),
.B2(n_21),
.Y(n_55)
);

CKINVDCx6p67_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_1),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_21),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_61),
.Y(n_73)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_50),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_54),
.B1(n_30),
.B2(n_47),
.Y(n_76)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_29),
.A2(n_22),
.B1(n_15),
.B2(n_13),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_22),
.B1(n_28),
.B2(n_14),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_68),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_29),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_77),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_69),
.B(n_26),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_33),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_74),
.C(n_78),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_35),
.C(n_41),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_79),
.C(n_47),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_55),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_17),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_7),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_50),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

AO22x1_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_59),
.B1(n_58),
.B2(n_50),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_59),
.B1(n_80),
.B2(n_71),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_68),
.B1(n_14),
.B2(n_27),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_83),
.B(n_95),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_89),
.B(n_78),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_72),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_101),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_65),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_104),
.B(n_45),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_106),
.B1(n_87),
.B2(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

AO221x1_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_94),
.B1(n_88),
.B2(n_82),
.C(n_81),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_112),
.C(n_114),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_63),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_113),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_75),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_97),
.C(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_119),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_103),
.C(n_102),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_104),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_121),
.B(n_125),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_108),
.C(n_113),
.Y(n_122)
);

OAI321xp33_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_112),
.A3(n_123),
.B1(n_121),
.B2(n_124),
.C(n_27),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_99),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_73),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_26),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_130),
.B(n_7),
.C(n_11),
.D(n_127),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_19),
.C(n_45),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_45),
.Y(n_132)
);


endmodule