module fake_jpeg_24184_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_6),
.B(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_7),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_40),
.B(n_25),
.C(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_6),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_22),
.B1(n_37),
.B2(n_38),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_36),
.B1(n_43),
.B2(n_21),
.Y(n_85)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_60),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_62),
.B(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_64),
.Y(n_119)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_22),
.B1(n_24),
.B2(n_17),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_69),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_44),
.B1(n_36),
.B2(n_22),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_85),
.B1(n_90),
.B2(n_34),
.Y(n_106)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_24),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_24),
.B1(n_17),
.B2(n_20),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_72),
.Y(n_107)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_78),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_34),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_87),
.Y(n_97)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_81),
.Y(n_105)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_86),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_34),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_39),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_42),
.B1(n_34),
.B2(n_17),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_40),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_106),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_16),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_77),
.B(n_34),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_64),
.C(n_74),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_62),
.A2(n_32),
.B1(n_30),
.B2(n_20),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_30),
.B1(n_26),
.B2(n_32),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_16),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_117),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_16),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_79),
.Y(n_118)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_71),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_84),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_125),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_85),
.B1(n_88),
.B2(n_82),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_142),
.B1(n_102),
.B2(n_112),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_135),
.C(n_93),
.Y(n_165)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_136),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_63),
.C(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_140),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_42),
.B1(n_71),
.B2(n_91),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_147),
.B1(n_148),
.B2(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_117),
.B1(n_120),
.B2(n_113),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_78),
.B1(n_65),
.B2(n_69),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_150),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_101),
.A2(n_73),
.B1(n_83),
.B2(n_81),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_97),
.A2(n_83),
.B1(n_86),
.B2(n_80),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_16),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_119),
.Y(n_151)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_174),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_153),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_97),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_154),
.B(n_172),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_155),
.A2(n_158),
.B1(n_162),
.B2(n_26),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_96),
.Y(n_156)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_160),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_121),
.B(n_115),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_161),
.A2(n_163),
.B(n_29),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_99),
.B1(n_94),
.B2(n_109),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_109),
.B(n_94),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_177),
.B(n_26),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_32),
.C(n_30),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_29),
.A3(n_84),
.B1(n_100),
.B2(n_23),
.C1(n_118),
.C2(n_19),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_166),
.B(n_145),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_178),
.B1(n_17),
.B2(n_28),
.Y(n_214)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_168),
.B(n_176),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_102),
.Y(n_169)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_102),
.Y(n_170)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_111),
.Y(n_171)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_16),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_131),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_111),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_21),
.B(n_20),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_126),
.A2(n_112),
.B1(n_21),
.B2(n_111),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_23),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_180),
.B(n_124),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_139),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_181),
.B(n_184),
.Y(n_197)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_163),
.B(n_135),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_185),
.B(n_187),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_148),
.B(n_141),
.C(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_146),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_206),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_209),
.B1(n_214),
.B2(n_171),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_191),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_203),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_198),
.C(n_210),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_144),
.C(n_128),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_207),
.B1(n_208),
.B2(n_212),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_29),
.Y(n_201)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_161),
.A2(n_25),
.B(n_19),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_18),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_173),
.A2(n_25),
.B1(n_28),
.B2(n_33),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_155),
.A2(n_184),
.B1(n_162),
.B2(n_152),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_170),
.B(n_174),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_33),
.C(n_28),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_156),
.B(n_33),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_160),
.A2(n_33),
.B1(n_28),
.B2(n_18),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_196),
.B(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_151),
.Y(n_222)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_199),
.B(n_168),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_226),
.A2(n_210),
.B1(n_242),
.B2(n_202),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_178),
.B1(n_176),
.B2(n_175),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_232),
.B1(n_239),
.B2(n_214),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_172),
.C(n_154),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_237),
.C(n_238),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_186),
.A2(n_182),
.B1(n_183),
.B2(n_159),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_204),
.A2(n_180),
.B1(n_159),
.B2(n_177),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_233),
.A2(n_241),
.B1(n_199),
.B2(n_11),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_212),
.Y(n_254)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_18),
.C(n_1),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_0),
.C(n_1),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_193),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_209),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_240),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_204),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_185),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_245),
.B(n_236),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_194),
.B(n_213),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_217),
.B(n_234),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_249),
.A2(n_257),
.B1(n_232),
.B2(n_244),
.Y(n_266)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_206),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_236),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_213),
.C(n_202),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_255),
.C(n_256),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_218),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_203),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_211),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_222),
.A2(n_193),
.B1(n_215),
.B2(n_187),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_215),
.C(n_188),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_260),
.C(n_239),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_205),
.C(n_191),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_227),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_262),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_263),
.B(n_218),
.Y(n_274)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_242),
.B1(n_230),
.B2(n_225),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_268),
.A2(n_278),
.B1(n_3),
.B2(n_4),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_269),
.B(n_280),
.Y(n_290)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_270),
.B(n_272),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_11),
.B(n_14),
.Y(n_291)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_2),
.Y(n_295)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_281),
.C(n_8),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_228),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_253),
.B1(n_252),
.B2(n_251),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_279),
.A2(n_258),
.B1(n_245),
.B2(n_246),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_0),
.C(n_2),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_264),
.A2(n_261),
.B1(n_260),
.B2(n_255),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_296),
.B1(n_267),
.B2(n_275),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_265),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_243),
.B1(n_246),
.B2(n_4),
.Y(n_287)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_288),
.B(n_4),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_11),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_295),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_291),
.A2(n_281),
.B(n_5),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_269),
.C(n_8),
.Y(n_304)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_298),
.B(n_304),
.Y(n_315)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_301),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_307),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_273),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_293),
.A2(n_278),
.B(n_280),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_302),
.A2(n_305),
.B(n_287),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_291),
.Y(n_316)
);

OAI321xp33_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_4),
.A3(n_12),
.B1(n_13),
.B2(n_15),
.C(n_286),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_13),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_285),
.Y(n_309)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_282),
.C(n_292),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_313),
.B(n_304),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_301),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_284),
.B1(n_294),
.B2(n_288),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_306),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_323),
.B(n_310),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_320),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_307),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_322),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_323),
.Y(n_327)
);

OAI21x1_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_324),
.B(n_326),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_319),
.B(n_315),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_314),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_312),
.B1(n_290),
.B2(n_15),
.Y(n_332)
);


endmodule