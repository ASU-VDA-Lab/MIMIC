module fake_jpeg_8300_n_144 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_25),
.Y(n_44)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_26),
.B1(n_22),
.B2(n_23),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_52),
.B1(n_37),
.B2(n_35),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_18),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_1),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_27),
.Y(n_63)
);

CKINVDCx6p67_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_51),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_33),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_61),
.B1(n_65),
.B2(n_73),
.Y(n_90)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_59),
.Y(n_91)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_66),
.Y(n_80)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_1),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_64),
.B(n_76),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_35),
.B1(n_32),
.B2(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_76),
.Y(n_81)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_39),
.B1(n_29),
.B2(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_50),
.C(n_45),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_3),
.C(n_4),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_1),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_87),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_53),
.A3(n_14),
.B1(n_4),
.B2(n_5),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_2),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_86),
.Y(n_108)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_67),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_2),
.B(n_3),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_7),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_5),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_10),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_7),
.B(n_8),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_9),
.B(n_10),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_73),
.B1(n_62),
.B2(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_103),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_97),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_70),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_73),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_81),
.C(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_85),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_62),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_96),
.B(n_80),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_111),
.B(n_112),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_108),
.C(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_107),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_85),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_124),
.C(n_125),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_109),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_102),
.C(n_101),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_112),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_101),
.B(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_114),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_128),
.A2(n_95),
.B(n_103),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_111),
.C(n_101),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_99),
.B1(n_119),
.B2(n_106),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_131),
.A2(n_127),
.B1(n_129),
.B2(n_68),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_89),
.B1(n_84),
.B2(n_10),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_125),
.C(n_83),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_134),
.C(n_11),
.Y(n_137)
);

AOI31xp67_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_78),
.A3(n_95),
.B(n_88),
.Y(n_135)
);

AOI31xp67_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_11),
.A3(n_13),
.B(n_54),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_136),
.B(n_138),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_139),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_142),
.B(n_140),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_137),
.Y(n_144)
);


endmodule