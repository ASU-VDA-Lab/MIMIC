module fake_netlist_1_6247_n_30 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NOR2x1_ASAP7_75t_L g13 ( .A(n_4), .B(n_5), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
AOI22xp5_ASAP7_75t_L g17 ( .A1(n_9), .A2(n_8), .B1(n_12), .B2(n_3), .Y(n_17) );
BUFx3_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_16), .B(n_0), .Y(n_19) );
OAI222xp33_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_17), .B1(n_13), .B2(n_4), .C1(n_5), .C2(n_6), .Y(n_20) );
OAI21x1_ASAP7_75t_L g21 ( .A1(n_18), .A2(n_10), .B(n_11), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
AOI211xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_20), .B(n_18), .C(n_21), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_24), .B(n_21), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_15), .Y(n_26) );
NAND4xp25_ASAP7_75t_SL g27 ( .A(n_25), .B(n_20), .C(n_2), .D(n_7), .Y(n_27) );
AOI21xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_21), .B(n_15), .Y(n_28) );
OAI22x1_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_27), .B1(n_2), .B2(n_7), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_1), .B1(n_8), .B2(n_27), .Y(n_30) );
endmodule