module real_jpeg_4544_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_1),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_1),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_1),
.A2(n_187),
.B1(n_243),
.B2(n_246),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_1),
.A2(n_187),
.B1(n_311),
.B2(n_313),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_1),
.A2(n_187),
.B1(n_322),
.B2(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_3),
.A2(n_137),
.B1(n_138),
.B2(n_140),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_3),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_140),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_3),
.A2(n_140),
.B1(n_198),
.B2(n_201),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_3),
.A2(n_140),
.B1(n_277),
.B2(n_358),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_4),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_4),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_4),
.A2(n_96),
.B1(n_132),
.B2(n_231),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_4),
.A2(n_96),
.B1(n_252),
.B2(n_256),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_4),
.A2(n_96),
.B1(n_209),
.B2(n_321),
.Y(n_320)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_5),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_5),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_5),
.Y(n_360)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_6),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_7),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_7),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_7),
.A2(n_266),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_7),
.A2(n_147),
.B1(n_266),
.B2(n_349),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_7),
.A2(n_80),
.B1(n_266),
.B2(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_8),
.A2(n_35),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_9),
.Y(n_93)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_9),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_10),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_10),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_10),
.A2(n_79),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_10),
.A2(n_79),
.B1(n_244),
.B2(n_285),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_10),
.A2(n_47),
.B1(n_79),
.B2(n_406),
.Y(n_405)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_12),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_12),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_12),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_12),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_12),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_12),
.Y(n_201)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_12),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_13),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_13),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_13),
.B(n_58),
.C(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_13),
.B(n_128),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_13),
.B(n_27),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_13),
.B(n_73),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_13),
.B(n_210),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_14),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_14),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_14),
.A2(n_69),
.B1(n_161),
.B2(n_165),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_14),
.A2(n_69),
.B1(n_147),
.B2(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_16),
.A2(n_42),
.B1(n_43),
.B2(n_47),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_16),
.A2(n_42),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_16),
.A2(n_39),
.B1(n_42),
.B2(n_64),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_215),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_213),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_190),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_20),
.B(n_190),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_111),
.C(n_157),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_21),
.A2(n_22),
.B1(n_111),
.B2(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_74),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_23),
.A2(n_24),
.B(n_76),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_24),
.A2(n_75),
.B1(n_76),
.B2(n_110),
.Y(n_74)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_24),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_24),
.A2(n_40),
.B1(n_110),
.B2(n_416),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_34),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_25),
.A2(n_34),
.B1(n_160),
.B2(n_168),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_25),
.A2(n_242),
.B(n_249),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_25),
.A2(n_228),
.B(n_249),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_25),
.A2(n_383),
.B1(n_384),
.B2(n_386),
.Y(n_382)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_26),
.B(n_251),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_26),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_26),
.A2(n_328),
.B1(n_357),
.B2(n_359),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_26),
.A2(n_387),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_31),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_31),
.Y(n_255)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_32),
.Y(n_250)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_37),
.Y(n_239)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_37),
.Y(n_259)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_40),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_68),
.B2(n_73),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_41),
.A2(n_49),
.B1(n_73),
.B2(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_43),
.Y(n_225)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_44),
.Y(n_173)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_45),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_45),
.Y(n_269)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_45),
.Y(n_407)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_46),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_46),
.Y(n_155)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_46),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_46),
.Y(n_233)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_49),
.A2(n_68),
.B1(n_73),
.B2(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_49),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_49),
.B(n_230),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_60),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_54),
.B1(n_57),
.B2(n_59),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_53),
.Y(n_313)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22x1_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_61),
.B1(n_64),
.B2(n_67),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_60),
.A2(n_152),
.B(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_60),
.A2(n_263),
.B(n_270),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_60),
.A2(n_204),
.B1(n_263),
.B2(n_310),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_60),
.A2(n_270),
.B(n_405),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_60),
.A2(n_204),
.B1(n_405),
.B2(n_420),
.Y(n_419)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_66),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g245 ( 
.A(n_66),
.Y(n_245)
);

BUFx8_ASAP7_75t_L g279 ( 
.A(n_66),
.Y(n_279)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_73),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_94),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_78),
.Y(n_195)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_80),
.B(n_228),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_82),
.B(n_95),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_82),
.Y(n_196)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_91),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_86),
.Y(n_372)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_87),
.Y(n_351)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_88),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_88),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_90),
.Y(n_379)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_94),
.A2(n_196),
.B(n_426),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_98),
.A2(n_105),
.B1(n_107),
.B2(n_109),
.Y(n_104)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_103),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_103),
.A2(n_394),
.B(n_397),
.Y(n_393)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_106),
.Y(n_373)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_111),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_149),
.B(n_156),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_150),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_128),
.B1(n_135),
.B2(n_141),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_114),
.A2(n_316),
.B(n_319),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_114),
.B(n_353),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_114),
.A2(n_128),
.B1(n_353),
.B2(n_431),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_114),
.A2(n_319),
.B(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_115),
.A2(n_136),
.B1(n_175),
.B2(n_181),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_115),
.A2(n_181),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_115),
.A2(n_181),
.B1(n_348),
.B2(n_400),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_128),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_121),
.B1(n_123),
.B2(n_126),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_119),
.Y(n_332)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_122),
.Y(n_403)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_125),
.Y(n_337)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_128),
.Y(n_181)
);

AO22x2_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_128)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_130),
.Y(n_236)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_130),
.Y(n_265)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_131),
.Y(n_312)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_139),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_SL g316 ( 
.A1(n_142),
.A2(n_228),
.B(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_156),
.B(n_191),
.CI(n_192),
.CON(n_190),
.SN(n_190)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_157),
.B(n_433),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_174),
.C(n_182),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_158),
.B(n_414),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_170),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_159),
.B(n_170),
.Y(n_441)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_160),
.Y(n_422)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_164),
.Y(n_248)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_165),
.Y(n_285)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_168),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_168),
.A2(n_291),
.B(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_168),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_169),
.Y(n_385)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_171),
.Y(n_420)
);

NAND2xp33_ASAP7_75t_SL g333 ( 
.A(n_172),
.B(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_174),
.B(n_182),
.Y(n_414)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_175),
.Y(n_431)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_181),
.B(n_320),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_181),
.A2(n_348),
.B(n_352),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B(n_189),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_183),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_183),
.A2(n_184),
.B1(n_196),
.B2(n_426),
.Y(n_425)
);

OAI32xp33_ASAP7_75t_L g369 ( 
.A1(n_185),
.A2(n_370),
.A3(n_373),
.B1(n_374),
.B2(n_380),
.Y(n_369)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx8_ASAP7_75t_L g429 ( 
.A(n_188),
.Y(n_429)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_189),
.Y(n_397)
);

BUFx24_ASAP7_75t_SL g474 ( 
.A(n_190),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_202),
.B2(n_212),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_196),
.B(n_228),
.Y(n_355)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_205),
.B1(n_206),
.B2(n_211),
.Y(n_202)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_204),
.A2(n_224),
.B(n_229),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_204),
.A2(n_229),
.B(n_310),
.Y(n_344)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI311xp33_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_410),
.A3(n_450),
.B1(n_468),
.C1(n_473),
.Y(n_216)
);

AOI21x1_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_363),
.B(n_409),
.Y(n_217)
);

AO21x1_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_339),
.B(n_362),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_304),
.B(n_338),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_273),
.B(n_303),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_240),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_222),
.B(n_240),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_234),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_223),
.A2(n_234),
.B1(n_235),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_223),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_SL g394 ( 
.A1(n_228),
.A2(n_380),
.B(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_260),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_241),
.B(n_261),
.C(n_272),
.Y(n_305)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_242),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_253),
.Y(n_358)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_271),
.B2(n_272),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_294),
.B(n_302),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_282),
.B(n_293),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_292),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_292),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_288),
.B(n_291),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_300),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_300),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_306),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_325),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_314),
.B2(n_315),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_314),
.C(n_325),
.Y(n_340)
);

AOI32xp33_ASAP7_75t_L g329 ( 
.A1(n_311),
.A2(n_318),
.A3(n_322),
.B1(n_330),
.B2(n_333),
.Y(n_329)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_320),
.Y(n_353)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_329),
.Y(n_345)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx8_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_340),
.B(n_341),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_346),
.B2(n_361),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_345),
.C(n_361),
.Y(n_364)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_346),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_354),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_355),
.C(n_356),
.Y(n_388)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_364),
.B(n_365),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_391),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_388),
.B1(n_389),
.B2(n_390),
.Y(n_366)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_367),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_381),
.B2(n_382),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_369),
.B(n_381),
.Y(n_445)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx12f_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_388),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_388),
.B(n_389),
.C(n_391),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_393),
.B1(n_398),
.B2(n_408),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_392),
.B(n_399),
.C(n_404),
.Y(n_459)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_398),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_404),
.Y(n_398)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx8_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

NAND2xp33_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_435),
.Y(n_410)
);

A2O1A1Ixp33_ASAP7_75t_SL g468 ( 
.A1(n_411),
.A2(n_435),
.B(n_469),
.C(n_472),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_432),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_412),
.B(n_432),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_415),
.C(n_417),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_415),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_449),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_424),
.C(n_430),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_419),
.B(n_421),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_421),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_424),
.A2(n_425),
.B1(n_430),
.B2(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_430),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_448),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_448),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_441),
.C(n_442),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_437),
.A2(n_438),
.B1(n_441),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_441),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_461),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_445),
.C(n_446),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_443),
.A2(n_444),
.B1(n_446),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_446),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_463),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_452),
.A2(n_470),
.B(n_471),
.Y(n_469)
);

NOR2x1_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_460),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_460),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_457),
.C(n_459),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_466),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_457),
.A2(n_458),
.B1(n_459),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_459),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_464),
.B(n_465),
.Y(n_470)
);


endmodule