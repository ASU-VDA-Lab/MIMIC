module fake_jpeg_20576_n_304 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_43),
.Y(n_51)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_59),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_19),
.B1(n_33),
.B2(n_24),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_62),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_44),
.B1(n_37),
.B2(n_20),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_20),
.B1(n_35),
.B2(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_19),
.B1(n_33),
.B2(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_22),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_69),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_86),
.Y(n_121)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_18),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_73),
.B(n_25),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_47),
.Y(n_74)
);

CKINVDCx10_ASAP7_75t_R g132 ( 
.A(n_74),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_40),
.C(n_26),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_32),
.C(n_30),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_22),
.B1(n_33),
.B2(n_24),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_54),
.B(n_48),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_78),
.A2(n_85),
.B(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_89),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_45),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_22),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_18),
.B(n_23),
.C(n_35),
.Y(n_89)
);

AO22x2_ASAP7_75t_SL g91 ( 
.A1(n_66),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_91)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_99),
.B1(n_32),
.B2(n_30),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_46),
.B(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_27),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_26),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_98),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_20),
.B1(n_36),
.B2(n_31),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_107),
.B1(n_108),
.B2(n_0),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_26),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_67),
.A2(n_42),
.B1(n_17),
.B2(n_35),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_58),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_101),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_61),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_39),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_67),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_50),
.A2(n_36),
.B1(n_31),
.B2(n_23),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_50),
.A2(n_29),
.B1(n_36),
.B2(n_31),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_51),
.B(n_29),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_27),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_32),
.B1(n_30),
.B2(n_27),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_110),
.A2(n_92),
.B1(n_87),
.B2(n_71),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_120),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_119),
.C(n_127),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_32),
.C(n_30),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_123),
.B(n_101),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_73),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_126),
.A2(n_138),
.B1(n_88),
.B2(n_82),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_25),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_72),
.B(n_27),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_130),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_25),
.C(n_21),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_136),
.C(n_91),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_84),
.B(n_25),
.C(n_21),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_70),
.B(n_15),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_13),
.Y(n_142)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_104),
.B(n_109),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_141),
.A2(n_143),
.B(n_149),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_146),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_86),
.B(n_79),
.Y(n_143)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_94),
.B1(n_79),
.B2(n_80),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_157),
.B1(n_161),
.B2(n_170),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_94),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_163),
.B(n_130),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_89),
.B(n_85),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_108),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_151),
.B(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_74),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_71),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_162),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_128),
.B1(n_139),
.B2(n_118),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_85),
.C(n_103),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_168),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_136),
.B1(n_115),
.B2(n_134),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_115),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g189 ( 
.A(n_160),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_120),
.A2(n_88),
.B1(n_91),
.B2(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_102),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_166),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_113),
.A2(n_91),
.B1(n_82),
.B2(n_106),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_132),
.B(n_125),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_171),
.A2(n_181),
.B(n_196),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_110),
.B1(n_138),
.B2(n_123),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_188),
.B1(n_199),
.B2(n_159),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_193),
.B1(n_195),
.B2(n_145),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_112),
.B(n_138),
.Y(n_181)
);

AO21x1_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_0),
.B(n_1),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_148),
.A2(n_133),
.B(n_116),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_10),
.B(n_9),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_134),
.B1(n_115),
.B2(n_106),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_83),
.C(n_124),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_163),
.C(n_150),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_124),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_168),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_140),
.A2(n_90),
.B1(n_105),
.B2(n_83),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_140),
.A2(n_90),
.B1(n_83),
.B2(n_13),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_148),
.B(n_143),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_144),
.B1(n_152),
.B2(n_146),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_160),
.B1(n_169),
.B2(n_164),
.Y(n_200)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_150),
.A2(n_83),
.B1(n_12),
.B2(n_10),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_205),
.B1(n_216),
.B2(n_219),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_203),
.C(n_215),
.Y(n_226)
);

BUFx12_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_211),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_174),
.B(n_156),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_204),
.B(n_206),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_183),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_142),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_141),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_208),
.B(n_213),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_155),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_165),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_214),
.B1(n_191),
.B2(n_1),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_183),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_151),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_158),
.C(n_145),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_175),
.A2(n_158),
.B1(n_162),
.B2(n_2),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_175),
.A2(n_196),
.B1(n_181),
.B2(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_222),
.C(n_189),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_0),
.C(n_1),
.Y(n_222)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

NAND5xp2_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_186),
.C(n_182),
.D(n_171),
.E(n_184),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_202),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_210),
.A2(n_178),
.B1(n_173),
.B2(n_194),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_231),
.B1(n_239),
.B2(n_240),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_172),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_230),
.B(n_213),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_198),
.B1(n_185),
.B2(n_189),
.Y(n_231)
);

NOR3xp33_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_199),
.C(n_189),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_232),
.B(n_237),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_191),
.B1(n_187),
.B2(n_2),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_0),
.C(n_1),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_203),
.C(n_208),
.Y(n_253)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_253),
.Y(n_262)
);

BUFx12f_ASAP7_75t_SL g246 ( 
.A(n_232),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_246),
.A2(n_261),
.B(n_228),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_255),
.Y(n_274)
);

OA22x2_ASAP7_75t_L g250 ( 
.A1(n_236),
.A2(n_211),
.B1(n_206),
.B2(n_212),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_250),
.A2(n_252),
.B1(n_239),
.B2(n_231),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_227),
.A2(n_216),
.B1(n_214),
.B2(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_233),
.C(n_215),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_257),
.B(n_260),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_221),
.C(n_209),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_258),
.B(n_259),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_226),
.B(n_223),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_229),
.B(n_220),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_234),
.A2(n_223),
.B(n_218),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_234),
.B1(n_228),
.B2(n_235),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_263),
.A2(n_251),
.B1(n_250),
.B2(n_253),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_236),
.B(n_244),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_267),
.B(n_261),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_271),
.B1(n_254),
.B2(n_250),
.Y(n_280)
);

FAx1_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_235),
.CI(n_202),
.CON(n_268),
.SN(n_268)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_273),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_251),
.A2(n_242),
.B1(n_225),
.B2(n_218),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_241),
.B(n_217),
.Y(n_272)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_249),
.B(n_2),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_278),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_265),
.B1(n_271),
.B2(n_269),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_263),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_250),
.B(n_258),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_280),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_257),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_3),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_3),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_3),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_268),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_289),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_275),
.A2(n_262),
.B(n_268),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_286),
.B(n_277),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_294),
.B(n_295),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_279),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_291),
.B(n_280),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_285),
.A3(n_276),
.B1(n_287),
.B2(n_7),
.C1(n_4),
.C2(n_6),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g298 ( 
.A(n_293),
.B(n_278),
.CI(n_288),
.CON(n_298),
.SN(n_298)
);

AOI322xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_299),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_297),
.A2(n_292),
.B(n_298),
.Y(n_300)
);

AOI321xp33_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_301),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_5),
.Y(n_304)
);


endmodule