module fake_jpeg_8691_n_174 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx11_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_12),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_34),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_27),
.B1(n_18),
.B2(n_19),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_19),
.B1(n_18),
.B2(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_44),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_34),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_13),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_35),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_29),
.B(n_25),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_58),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_28),
.B1(n_34),
.B2(n_17),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_25),
.B1(n_17),
.B2(n_24),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_35),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_28),
.B1(n_26),
.B2(n_23),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_68),
.B1(n_48),
.B2(n_54),
.Y(n_84)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_49),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_28),
.B1(n_33),
.B2(n_29),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_80),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_88),
.B(n_50),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_22),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_67),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_42),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_58),
.C(n_66),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_85),
.B1(n_21),
.B2(n_73),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_24),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_60),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_59),
.B(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_101),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_69),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_95),
.B1(n_75),
.B2(n_70),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_94),
.B(n_106),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_106),
.C(n_90),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_44),
.B1(n_65),
.B2(n_42),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_64),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_104),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_42),
.B1(n_21),
.B2(n_68),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_68),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_83),
.B(n_88),
.Y(n_108)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_107),
.B(n_78),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_102),
.B1(n_94),
.B2(n_97),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_116),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_72),
.C(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_102),
.C(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_120),
.B(n_122),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_130),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_118),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_133),
.Y(n_146)
);

XOR2x2_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_96),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_136),
.B1(n_121),
.B2(n_49),
.Y(n_144)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_134),
.A2(n_135),
.B1(n_121),
.B2(n_22),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_93),
.B1(n_71),
.B2(n_70),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_138),
.B(n_142),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_112),
.C(n_113),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_140),
.C(n_141),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_110),
.C(n_111),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_114),
.C(n_52),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_136),
.B(n_131),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_145),
.B(n_99),
.Y(n_150)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_126),
.C(n_129),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_137),
.C(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_154),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_140),
.B(n_142),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_156),
.C(n_157),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_99),
.B(n_10),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_153),
.C(n_152),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_163),
.B(n_164),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_160),
.B(n_9),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_158),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_158),
.B(n_63),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_166),
.A2(n_161),
.B1(n_2),
.B2(n_3),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.C(n_1),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_161),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_171),
.A3(n_1),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_172)
);

OAI221xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.C(n_14),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_169),
.Y(n_174)
);


endmodule