module real_jpeg_8314_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

AOI21xp33_ASAP7_75t_L g28 ( 
.A1(n_3),
.A2(n_27),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_3),
.B(n_64),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_25),
.B1(n_30),
.B2(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_3),
.A2(n_55),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_3),
.B(n_55),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_3),
.A2(n_38),
.B1(n_43),
.B2(n_143),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_7),
.A2(n_55),
.B(n_79),
.C(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_7),
.B(n_55),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

BUFx6f_ASAP7_75t_SL g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_10),
.A2(n_53),
.B1(n_55),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_10),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_83),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_11),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_11),
.A2(n_53),
.B1(n_55),
.B2(n_70),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_13),
.A2(n_29),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_13),
.A2(n_30),
.B1(n_58),
.B2(n_95),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_13),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_58),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_14),
.A2(n_29),
.B1(n_59),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_61),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_14),
.A2(n_53),
.B1(n_55),
.B2(n_61),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_15),
.A2(n_29),
.B1(n_59),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_15),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_15),
.A2(n_53),
.B1(n_55),
.B2(n_89),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_89),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_118),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_117),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_98),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_20),
.B(n_98),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_44),
.B1(n_71),
.B2(n_72),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.C(n_30),
.Y(n_24)
);

HAxp5_ASAP7_75t_SL g111 ( 
.A(n_25),
.B(n_29),
.CON(n_111),
.SN(n_111)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_25),
.B(n_80),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_25),
.B(n_43),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_25),
.B(n_62),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_59),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_26),
.A2(n_30),
.B(n_65),
.C(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_26),
.B(n_30),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_49),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_30),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_33),
.A2(n_43),
.B(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_34),
.B(n_81),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_34),
.B(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_35),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_38),
.A2(n_114),
.B(n_116),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_38),
.A2(n_43),
.B1(n_125),
.B2(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_38),
.A2(n_127),
.B(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_39),
.B(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_39),
.A2(n_40),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_40),
.B(n_69),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_40),
.B(n_115),
.Y(n_158)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_63),
.C(n_66),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_45),
.A2(n_46),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_56),
.B1(n_60),
.B2(n_62),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_60),
.B1(n_62),
.B2(n_88),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_48),
.A2(n_52),
.B1(n_57),
.B2(n_111),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_50),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_49),
.B(n_55),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_51),
.A2(n_53),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_63),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_64),
.A2(n_91),
.B1(n_94),
.B2(n_96),
.Y(n_90)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_90),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_86),
.B2(n_87),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_82),
.B(n_84),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_78),
.A2(n_80),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_78),
.A2(n_80),
.B1(n_133),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_78),
.A2(n_80),
.B1(n_105),
.B2(n_156),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.C(n_108),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_99),
.A2(n_100),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_104),
.A2(n_108),
.B1(n_109),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_104),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_110),
.B(n_113),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_171),
.B(n_177),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_160),
.B(n_170),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_150),
.B(n_159),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_139),
.B(n_149),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_128),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_128),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_134),
.B2(n_138),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_138),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_132),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_144),
.B(n_148),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_141),
.B(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_151),
.B(n_152),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_153),
.B(n_161),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_155),
.CI(n_157),
.CON(n_153),
.SN(n_153)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_169),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_164),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_165),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_167),
.C(n_169),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_168),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_172),
.B(n_173),
.Y(n_177)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);


endmodule