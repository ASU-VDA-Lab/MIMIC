module fake_jpeg_3516_n_137 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_0),
.B(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_28),
.B(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_6),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_11),
.B(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_46),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_2),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_45),
.Y(n_56)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_7),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_22),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_25),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_23),
.C(n_27),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_17),
.C(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_9),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_51),
.B(n_68),
.Y(n_91)
);

NAND2x1_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_69),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_22),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_70),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_28),
.A2(n_27),
.B1(n_16),
.B2(n_12),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_67),
.B1(n_56),
.B2(n_74),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_36),
.A2(n_16),
.B1(n_12),
.B2(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_25),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_35),
.A2(n_38),
.B(n_48),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NAND2xp67_ASAP7_75t_SL g72 ( 
.A(n_37),
.B(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_43),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_65),
.A2(n_40),
.B1(n_33),
.B2(n_44),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_89),
.B1(n_93),
.B2(n_55),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_56),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_92),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_52),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_64),
.B1(n_52),
.B2(n_67),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_66),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_75),
.B1(n_55),
.B2(n_54),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_89),
.B1(n_94),
.B2(n_92),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_53),
.B(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_77),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_103),
.B1(n_92),
.B2(n_99),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_66),
.B1(n_79),
.B2(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_93),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_114),
.B1(n_102),
.B2(n_107),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_76),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_105),
.B(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_113),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_84),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_115),
.Y(n_117)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_99),
.C(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_103),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_111),
.B(n_109),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_120),
.B(n_121),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_122),
.B(n_123),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_117),
.B(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_118),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_95),
.C(n_98),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_98),
.C(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_128),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_124),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_132),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.C(n_130),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_127),
.Y(n_137)
);


endmodule