module real_aes_7204_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g107 ( .A(n_0), .Y(n_107) );
INVx1_ASAP7_75t_L g533 ( .A(n_1), .Y(n_533) );
INVx1_ASAP7_75t_L g154 ( .A(n_2), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_3), .A2(n_38), .B1(n_179), .B2(n_479), .Y(n_502) );
AOI21xp33_ASAP7_75t_L g186 ( .A1(n_4), .A2(n_170), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_5), .B(n_168), .Y(n_545) );
AND2x6_ASAP7_75t_L g147 ( .A(n_6), .B(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_7), .A2(n_257), .B(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_8), .B(n_113), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_8), .B(n_39), .Y(n_121) );
INVx1_ASAP7_75t_L g192 ( .A(n_9), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_10), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g139 ( .A(n_11), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_12), .B(n_160), .Y(n_488) );
INVx1_ASAP7_75t_L g263 ( .A(n_13), .Y(n_263) );
INVx1_ASAP7_75t_L g527 ( .A(n_14), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_15), .B(n_135), .Y(n_516) );
AO32x2_ASAP7_75t_L g500 ( .A1(n_16), .A2(n_134), .A3(n_168), .B1(n_481), .B2(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_17), .B(n_179), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_18), .B(n_175), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_19), .B(n_135), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_20), .A2(n_49), .B1(n_179), .B2(n_479), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_21), .B(n_170), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_22), .A2(n_98), .B1(n_735), .B2(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_22), .Y(n_736) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_23), .A2(n_76), .B1(n_160), .B2(n_179), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_24), .B(n_179), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_25), .B(n_182), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_26), .A2(n_261), .B(n_262), .C(n_264), .Y(n_260) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_27), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_28), .B(n_165), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_29), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_30), .B(n_116), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_31), .A2(n_88), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_31), .Y(n_125) );
INVx1_ASAP7_75t_L g207 ( .A(n_32), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_33), .B(n_165), .Y(n_472) );
INVx2_ASAP7_75t_L g145 ( .A(n_34), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_35), .B(n_179), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_36), .B(n_165), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_37), .A2(n_147), .B(n_150), .C(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g113 ( .A(n_39), .Y(n_113) );
INVx1_ASAP7_75t_L g205 ( .A(n_40), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_41), .B(n_158), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_42), .B(n_179), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_43), .A2(n_86), .B1(n_227), .B2(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_44), .B(n_179), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_45), .B(n_179), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g208 ( .A(n_46), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_47), .B(n_532), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_48), .B(n_170), .Y(n_251) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_50), .A2(n_60), .B1(n_160), .B2(n_179), .Y(n_520) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_51), .A2(n_733), .B1(n_734), .B2(n_737), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_51), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_52), .A2(n_150), .B1(n_160), .B2(n_203), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_53), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_54), .B(n_179), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g141 ( .A(n_55), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_56), .B(n_179), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_57), .A2(n_178), .B(n_190), .C(n_191), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_58), .Y(n_240) );
INVx1_ASAP7_75t_L g188 ( .A(n_59), .Y(n_188) );
INVx1_ASAP7_75t_L g148 ( .A(n_61), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_62), .B(n_179), .Y(n_534) );
INVx1_ASAP7_75t_L g138 ( .A(n_63), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_64), .Y(n_444) );
AO32x2_ASAP7_75t_L g476 ( .A1(n_65), .A2(n_168), .A3(n_243), .B1(n_477), .B2(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g552 ( .A(n_66), .Y(n_552) );
INVx1_ASAP7_75t_L g467 ( .A(n_67), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_68), .A2(n_123), .B1(n_439), .B2(n_440), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_68), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_SL g174 ( .A1(n_69), .A2(n_175), .B(n_176), .C(n_178), .Y(n_174) );
INVxp67_ASAP7_75t_L g177 ( .A(n_70), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_71), .B(n_160), .Y(n_468) );
INVx1_ASAP7_75t_L g111 ( .A(n_72), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_73), .Y(n_210) );
INVx1_ASAP7_75t_L g233 ( .A(n_74), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_75), .A2(n_104), .B1(n_114), .B2(n_743), .Y(n_103) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_77), .A2(n_147), .B(n_150), .C(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_78), .B(n_479), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_79), .B(n_160), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_80), .B(n_155), .Y(n_223) );
INVx2_ASAP7_75t_L g136 ( .A(n_81), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_82), .B(n_175), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_83), .B(n_160), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g149 ( .A1(n_84), .A2(n_147), .B(n_150), .C(n_153), .Y(n_149) );
INVx2_ASAP7_75t_L g108 ( .A(n_85), .Y(n_108) );
OR2x2_ASAP7_75t_L g118 ( .A(n_85), .B(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g450 ( .A(n_85), .B(n_120), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_87), .A2(n_102), .B1(n_160), .B2(n_161), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_88), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_89), .B(n_165), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_90), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_91), .A2(n_147), .B(n_150), .C(n_246), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_92), .Y(n_253) );
INVx1_ASAP7_75t_L g173 ( .A(n_93), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_94), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_95), .B(n_155), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_96), .B(n_160), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_97), .B(n_168), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_98), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_99), .B(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_100), .A2(n_170), .B(n_171), .Y(n_169) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_101), .A2(n_447), .B1(n_731), .B2(n_732), .C1(n_738), .C2(n_741), .Y(n_446) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g744 ( .A(n_105), .Y(n_744) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_112), .Y(n_105) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_108), .C(n_109), .Y(n_106) );
AND2x2_ASAP7_75t_L g120 ( .A(n_107), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g454 ( .A(n_108), .B(n_120), .Y(n_454) );
NOR2x2_ASAP7_75t_L g740 ( .A(n_108), .B(n_119), .Y(n_740) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AO21x1_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_442), .B(n_445), .Y(n_114) );
OAI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_122), .B(n_441), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g440 ( .A(n_123), .Y(n_440) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_127), .Y(n_123) );
INVx1_ASAP7_75t_L g451 ( .A(n_127), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g741 ( .A1(n_127), .A2(n_452), .B1(n_456), .B2(n_742), .Y(n_741) );
NAND2x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_355), .Y(n_127) );
NOR5xp2_ASAP7_75t_L g128 ( .A(n_129), .B(n_278), .C(n_310), .D(n_325), .E(n_342), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_194), .B(n_215), .C(n_266), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_166), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_131), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_131), .B(n_330), .Y(n_393) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_132), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_132), .B(n_212), .Y(n_279) );
AND2x2_ASAP7_75t_L g320 ( .A(n_132), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_132), .B(n_289), .Y(n_324) );
OR2x2_ASAP7_75t_L g361 ( .A(n_132), .B(n_200), .Y(n_361) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g199 ( .A(n_133), .B(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g269 ( .A(n_133), .Y(n_269) );
OR2x2_ASAP7_75t_L g432 ( .A(n_133), .B(n_272), .Y(n_432) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_140), .B(n_162), .Y(n_133) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_134), .A2(n_201), .B(n_209), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_134), .B(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g228 ( .A(n_134), .Y(n_228) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_136), .B(n_137), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
OAI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_149), .Y(n_140) );
OAI22xp33_ASAP7_75t_L g201 ( .A1(n_142), .A2(n_180), .B1(n_202), .B2(n_208), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_142), .A2(n_233), .B(n_234), .Y(n_232) );
NAND2x1p5_ASAP7_75t_L g142 ( .A(n_143), .B(n_147), .Y(n_142) );
AND2x4_ASAP7_75t_L g170 ( .A(n_143), .B(n_147), .Y(n_170) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx1_ASAP7_75t_L g532 ( .A(n_144), .Y(n_532) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
INVx1_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
INVx1_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
INVx3_ASAP7_75t_L g156 ( .A(n_146), .Y(n_156) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_146), .Y(n_158) );
INVx1_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_146), .Y(n_204) );
INVx4_ASAP7_75t_SL g180 ( .A(n_147), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_147), .A2(n_466), .B(n_469), .Y(n_465) );
BUFx3_ASAP7_75t_L g481 ( .A(n_147), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_147), .A2(n_486), .B(n_490), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_147), .A2(n_526), .B(n_530), .Y(n_525) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_147), .A2(n_539), .B(n_542), .Y(n_538) );
INVx5_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
AND2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
BUFx3_ASAP7_75t_L g227 ( .A(n_151), .Y(n_227) );
INVx1_ASAP7_75t_L g479 ( .A(n_151), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_157), .C(n_159), .Y(n_153) );
O2A1O1Ixp5_ASAP7_75t_SL g466 ( .A1(n_155), .A2(n_178), .B(n_467), .C(n_468), .Y(n_466) );
INVx2_ASAP7_75t_L g503 ( .A(n_155), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_155), .A2(n_540), .B(n_541), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_155), .A2(n_549), .B(n_550), .Y(n_548) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_156), .B(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_156), .B(n_192), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g477 ( .A1(n_156), .A2(n_158), .B1(n_478), .B2(n_480), .Y(n_477) );
INVx2_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
INVx4_ASAP7_75t_L g249 ( .A(n_158), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_158), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_158), .A2(n_503), .B1(n_519), .B2(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_159), .A2(n_527), .B(n_528), .C(n_529), .Y(n_526) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_164), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_164), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g243 ( .A(n_165), .Y(n_243) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_165), .A2(n_256), .B(n_265), .Y(n_255) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_165), .A2(n_465), .B(n_472), .Y(n_464) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_165), .A2(n_485), .B(n_493), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_166), .A2(n_335), .B1(n_336), .B2(n_339), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_166), .B(n_269), .Y(n_418) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_184), .Y(n_166) );
AND2x2_ASAP7_75t_L g214 ( .A(n_167), .B(n_200), .Y(n_214) );
AND2x2_ASAP7_75t_L g271 ( .A(n_167), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g276 ( .A(n_167), .Y(n_276) );
INVx3_ASAP7_75t_L g289 ( .A(n_167), .Y(n_289) );
OR2x2_ASAP7_75t_L g309 ( .A(n_167), .B(n_272), .Y(n_309) );
AND2x2_ASAP7_75t_L g328 ( .A(n_167), .B(n_185), .Y(n_328) );
BUFx2_ASAP7_75t_L g360 ( .A(n_167), .Y(n_360) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_181), .Y(n_167) );
INVx4_ASAP7_75t_L g183 ( .A(n_168), .Y(n_183) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_168), .A2(n_538), .B(n_545), .Y(n_537) );
BUFx2_ASAP7_75t_L g257 ( .A(n_170), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_174), .C(n_180), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_172), .A2(n_180), .B(n_188), .C(n_189), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_172), .A2(n_180), .B(n_259), .C(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g489 ( .A(n_175), .Y(n_489) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_179), .Y(n_250) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_182), .A2(n_186), .B(n_193), .Y(n_185) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_SL g229 ( .A(n_183), .B(n_230), .Y(n_229) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_183), .B(n_481), .C(n_518), .Y(n_517) );
AO21x1_ASAP7_75t_L g607 ( .A1(n_183), .A2(n_518), .B(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g275 ( .A(n_184), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
BUFx2_ASAP7_75t_L g198 ( .A(n_185), .Y(n_198) );
INVx2_ASAP7_75t_L g213 ( .A(n_185), .Y(n_213) );
OR2x2_ASAP7_75t_L g291 ( .A(n_185), .B(n_272), .Y(n_291) );
AND2x2_ASAP7_75t_L g321 ( .A(n_185), .B(n_200), .Y(n_321) );
AND2x2_ASAP7_75t_L g338 ( .A(n_185), .B(n_269), .Y(n_338) );
AND2x2_ASAP7_75t_L g378 ( .A(n_185), .B(n_289), .Y(n_378) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_185), .B(n_214), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_190), .A2(n_491), .B(n_492), .Y(n_490) );
O2A1O1Ixp5_ASAP7_75t_L g551 ( .A1(n_190), .A2(n_531), .B(n_552), .C(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp33_ASAP7_75t_SL g195 ( .A(n_196), .B(n_211), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_199), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_197), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
OAI21xp33_ASAP7_75t_L g352 ( .A1(n_198), .A2(n_214), .B(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_198), .B(n_200), .Y(n_408) );
AND2x2_ASAP7_75t_L g344 ( .A(n_199), .B(n_345), .Y(n_344) );
INVx3_ASAP7_75t_L g272 ( .A(n_200), .Y(n_272) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_200), .Y(n_370) );
OAI22xp5_ASAP7_75t_SL g203 ( .A1(n_204), .A2(n_205), .B1(n_206), .B2(n_207), .Y(n_203) );
INVx2_ASAP7_75t_L g206 ( .A(n_204), .Y(n_206) );
INVx4_ASAP7_75t_L g261 ( .A(n_204), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_211), .B(n_269), .Y(n_437) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_212), .A2(n_380), .B1(n_381), .B2(n_386), .Y(n_379) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AND2x2_ASAP7_75t_L g270 ( .A(n_213), .B(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g308 ( .A(n_213), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_SL g345 ( .A(n_213), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_214), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g399 ( .A(n_214), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_241), .Y(n_216) );
INVx4_ASAP7_75t_L g285 ( .A(n_217), .Y(n_285) );
AND2x2_ASAP7_75t_L g363 ( .A(n_217), .B(n_330), .Y(n_363) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_231), .Y(n_217) );
INVx3_ASAP7_75t_L g282 ( .A(n_218), .Y(n_282) );
AND2x2_ASAP7_75t_L g296 ( .A(n_218), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g300 ( .A(n_218), .Y(n_300) );
INVx2_ASAP7_75t_L g314 ( .A(n_218), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_218), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g371 ( .A(n_218), .B(n_366), .Y(n_371) );
AND2x2_ASAP7_75t_L g436 ( .A(n_218), .B(n_406), .Y(n_436) );
OR2x6_ASAP7_75t_L g218 ( .A(n_219), .B(n_229), .Y(n_218) );
AOI21xp5_ASAP7_75t_SL g219 ( .A1(n_220), .A2(n_221), .B(n_228), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_225), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_225), .A2(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g264 ( .A(n_227), .Y(n_264) );
INVx1_ASAP7_75t_L g238 ( .A(n_228), .Y(n_238) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_228), .A2(n_525), .B(n_535), .Y(n_524) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_228), .A2(n_547), .B(n_554), .Y(n_546) );
AND2x2_ASAP7_75t_L g277 ( .A(n_231), .B(n_255), .Y(n_277) );
INVx2_ASAP7_75t_L g297 ( .A(n_231), .Y(n_297) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_238), .B(n_239), .Y(n_231) );
INVx1_ASAP7_75t_L g302 ( .A(n_241), .Y(n_302) );
AND2x2_ASAP7_75t_L g348 ( .A(n_241), .B(n_296), .Y(n_348) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_254), .Y(n_241) );
INVx2_ASAP7_75t_L g287 ( .A(n_242), .Y(n_287) );
INVx1_ASAP7_75t_L g295 ( .A(n_242), .Y(n_295) );
AND2x2_ASAP7_75t_L g313 ( .A(n_242), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_242), .B(n_297), .Y(n_351) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_252), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_251), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_250), .Y(n_246) );
AND2x2_ASAP7_75t_L g330 ( .A(n_254), .B(n_287), .Y(n_330) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g283 ( .A(n_255), .Y(n_283) );
AND2x2_ASAP7_75t_L g366 ( .A(n_255), .B(n_297), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_261), .B(n_263), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_261), .A2(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g529 ( .A(n_261), .Y(n_529) );
OAI21xp5_ASAP7_75t_SL g266 ( .A1(n_267), .A2(n_273), .B(n_277), .Y(n_266) );
INVx1_ASAP7_75t_SL g311 ( .A(n_267), .Y(n_311) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_268), .B(n_275), .Y(n_368) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g317 ( .A(n_269), .B(n_272), .Y(n_317) );
AND2x2_ASAP7_75t_L g346 ( .A(n_269), .B(n_290), .Y(n_346) );
OR2x2_ASAP7_75t_L g349 ( .A(n_269), .B(n_309), .Y(n_349) );
AOI222xp33_ASAP7_75t_L g413 ( .A1(n_270), .A2(n_362), .B1(n_414), .B2(n_415), .C1(n_417), .C2(n_419), .Y(n_413) );
BUFx2_ASAP7_75t_L g327 ( .A(n_272), .Y(n_327) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g316 ( .A(n_275), .B(n_317), .Y(n_316) );
INVx3_ASAP7_75t_SL g333 ( .A(n_275), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_275), .B(n_327), .Y(n_387) );
AND2x2_ASAP7_75t_L g322 ( .A(n_277), .B(n_282), .Y(n_322) );
INVx1_ASAP7_75t_L g341 ( .A(n_277), .Y(n_341) );
OAI221xp5_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_280), .B1(n_284), .B2(n_288), .C(n_292), .Y(n_278) );
OR2x2_ASAP7_75t_L g350 ( .A(n_280), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g335 ( .A(n_282), .B(n_305), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_282), .B(n_295), .Y(n_375) );
AND2x2_ASAP7_75t_L g380 ( .A(n_282), .B(n_330), .Y(n_380) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_282), .Y(n_390) );
NAND2x1_ASAP7_75t_SL g401 ( .A(n_282), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g286 ( .A(n_283), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_283), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_283), .B(n_301), .Y(n_332) );
INVx1_ASAP7_75t_L g398 ( .A(n_283), .Y(n_398) );
INVx1_ASAP7_75t_L g373 ( .A(n_284), .Y(n_373) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g385 ( .A(n_285), .Y(n_385) );
NOR2xp67_ASAP7_75t_L g397 ( .A(n_285), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g402 ( .A(n_286), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_286), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g305 ( .A(n_287), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_287), .B(n_297), .Y(n_318) );
INVx1_ASAP7_75t_L g384 ( .A(n_287), .Y(n_384) );
INVx1_ASAP7_75t_L g405 ( .A(n_288), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_298), .B(n_307), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
AND2x2_ASAP7_75t_L g438 ( .A(n_294), .B(n_371), .Y(n_438) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g406 ( .A(n_295), .B(n_366), .Y(n_406) );
AOI32xp33_ASAP7_75t_L g319 ( .A1(n_296), .A2(n_302), .A3(n_320), .B1(n_322), .B2(n_323), .Y(n_319) );
AOI322xp5_ASAP7_75t_L g421 ( .A1(n_296), .A2(n_328), .A3(n_411), .B1(n_422), .B2(n_423), .C1(n_424), .C2(n_426), .Y(n_421) );
INVx2_ASAP7_75t_L g301 ( .A(n_297), .Y(n_301) );
INVx1_ASAP7_75t_L g411 ( .A(n_297), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B1(n_303), .B2(n_304), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_299), .B(n_305), .Y(n_354) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_300), .B(n_366), .Y(n_416) );
INVx1_ASAP7_75t_L g303 ( .A(n_301), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_301), .B(n_330), .Y(n_420) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_309), .B(n_404), .Y(n_403) );
OAI221xp5_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_312), .B1(n_315), .B2(n_318), .C(n_319), .Y(n_310) );
OR2x2_ASAP7_75t_L g331 ( .A(n_312), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g340 ( .A(n_312), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g365 ( .A(n_313), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g369 ( .A(n_323), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI221xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B1(n_331), .B2(n_333), .C(n_334), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_327), .A2(n_358), .B1(n_362), .B2(n_363), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_328), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_328), .Y(n_433) );
INVx1_ASAP7_75t_L g427 ( .A(n_330), .Y(n_427) );
INVx1_ASAP7_75t_SL g362 ( .A(n_331), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_333), .B(n_361), .Y(n_423) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_338), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g404 ( .A(n_338), .Y(n_404) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
OAI221xp5_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_347), .B1(n_349), .B2(n_350), .C(n_352), .Y(n_342) );
NOR2xp33_ASAP7_75t_SL g343 ( .A(n_344), .B(n_346), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_344), .A2(n_362), .B1(n_408), .B2(n_409), .Y(n_407) );
CKINVDCx14_ASAP7_75t_R g347 ( .A(n_348), .Y(n_347) );
OAI21xp33_ASAP7_75t_L g426 ( .A1(n_349), .A2(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR3xp33_ASAP7_75t_SL g355 ( .A(n_356), .B(n_388), .C(n_412), .Y(n_355) );
NAND4xp25_ASAP7_75t_L g356 ( .A(n_357), .B(n_364), .C(n_372), .D(n_379), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g435 ( .A(n_360), .Y(n_435) );
INVx3_ASAP7_75t_SL g429 ( .A(n_361), .Y(n_429) );
OR2x2_ASAP7_75t_L g434 ( .A(n_361), .B(n_435), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B1(n_369), .B2(n_371), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_366), .B(n_384), .Y(n_425) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI21xp5_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_374), .B(n_376), .Y(n_372) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI211xp5_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_391), .B(n_394), .C(n_407), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g422 ( .A(n_393), .Y(n_422) );
AOI222xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_399), .B1(n_400), .B2(n_403), .C1(n_405), .C2(n_406), .Y(n_394) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND4xp25_ASAP7_75t_SL g431 ( .A(n_404), .B(n_432), .C(n_433), .D(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND3xp33_ASAP7_75t_SL g412 ( .A(n_413), .B(n_421), .C(n_430), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_436), .B1(n_437), .B2(n_438), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g445 ( .A1(n_441), .A2(n_442), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_451), .B1(n_452), .B2(n_455), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g742 ( .A(n_449), .Y(n_742) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_652), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_601), .C(n_643), .Y(n_457) );
AOI211xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_510), .B(n_555), .C(n_577), .Y(n_458) );
OAI211xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_473), .B(n_494), .C(n_505), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_461), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g664 ( .A(n_461), .B(n_581), .Y(n_664) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g566 ( .A(n_462), .B(n_497), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_462), .B(n_484), .Y(n_683) );
INVx1_ASAP7_75t_L g701 ( .A(n_462), .Y(n_701) );
AND2x2_ASAP7_75t_L g710 ( .A(n_462), .B(n_598), .Y(n_710) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g593 ( .A(n_463), .B(n_484), .Y(n_593) );
AND2x2_ASAP7_75t_L g651 ( .A(n_463), .B(n_598), .Y(n_651) );
INVx1_ASAP7_75t_L g695 ( .A(n_463), .Y(n_695) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g572 ( .A(n_464), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g580 ( .A(n_464), .Y(n_580) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_464), .Y(n_620) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_482), .Y(n_474) );
AND2x2_ASAP7_75t_L g559 ( .A(n_475), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g592 ( .A(n_475), .Y(n_592) );
OR2x2_ASAP7_75t_L g718 ( .A(n_475), .B(n_719), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_475), .B(n_484), .Y(n_722) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g497 ( .A(n_476), .Y(n_497) );
INVx1_ASAP7_75t_L g508 ( .A(n_476), .Y(n_508) );
AND2x2_ASAP7_75t_L g581 ( .A(n_476), .B(n_499), .Y(n_581) );
AND2x2_ASAP7_75t_L g621 ( .A(n_476), .B(n_500), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_481), .A2(n_548), .B(n_551), .Y(n_547) );
INVxp67_ASAP7_75t_L g663 ( .A(n_482), .Y(n_663) );
AND2x4_ASAP7_75t_L g688 ( .A(n_482), .B(n_581), .Y(n_688) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_SL g579 ( .A(n_483), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g498 ( .A(n_484), .B(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g567 ( .A(n_484), .B(n_500), .Y(n_567) );
INVx1_ASAP7_75t_L g573 ( .A(n_484), .Y(n_573) );
INVx2_ASAP7_75t_L g599 ( .A(n_484), .Y(n_599) );
AND2x2_ASAP7_75t_L g615 ( .A(n_484), .B(n_616), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_495), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g570 ( .A(n_497), .Y(n_570) );
AND2x2_ASAP7_75t_L g678 ( .A(n_497), .B(n_499), .Y(n_678) );
AND2x2_ASAP7_75t_L g595 ( .A(n_498), .B(n_580), .Y(n_595) );
AND2x2_ASAP7_75t_L g694 ( .A(n_498), .B(n_695), .Y(n_694) );
NOR2xp67_ASAP7_75t_L g616 ( .A(n_499), .B(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g719 ( .A(n_499), .B(n_580), .Y(n_719) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g509 ( .A(n_500), .Y(n_509) );
AND2x2_ASAP7_75t_L g598 ( .A(n_500), .B(n_599), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_503), .A2(n_531), .B(n_533), .C(n_534), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_503), .A2(n_543), .B(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
AND2x2_ASAP7_75t_L g644 ( .A(n_507), .B(n_579), .Y(n_644) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_508), .B(n_580), .Y(n_629) );
INVx2_ASAP7_75t_L g628 ( .A(n_509), .Y(n_628) );
OAI222xp33_ASAP7_75t_L g632 ( .A1(n_509), .A2(n_572), .B1(n_633), .B2(n_635), .C1(n_636), .C2(n_639), .Y(n_632) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_521), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g557 ( .A(n_514), .Y(n_557) );
OR2x2_ASAP7_75t_L g668 ( .A(n_514), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx3_ASAP7_75t_L g590 ( .A(n_515), .Y(n_590) );
NOR2x1_ASAP7_75t_L g641 ( .A(n_515), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g647 ( .A(n_515), .B(n_561), .Y(n_647) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g608 ( .A(n_516), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_521), .A2(n_611), .B1(n_650), .B2(n_651), .Y(n_649) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_536), .Y(n_521) );
INVx3_ASAP7_75t_L g583 ( .A(n_522), .Y(n_583) );
OR2x2_ASAP7_75t_L g716 ( .A(n_522), .B(n_592), .Y(n_716) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g589 ( .A(n_523), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g605 ( .A(n_523), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g613 ( .A(n_523), .B(n_561), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_523), .B(n_537), .Y(n_669) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g560 ( .A(n_524), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g564 ( .A(n_524), .B(n_537), .Y(n_564) );
AND2x2_ASAP7_75t_L g640 ( .A(n_524), .B(n_587), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_524), .B(n_546), .Y(n_680) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_536), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g596 ( .A(n_536), .B(n_557), .Y(n_596) );
AND2x2_ASAP7_75t_L g600 ( .A(n_536), .B(n_590), .Y(n_600) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_546), .Y(n_536) );
INVx3_ASAP7_75t_L g561 ( .A(n_537), .Y(n_561) );
AND2x2_ASAP7_75t_L g586 ( .A(n_537), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g721 ( .A(n_537), .B(n_704), .Y(n_721) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_546), .Y(n_575) );
INVx2_ASAP7_75t_L g587 ( .A(n_546), .Y(n_587) );
AND2x2_ASAP7_75t_L g631 ( .A(n_546), .B(n_607), .Y(n_631) );
INVx1_ASAP7_75t_L g674 ( .A(n_546), .Y(n_674) );
OR2x2_ASAP7_75t_L g705 ( .A(n_546), .B(n_607), .Y(n_705) );
AND2x2_ASAP7_75t_L g725 ( .A(n_546), .B(n_561), .Y(n_725) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_558), .B(n_562), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g563 ( .A(n_557), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_557), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g682 ( .A(n_559), .Y(n_682) );
INVx2_ASAP7_75t_SL g576 ( .A(n_560), .Y(n_576) );
AND2x2_ASAP7_75t_L g696 ( .A(n_560), .B(n_590), .Y(n_696) );
INVx2_ASAP7_75t_L g642 ( .A(n_561), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_561), .B(n_674), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_565), .B1(n_568), .B2(n_574), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_564), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g730 ( .A(n_564), .Y(n_730) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g655 ( .A(n_566), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_566), .B(n_598), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_567), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g671 ( .A(n_567), .B(n_620), .Y(n_671) );
INVx2_ASAP7_75t_L g727 ( .A(n_567), .Y(n_727) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AND2x2_ASAP7_75t_L g597 ( .A(n_570), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_570), .B(n_615), .Y(n_648) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_572), .B(n_592), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g709 ( .A(n_575), .Y(n_709) );
O2A1O1Ixp33_ASAP7_75t_SL g659 ( .A1(n_576), .A2(n_660), .B(n_662), .C(n_665), .Y(n_659) );
OR2x2_ASAP7_75t_L g686 ( .A(n_576), .B(n_590), .Y(n_686) );
OAI221xp5_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_582), .B1(n_584), .B2(n_591), .C(n_594), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_579), .B(n_581), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_579), .B(n_628), .Y(n_635) );
AND2x2_ASAP7_75t_L g677 ( .A(n_579), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g713 ( .A(n_579), .Y(n_713) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_580), .Y(n_604) );
INVx1_ASAP7_75t_L g617 ( .A(n_580), .Y(n_617) );
NOR2xp67_ASAP7_75t_L g637 ( .A(n_583), .B(n_638), .Y(n_637) );
INVxp67_ASAP7_75t_L g691 ( .A(n_583), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_583), .B(n_631), .Y(n_707) );
INVx2_ASAP7_75t_L g693 ( .A(n_584), .Y(n_693) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g634 ( .A(n_586), .B(n_605), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_586), .A2(n_602), .B(n_644), .C(n_645), .Y(n_643) );
AND2x2_ASAP7_75t_L g612 ( .A(n_587), .B(n_607), .Y(n_612) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_591), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
OR2x2_ASAP7_75t_L g660 ( .A(n_592), .B(n_661), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_597), .B2(n_600), .Y(n_594) );
INVx1_ASAP7_75t_L g714 ( .A(n_596), .Y(n_714) );
INVx1_ASAP7_75t_L g661 ( .A(n_598), .Y(n_661) );
INVx1_ASAP7_75t_L g712 ( .A(n_600), .Y(n_712) );
AOI211xp5_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_605), .B(n_609), .C(n_632), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g624 ( .A(n_604), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g675 ( .A(n_605), .Y(n_675) );
AND2x2_ASAP7_75t_L g724 ( .A(n_605), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI21xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_614), .B(n_622), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx2_ASAP7_75t_L g638 ( .A(n_612), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_612), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g630 ( .A(n_613), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g706 ( .A(n_613), .Y(n_706) );
OAI32xp33_ASAP7_75t_L g717 ( .A1(n_613), .A2(n_665), .A3(n_672), .B1(n_713), .B2(n_718), .Y(n_717) );
NOR2xp33_ASAP7_75t_SL g614 ( .A(n_615), .B(n_618), .Y(n_614) );
INVx1_ASAP7_75t_SL g685 ( .A(n_615), .Y(n_685) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g625 ( .A(n_621), .Y(n_625) );
OAI21xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B(n_630), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_624), .A2(n_672), .B1(n_698), .B2(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_628), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g665 ( .A(n_631), .Y(n_665) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2x1p5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g658 ( .A(n_642), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_648), .B(n_649), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_651), .A2(n_693), .B1(n_694), .B2(n_696), .C(n_697), .Y(n_692) );
NAND5xp2_ASAP7_75t_L g652 ( .A(n_653), .B(n_676), .C(n_692), .D(n_702), .E(n_720), .Y(n_652) );
AOI211xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_656), .B(n_659), .C(n_666), .Y(n_653) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g723 ( .A(n_660), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_670), .B2(n_672), .Y(n_666) );
INVx1_ASAP7_75t_SL g699 ( .A(n_669), .Y(n_699) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI322xp33_ASAP7_75t_L g681 ( .A1(n_672), .A2(n_682), .A3(n_683), .B1(n_684), .B2(n_685), .C1(n_686), .C2(n_687), .Y(n_681) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVx1_ASAP7_75t_L g684 ( .A(n_674), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_674), .B(n_699), .Y(n_698) );
AOI211xp5_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_679), .B(n_681), .C(n_689), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_685), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_711) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g728 ( .A(n_695), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_710), .B1(n_711), .B2(n_715), .C(n_717), .Y(n_702) );
OAI211xp5_ASAP7_75t_SL g703 ( .A1(n_704), .A2(n_706), .B(n_707), .C(n_708), .Y(n_703) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g729 ( .A(n_705), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_723), .B2(n_724), .C(n_726), .Y(n_720) );
AOI21xp33_ASAP7_75t_SL g726 ( .A1(n_727), .A2(n_728), .B(n_729), .Y(n_726) );
CKINVDCx16_ASAP7_75t_R g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
endmodule