module fake_jpeg_21671_n_163 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_163);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_18),
.C(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_22),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_25),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_47),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_48),
.B(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_18),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_36),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_46),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_17),
.B1(n_31),
.B2(n_25),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_66),
.B1(n_31),
.B2(n_19),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_29),
.B(n_23),
.C(n_19),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_29),
.B(n_24),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_17),
.B1(n_22),
.B2(n_24),
.Y(n_66)
);

HAxp5_ASAP7_75t_SL g68 ( 
.A(n_65),
.B(n_29),
.CON(n_68),
.SN(n_68)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_68),
.B(n_75),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_79),
.B1(n_61),
.B2(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_30),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_80),
.B(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_30),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_26),
.B1(n_28),
.B2(n_44),
.Y(n_79)
);

HAxp5_ASAP7_75t_SL g80 ( 
.A(n_50),
.B(n_23),
.CON(n_80),
.SN(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_14),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_84),
.B(n_86),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_44),
.B(n_38),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_13),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_52),
.B1(n_60),
.B2(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_95),
.B1(n_106),
.B2(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_52),
.B1(n_60),
.B2(n_53),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_67),
.C(n_34),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_88),
.C(n_84),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_70),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_52),
.B1(n_54),
.B2(n_43),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_111),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_88),
.C(n_90),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_117),
.B(n_102),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_93),
.C(n_98),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_116),
.C(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_90),
.C(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_89),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_74),
.B1(n_72),
.B2(n_85),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_125),
.C(n_127),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_94),
.B(n_104),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_122),
.A2(n_128),
.B(n_117),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_110),
.C(n_108),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_15),
.A3(n_14),
.B1(n_12),
.B2(n_11),
.C1(n_9),
.C2(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_28),
.C(n_26),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_139),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_124),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_136),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_107),
.B1(n_85),
.B2(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_82),
.B(n_97),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_97),
.B1(n_101),
.B2(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_138),
.Y(n_146)
);

OAI321xp33_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_87),
.A3(n_103),
.B1(n_69),
.B2(n_11),
.C(n_32),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_121),
.C(n_125),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_28),
.B1(n_26),
.B2(n_54),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_122),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_133),
.Y(n_149)
);

AOI21x1_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_1),
.B(n_2),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_144),
.A2(n_147),
.B(n_5),
.Y(n_152)
);

AOI321xp33_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_152),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_139),
.B(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_146),
.B(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_6),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_153),
.B(n_154),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_143),
.B(n_6),
.Y(n_154)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_151),
.B(n_141),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_155),
.B(n_156),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_148),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_158),
.C(n_69),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.Y(n_163)
);


endmodule