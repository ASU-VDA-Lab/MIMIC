module fake_jpeg_10338_n_253 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_37),
.Y(n_53)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_0),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_24),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_49),
.B(n_56),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_30),
.B(n_29),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_51),
.A2(n_55),
.B(n_59),
.C(n_53),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_62),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_30),
.B1(n_37),
.B2(n_26),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_55),
.B1(n_24),
.B2(n_33),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_28),
.B(n_18),
.C(n_23),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_34),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_30),
.B1(n_37),
.B2(n_26),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_45),
.B1(n_33),
.B2(n_24),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_32),
.B1(n_27),
.B2(n_23),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_22),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_32),
.B1(n_27),
.B2(n_23),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_27),
.B1(n_17),
.B2(n_18),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_41),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_43),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_17),
.Y(n_66)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_20),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_35),
.A2(n_27),
.B1(n_17),
.B2(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_21),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_71),
.B(n_87),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_73),
.A2(n_91),
.B(n_92),
.Y(n_116)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_81),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_75),
.B(n_5),
.Y(n_124)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_31),
.B1(n_25),
.B2(n_19),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_20),
.B1(n_19),
.B2(n_25),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_78),
.A2(n_82),
.B1(n_100),
.B2(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_45),
.B1(n_35),
.B2(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_22),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_96),
.Y(n_106)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_93),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_65),
.B(n_47),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_21),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_22),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_1),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_95),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_1),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_41),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_97),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_33),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_65),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_70),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_2),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_114),
.B(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_72),
.B(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_124),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_112),
.B(n_92),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_53),
.B(n_54),
.Y(n_114)
);

AOI32xp33_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_50),
.A3(n_60),
.B1(n_9),
.B2(n_10),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_127),
.B1(n_101),
.B2(n_102),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_129),
.Y(n_133)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_72),
.B(n_11),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_100),
.C(n_83),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_132),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_91),
.B1(n_88),
.B2(n_80),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_141),
.Y(n_171)
);

AO21x2_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_73),
.B(n_82),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_138),
.B1(n_144),
.B2(n_151),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_89),
.B1(n_84),
.B2(n_75),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_85),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_89),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_103),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_143),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_123),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_73),
.B1(n_94),
.B2(n_83),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_103),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_147),
.A2(n_155),
.B(n_156),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_152),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_76),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_154),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_126),
.B1(n_116),
.B2(n_108),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_92),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_157),
.A2(n_121),
.B(n_119),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_166),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_151),
.A2(n_112),
.B(n_116),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_164),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_119),
.B(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_149),
.B(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_179),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_74),
.B1(n_111),
.B2(n_105),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_118),
.B1(n_136),
.B2(n_143),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_118),
.B1(n_111),
.B2(n_99),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_177),
.A2(n_134),
.B1(n_139),
.B2(n_131),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_144),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_137),
.C(n_147),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_135),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_187),
.C(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_136),
.B1(n_155),
.B2(n_154),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_186),
.A2(n_191),
.B1(n_171),
.B2(n_177),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_135),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_196),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_131),
.C(n_153),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_159),
.C(n_192),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_148),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_167),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_194),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_159),
.B(n_171),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_15),
.C(n_16),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_164),
.C(n_160),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

OA21x2_ASAP7_75t_SL g209 ( 
.A1(n_183),
.A2(n_185),
.B(n_187),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_SL g222 ( 
.A(n_209),
.B(n_197),
.C(n_178),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_190),
.C(n_191),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_211),
.A2(n_179),
.B1(n_175),
.B2(n_170),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_161),
.C(n_169),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.C(n_192),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_217),
.C(n_221),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_185),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_211),
.A2(n_197),
.B(n_165),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_219),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_158),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_222),
.C(n_210),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_178),
.C(n_172),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_212),
.C(n_214),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_206),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_203),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_203),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_208),
.B1(n_204),
.B2(n_201),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_226),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_200),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_232),
.B1(n_220),
.B2(n_222),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_223),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_SL g240 ( 
.A(n_231),
.B(n_168),
.C(n_207),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_219),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_236),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_239),
.Y(n_243)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_238),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_239),
.A2(n_227),
.B1(n_230),
.B2(n_226),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_242),
.A2(n_244),
.B1(n_243),
.B2(n_238),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_233),
.B(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_233),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_237),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_246),
.A2(n_242),
.B(n_166),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_248),
.Y(n_249)
);

OAI211xp5_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_249),
.B(n_198),
.C(n_16),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_12),
.B(n_13),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_13),
.Y(n_253)
);


endmodule