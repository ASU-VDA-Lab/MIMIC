module fake_netlist_1_12076_n_46 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_46);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_46;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_L g16 ( .A(n_14), .B(n_7), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_9), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_8), .B(n_6), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_0), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_5), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_1), .B(n_10), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_11), .B(n_3), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_4), .B(n_0), .Y(n_23) );
BUFx6f_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
INVx2_ASAP7_75t_SL g25 ( .A(n_19), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_17), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_18), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g28 ( .A(n_27), .Y(n_28) );
OAI21xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_18), .B(n_16), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_24), .Y(n_30) );
AND2x2_ASAP7_75t_SL g31 ( .A(n_28), .B(n_23), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_29), .B(n_25), .Y(n_32) );
INVx1_ASAP7_75t_SL g33 ( .A(n_31), .Y(n_33) );
NAND4xp25_ASAP7_75t_L g34 ( .A(n_32), .B(n_22), .C(n_21), .D(n_16), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_34), .B(n_24), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
OAI221xp5_ASAP7_75t_L g38 ( .A1(n_36), .A2(n_24), .B1(n_30), .B2(n_3), .C(n_1), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_35), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_37), .Y(n_40) );
O2A1O1Ixp5_ASAP7_75t_L g41 ( .A1(n_39), .A2(n_30), .B(n_24), .C(n_13), .Y(n_41) );
NAND3x1_ASAP7_75t_L g42 ( .A(n_38), .B(n_2), .C(n_12), .Y(n_42) );
HB1xp67_ASAP7_75t_L g43 ( .A(n_40), .Y(n_43) );
INVx1_ASAP7_75t_L g44 ( .A(n_41), .Y(n_44) );
OAI22xp33_ASAP7_75t_L g45 ( .A1(n_43), .A2(n_42), .B1(n_2), .B2(n_15), .Y(n_45) );
XNOR2xp5_ASAP7_75t_L g46 ( .A(n_45), .B(n_44), .Y(n_46) );
endmodule