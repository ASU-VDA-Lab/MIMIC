module fake_netlist_1_6603_n_1328 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1328);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1328;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_271;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_1321;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_272;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1271;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_270;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_269;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_274;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1219;
wire n_1120;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g269 ( .A(n_54), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_47), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_155), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_204), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_177), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_181), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_184), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_86), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_253), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_259), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g279 ( .A(n_159), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_137), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_206), .Y(n_281) );
INVxp67_ASAP7_75t_L g282 ( .A(n_161), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_32), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_200), .Y(n_284) );
CKINVDCx14_ASAP7_75t_R g285 ( .A(n_227), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_6), .Y(n_286) );
NOR2xp67_ASAP7_75t_L g287 ( .A(n_9), .B(n_256), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_29), .Y(n_288) );
INVxp33_ASAP7_75t_SL g289 ( .A(n_16), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_93), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_226), .Y(n_291) );
BUFx2_ASAP7_75t_SL g292 ( .A(n_170), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_176), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_57), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_205), .Y(n_295) );
INVxp67_ASAP7_75t_SL g296 ( .A(n_26), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_246), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_140), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_139), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_254), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_221), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_237), .Y(n_302) );
INVxp33_ASAP7_75t_L g303 ( .A(n_20), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_122), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_35), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_73), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_91), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_119), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_144), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_135), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_5), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_143), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_109), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_76), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_106), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_182), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_146), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_185), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_145), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_255), .Y(n_320) );
CKINVDCx16_ASAP7_75t_R g321 ( .A(n_207), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_223), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_82), .Y(n_323) );
INVxp67_ASAP7_75t_L g324 ( .A(n_78), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_250), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_53), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_131), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_154), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_104), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_43), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_64), .Y(n_331) );
CKINVDCx14_ASAP7_75t_R g332 ( .A(n_76), .Y(n_332) );
BUFx3_ASAP7_75t_L g333 ( .A(n_215), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_153), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_172), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_202), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_106), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_25), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_39), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_165), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_212), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_189), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_262), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_136), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_92), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_81), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_132), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_265), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_12), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_45), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_128), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_164), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_266), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_245), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_59), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_152), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_260), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_87), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_66), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_85), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_26), .Y(n_361) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_233), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_20), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_72), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_263), .Y(n_365) );
CKINVDCx16_ASAP7_75t_R g366 ( .A(n_99), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_121), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_123), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_174), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_126), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_231), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_103), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_129), .Y(n_373) );
CKINVDCx14_ASAP7_75t_R g374 ( .A(n_203), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_104), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_238), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_149), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_29), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_111), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_264), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_13), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_24), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_62), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_168), .Y(n_384) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_133), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_73), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_192), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_34), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_234), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_216), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_141), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_150), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_116), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_120), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_130), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_17), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_175), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_2), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_53), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_193), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_243), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_239), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_82), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_12), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_198), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_27), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_171), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_2), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_103), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_183), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_86), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_4), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_195), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_48), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_142), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_97), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_66), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_21), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_148), .Y(n_419) );
CKINVDCx16_ASAP7_75t_R g420 ( .A(n_107), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_125), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_99), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_32), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_197), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_92), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_371), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_371), .Y(n_427) );
OA21x2_ASAP7_75t_L g428 ( .A1(n_277), .A2(n_110), .B(n_108), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_332), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_371), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_366), .B(n_0), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_371), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_321), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_277), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_291), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_291), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_303), .B(n_0), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_356), .B(n_1), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_270), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_391), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_289), .A2(n_4), .B1(n_1), .B2(n_3), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_301), .B(n_3), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_350), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_295), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_289), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_280), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_350), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_363), .B(n_7), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_363), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_411), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_362), .B(n_8), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g452 ( .A1(n_276), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_411), .Y(n_453) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_280), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_295), .Y(n_455) );
OAI22xp5_ASAP7_75t_SL g456 ( .A1(n_276), .A2(n_13), .B1(n_10), .B2(n_11), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_312), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_310), .Y(n_458) );
INVx6_ASAP7_75t_L g459 ( .A(n_312), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_270), .A2(n_15), .B1(n_11), .B2(n_14), .Y(n_460) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_320), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_310), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_306), .Y(n_463) );
OR2x6_ASAP7_75t_L g464 ( .A(n_452), .B(n_292), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_429), .B(n_420), .Y(n_465) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_428), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_439), .Y(n_467) );
INVx4_ASAP7_75t_L g468 ( .A(n_448), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_448), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_446), .Y(n_470) );
BUFx4f_ASAP7_75t_L g471 ( .A(n_448), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_446), .Y(n_472) );
OAI22xp33_ASAP7_75t_L g473 ( .A1(n_431), .A2(n_288), .B1(n_307), .B2(n_283), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_440), .B(n_327), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_439), .B(n_285), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_459), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_448), .A2(n_286), .B1(n_290), .B2(n_269), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_438), .A2(n_305), .B1(n_314), .B2(n_294), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_446), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_438), .A2(n_315), .B1(n_331), .B2(n_326), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_459), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_434), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_433), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_440), .B(n_389), .Y(n_484) );
INVx4_ASAP7_75t_L g485 ( .A(n_459), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_438), .B(n_437), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_446), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_437), .B(n_298), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_446), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_451), .B(n_288), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_434), .Y(n_491) );
INVx4_ASAP7_75t_L g492 ( .A(n_459), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_446), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_451), .A2(n_279), .B1(n_297), .B2(n_275), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_431), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_452), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_434), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_435), .Y(n_498) );
OR2x6_ASAP7_75t_L g499 ( .A(n_456), .B(n_337), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_441), .A2(n_279), .B1(n_297), .B2(n_275), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_443), .B(n_391), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_446), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_443), .B(n_307), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_447), .B(n_282), .Y(n_504) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_428), .Y(n_505) );
OR2x6_ASAP7_75t_L g506 ( .A(n_442), .B(n_425), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_435), .Y(n_507) );
BUFx10_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_435), .Y(n_509) );
NOR2xp33_ASAP7_75t_SL g510 ( .A(n_442), .B(n_302), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_472), .Y(n_511) );
BUFx8_ASAP7_75t_SL g512 ( .A(n_483), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_488), .B(n_340), .Y(n_513) );
BUFx3_ASAP7_75t_L g514 ( .A(n_508), .Y(n_514) );
BUFx3_ASAP7_75t_L g515 ( .A(n_508), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_471), .B(n_271), .Y(n_516) );
NOR2x1p5_ASAP7_75t_L g517 ( .A(n_490), .B(n_311), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_501), .Y(n_518) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_466), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_501), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_501), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_501), .Y(n_522) );
INVxp67_ASAP7_75t_L g523 ( .A(n_467), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_472), .Y(n_524) );
OAI22xp5_ASAP7_75t_SL g525 ( .A1(n_496), .A2(n_330), .B1(n_422), .B2(n_329), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_506), .B(n_304), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_479), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_468), .Y(n_528) );
NOR2xp67_ASAP7_75t_L g529 ( .A(n_500), .B(n_441), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_465), .B(n_304), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_468), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_471), .A2(n_339), .B1(n_346), .B2(n_338), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_471), .B(n_272), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_506), .B(n_316), .Y(n_534) );
NOR2x1p5_ASAP7_75t_L g535 ( .A(n_475), .B(n_311), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_486), .B(n_316), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_495), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g538 ( .A1(n_473), .A2(n_324), .B(n_416), .C(n_436), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_506), .B(n_318), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_479), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_506), .B(n_318), .Y(n_541) );
NOR2xp67_ASAP7_75t_L g542 ( .A(n_500), .B(n_445), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_468), .B(n_273), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_502), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_475), .B(n_319), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_484), .B(n_468), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_503), .B(n_323), .Y(n_547) );
BUFx2_ASAP7_75t_L g548 ( .A(n_495), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_494), .B(n_445), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_502), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_470), .Y(n_551) );
BUFx3_ASAP7_75t_L g552 ( .A(n_508), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_510), .Y(n_553) );
BUFx12f_ASAP7_75t_L g554 ( .A(n_464), .Y(n_554) );
NAND2x1p5_ASAP7_75t_L g555 ( .A(n_469), .B(n_460), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_494), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_469), .A2(n_477), .B1(n_504), .B2(n_480), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_470), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_466), .B(n_505), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_478), .A2(n_302), .B1(n_394), .B2(n_379), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_491), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_474), .B(n_344), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_482), .B(n_428), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_470), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_466), .B(n_505), .Y(n_565) );
CKINVDCx14_ASAP7_75t_R g566 ( .A(n_464), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_491), .B(n_348), .Y(n_567) );
NAND2x1p5_ASAP7_75t_L g568 ( .A(n_482), .B(n_460), .Y(n_568) );
BUFx8_ASAP7_75t_L g569 ( .A(n_497), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_482), .A2(n_355), .B1(n_358), .B2(n_349), .Y(n_570) );
AND2x6_ASAP7_75t_SL g571 ( .A(n_499), .B(n_360), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_497), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_498), .B(n_354), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_498), .B(n_323), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_507), .B(n_354), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_507), .B(n_369), .Y(n_576) );
BUFx3_ASAP7_75t_L g577 ( .A(n_508), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_509), .B(n_369), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_509), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_482), .B(n_380), .Y(n_580) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_505), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_485), .B(n_387), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_476), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_466), .B(n_274), .Y(n_584) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_464), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_466), .A2(n_364), .B1(n_375), .B2(n_361), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_487), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_485), .B(n_392), .Y(n_588) );
INVx3_ASAP7_75t_L g589 ( .A(n_492), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_476), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_492), .B(n_392), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_464), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_481), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_481), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_464), .A2(n_345), .B1(n_372), .B2(n_359), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_505), .B(n_449), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_487), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_492), .B(n_395), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_492), .B(n_395), .Y(n_599) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_505), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_487), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_499), .B(n_345), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_489), .B(n_278), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_489), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_493), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_548), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_596), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_574), .B(n_359), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_523), .B(n_499), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_555), .B(n_499), .Y(n_610) );
OAI22xp5_ASAP7_75t_SL g611 ( .A1(n_537), .A2(n_499), .B1(n_329), .B2(n_422), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_556), .A2(n_330), .B1(n_396), .B2(n_381), .C(n_372), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_529), .A2(n_381), .B1(n_398), .B2(n_396), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_574), .B(n_398), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_596), .Y(n_615) );
OAI22x1_ASAP7_75t_L g616 ( .A1(n_560), .A2(n_404), .B1(n_423), .B2(n_296), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_542), .A2(n_444), .B1(n_455), .B2(n_436), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_547), .B(n_378), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_512), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_518), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_538), .A2(n_383), .B(n_386), .C(n_382), .Y(n_621) );
O2A1O1Ixp33_ASAP7_75t_L g622 ( .A1(n_549), .A2(n_399), .B(n_403), .C(n_388), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_519), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_520), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_555), .B(n_404), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_545), .B(n_423), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_557), .A2(n_444), .B1(n_455), .B2(n_436), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_547), .B(n_418), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g629 ( .A1(n_521), .A2(n_455), .B(n_458), .C(n_444), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_548), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_522), .B(n_458), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_514), .B(n_397), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_596), .Y(n_633) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_549), .A2(n_408), .B(n_409), .C(n_406), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_559), .A2(n_493), .B(n_385), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_559), .A2(n_284), .B(n_281), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_512), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_514), .B(n_397), .Y(n_638) );
OAI21xp5_ASAP7_75t_L g639 ( .A1(n_584), .A2(n_299), .B(n_293), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_569), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_586), .A2(n_462), .B1(n_458), .B2(n_414), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_565), .A2(n_308), .B(n_300), .Y(n_642) );
BUFx2_ASAP7_75t_L g643 ( .A(n_569), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_528), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_515), .B(n_405), .Y(n_645) );
BUFx3_ASAP7_75t_L g646 ( .A(n_569), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_531), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_517), .B(n_417), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_565), .A2(n_313), .B(n_309), .Y(n_649) );
INVx8_ASAP7_75t_L g650 ( .A(n_554), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_526), .B(n_405), .Y(n_651) );
CKINVDCx6p67_ASAP7_75t_R g652 ( .A(n_554), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_515), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_552), .B(n_410), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_535), .B(n_450), .Y(n_655) );
A2O1A1Ixp33_ASAP7_75t_L g656 ( .A1(n_561), .A2(n_287), .B(n_453), .C(n_450), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_534), .B(n_410), .Y(n_657) );
INVx8_ASAP7_75t_L g658 ( .A(n_571), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_595), .A2(n_415), .B1(n_421), .B2(n_374), .Y(n_659) );
INVx5_ASAP7_75t_L g660 ( .A(n_589), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_532), .A2(n_453), .B1(n_306), .B2(n_322), .Y(n_661) );
O2A1O1Ixp33_ASAP7_75t_SL g662 ( .A1(n_584), .A2(n_328), .B(n_334), .C(n_317), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_552), .B(n_421), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_543), .A2(n_336), .B(n_335), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_539), .B(n_341), .Y(n_665) );
OAI21x1_ASAP7_75t_L g666 ( .A1(n_563), .A2(n_384), .B(n_343), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_572), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_L g668 ( .A1(n_579), .A2(n_347), .B(n_352), .C(n_342), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_537), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_543), .A2(n_357), .B(n_353), .Y(n_670) );
NOR2xp33_ASAP7_75t_R g671 ( .A(n_566), .B(n_14), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g672 ( .A1(n_563), .A2(n_367), .B(n_365), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_546), .A2(n_373), .B(n_370), .Y(n_673) );
OAI22x1_ASAP7_75t_L g674 ( .A1(n_553), .A2(n_368), .B1(n_351), .B2(n_376), .Y(n_674) );
BUFx2_ASAP7_75t_L g675 ( .A(n_525), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_577), .B(n_377), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_568), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_602), .B(n_566), .Y(n_678) );
NAND2xp33_ASAP7_75t_SL g679 ( .A(n_592), .B(n_306), .Y(n_679) );
CKINVDCx11_ASAP7_75t_R g680 ( .A(n_577), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_516), .A2(n_393), .B(n_390), .Y(n_681) );
NOR2xp33_ASAP7_75t_R g682 ( .A(n_592), .B(n_15), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_602), .B(n_412), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_585), .B(n_401), .C(n_400), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_516), .A2(n_407), .B(n_402), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_530), .B(n_413), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_589), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_562), .B(n_412), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_533), .A2(n_424), .B(n_419), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_541), .B(n_384), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_568), .B(n_412), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_536), .B(n_412), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_580), .Y(n_693) );
BUFx12f_ASAP7_75t_L g694 ( .A(n_519), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_533), .A2(n_325), .B(n_320), .Y(n_695) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_567), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_573), .Y(n_697) );
AND2x4_ASAP7_75t_SL g698 ( .A(n_570), .B(n_454), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_575), .B(n_576), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_582), .A2(n_333), .B(n_325), .Y(n_700) );
BUFx2_ASAP7_75t_L g701 ( .A(n_588), .Y(n_701) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_578), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_583), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_590), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_SL g705 ( .A1(n_513), .A2(n_463), .B(n_426), .C(n_430), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_599), .B(n_16), .Y(n_706) );
OAI21xp33_ASAP7_75t_L g707 ( .A1(n_591), .A2(n_333), .B(n_454), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_593), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_594), .Y(n_709) );
INVxp67_ASAP7_75t_L g710 ( .A(n_598), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_519), .A2(n_457), .B(n_454), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_603), .A2(n_463), .B(n_427), .C(n_430), .Y(n_712) );
INVx3_ASAP7_75t_L g713 ( .A(n_519), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_551), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_551), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_519), .A2(n_457), .B(n_454), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_558), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_581), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_581), .B(n_457), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_581), .B(n_17), .Y(n_720) );
BUFx10_ASAP7_75t_L g721 ( .A(n_604), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_600), .A2(n_461), .B1(n_457), .B2(n_463), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_600), .B(n_18), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_600), .B(n_457), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_600), .B(n_18), .Y(n_725) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_600), .Y(n_726) );
AOI33xp33_ASAP7_75t_L g727 ( .A1(n_511), .A2(n_426), .A3(n_427), .B1(n_430), .B2(n_432), .B3(n_24), .Y(n_727) );
INVx4_ASAP7_75t_L g728 ( .A(n_564), .Y(n_728) );
INVxp67_ASAP7_75t_L g729 ( .A(n_587), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_597), .A2(n_461), .B(n_432), .Y(n_730) );
AOI21x1_ASAP7_75t_L g731 ( .A1(n_597), .A2(n_432), .B(n_461), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_601), .B(n_461), .Y(n_732) );
NOR3xp33_ASAP7_75t_L g733 ( .A(n_601), .B(n_463), .C(n_19), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_605), .B(n_461), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_605), .A2(n_22), .B1(n_19), .B2(n_21), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g736 ( .A1(n_511), .A2(n_25), .B(n_22), .C(n_23), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_524), .B(n_23), .Y(n_737) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_527), .Y(n_738) );
BUFx2_ASAP7_75t_L g739 ( .A(n_540), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_540), .A2(n_113), .B(n_112), .Y(n_740) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_544), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_550), .A2(n_27), .B1(n_28), .B2(n_30), .Y(n_742) );
AOI21x1_ASAP7_75t_L g743 ( .A1(n_559), .A2(n_115), .B(n_114), .Y(n_743) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_537), .A2(n_28), .B1(n_30), .B2(n_31), .Y(n_744) );
BUFx12f_ASAP7_75t_L g745 ( .A(n_619), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_699), .A2(n_118), .B(n_117), .Y(n_746) );
AO31x2_ASAP7_75t_L g747 ( .A1(n_627), .A2(n_31), .A3(n_33), .B(n_34), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_683), .Y(n_748) );
INVx2_ASAP7_75t_SL g749 ( .A(n_646), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_691), .Y(n_750) );
AO31x2_ASAP7_75t_L g751 ( .A1(n_627), .A2(n_33), .A3(n_35), .B(n_36), .Y(n_751) );
INVxp67_ASAP7_75t_L g752 ( .A(n_606), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_667), .Y(n_753) );
AO31x2_ASAP7_75t_L g754 ( .A1(n_656), .A2(n_37), .A3(n_38), .B(n_40), .Y(n_754) );
OR2x6_ASAP7_75t_L g755 ( .A(n_643), .B(n_41), .Y(n_755) );
AOI21xp33_ASAP7_75t_L g756 ( .A1(n_625), .A2(n_628), .B(n_614), .Y(n_756) );
O2A1O1Ixp33_ASAP7_75t_L g757 ( .A1(n_617), .A2(n_42), .B(n_43), .C(n_44), .Y(n_757) );
OAI21xp5_ASAP7_75t_L g758 ( .A1(n_672), .A2(n_127), .B(n_124), .Y(n_758) );
O2A1O1Ixp33_ASAP7_75t_L g759 ( .A1(n_622), .A2(n_44), .B(n_45), .C(n_46), .Y(n_759) );
AOI221x1_ASAP7_75t_L g760 ( .A1(n_674), .A2(n_46), .B1(n_47), .B2(n_48), .C(n_49), .Y(n_760) );
CKINVDCx5p33_ASAP7_75t_R g761 ( .A(n_637), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_608), .B(n_614), .Y(n_762) );
NOR2xp33_ASAP7_75t_SL g763 ( .A(n_640), .B(n_49), .Y(n_763) );
AND2x4_ASAP7_75t_L g764 ( .A(n_677), .B(n_50), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_608), .B(n_50), .Y(n_765) );
OAI21xp5_ASAP7_75t_L g766 ( .A1(n_636), .A2(n_138), .B(n_134), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_607), .Y(n_767) );
O2A1O1Ixp33_ASAP7_75t_SL g768 ( .A1(n_705), .A2(n_191), .B(n_268), .C(n_267), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_688), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_675), .A2(n_51), .B1(n_52), .B2(n_54), .Y(n_770) );
INVx8_ASAP7_75t_L g771 ( .A(n_650), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_615), .Y(n_772) );
AOI32xp33_ASAP7_75t_L g773 ( .A1(n_610), .A2(n_51), .A3(n_52), .B1(n_55), .B2(n_56), .Y(n_773) );
OAI22xp5_ASAP7_75t_SL g774 ( .A1(n_611), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_774) );
BUFx3_ASAP7_75t_L g775 ( .A(n_680), .Y(n_775) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_630), .Y(n_776) );
O2A1O1Ixp33_ASAP7_75t_L g777 ( .A1(n_634), .A2(n_58), .B(n_59), .C(n_60), .Y(n_777) );
NOR2x1_ASAP7_75t_R g778 ( .A(n_671), .B(n_58), .Y(n_778) );
A2O1A1Ixp33_ASAP7_75t_L g779 ( .A1(n_706), .A2(n_61), .B(n_62), .C(n_63), .Y(n_779) );
INVx4_ASAP7_75t_L g780 ( .A(n_694), .Y(n_780) );
OAI22xp33_ASAP7_75t_L g781 ( .A1(n_616), .A2(n_61), .B1(n_63), .B2(n_64), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_609), .A2(n_65), .B1(n_67), .B2(n_68), .Y(n_782) );
AOI22xp33_ASAP7_75t_SL g783 ( .A1(n_682), .A2(n_65), .B1(n_67), .B2(n_68), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g784 ( .A1(n_710), .A2(n_69), .B1(n_70), .B2(n_71), .Y(n_784) );
OA21x2_ASAP7_75t_L g785 ( .A1(n_666), .A2(n_201), .B(n_261), .Y(n_785) );
A2O1A1Ixp33_ASAP7_75t_L g786 ( .A1(n_686), .A2(n_69), .B(n_70), .C(n_71), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_612), .A2(n_72), .B1(n_74), .B2(n_75), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_652), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_644), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_633), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_696), .A2(n_74), .B1(n_75), .B2(n_77), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_647), .Y(n_792) );
INVx4_ASAP7_75t_L g793 ( .A(n_650), .Y(n_793) );
A2O1A1Ixp33_ASAP7_75t_L g794 ( .A1(n_673), .A2(n_727), .B(n_621), .C(n_690), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_631), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_714), .Y(n_796) );
INVxp67_ASAP7_75t_SL g797 ( .A(n_741), .Y(n_797) );
A2O1A1Ixp33_ASAP7_75t_L g798 ( .A1(n_690), .A2(n_77), .B(n_78), .C(n_79), .Y(n_798) );
A2O1A1Ixp33_ASAP7_75t_L g799 ( .A1(n_664), .A2(n_79), .B(n_80), .C(n_81), .Y(n_799) );
AO32x2_ASAP7_75t_L g800 ( .A1(n_661), .A2(n_80), .A3(n_83), .B1(n_84), .B2(n_85), .Y(n_800) );
INVxp67_ASAP7_75t_L g801 ( .A(n_702), .Y(n_801) );
OAI21xp5_ASAP7_75t_L g802 ( .A1(n_642), .A2(n_209), .B(n_258), .Y(n_802) );
INVx2_ASAP7_75t_SL g803 ( .A(n_650), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_618), .A2(n_83), .B1(n_84), .B2(n_87), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_620), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_649), .A2(n_211), .B(n_257), .Y(n_806) );
A2O1A1Ixp33_ASAP7_75t_L g807 ( .A1(n_670), .A2(n_88), .B(n_89), .C(n_90), .Y(n_807) );
O2A1O1Ixp33_ASAP7_75t_L g808 ( .A1(n_668), .A2(n_88), .B(n_89), .C(n_90), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_618), .B(n_91), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_669), .B(n_93), .Y(n_810) );
AO32x2_ASAP7_75t_L g811 ( .A1(n_661), .A2(n_94), .A3(n_95), .B1(n_96), .B2(n_97), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_631), .Y(n_812) );
NOR2xp33_ASAP7_75t_SL g813 ( .A(n_658), .B(n_94), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_613), .B(n_95), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_715), .Y(n_815) );
OR2x2_ASAP7_75t_L g816 ( .A(n_678), .B(n_98), .Y(n_816) );
A2O1A1Ixp33_ASAP7_75t_L g817 ( .A1(n_681), .A2(n_98), .B(n_100), .C(n_101), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_655), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_626), .B(n_102), .Y(n_819) );
AND2x4_ASAP7_75t_L g820 ( .A(n_655), .B(n_701), .Y(n_820) );
A2O1A1Ixp33_ASAP7_75t_L g821 ( .A1(n_685), .A2(n_105), .B(n_147), .C(n_151), .Y(n_821) );
A2O1A1Ixp33_ASAP7_75t_L g822 ( .A1(n_689), .A2(n_105), .B(n_156), .C(n_157), .Y(n_822) );
OR2x2_ASAP7_75t_L g823 ( .A(n_658), .B(n_158), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_717), .Y(n_824) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_623), .Y(n_825) );
OAI22xp33_ASAP7_75t_L g826 ( .A1(n_659), .A2(n_160), .B1(n_162), .B2(n_163), .Y(n_826) );
NOR2xp33_ASAP7_75t_SL g827 ( .A(n_658), .B(n_166), .Y(n_827) );
BUFx3_ASAP7_75t_L g828 ( .A(n_721), .Y(n_828) );
AO31x2_ASAP7_75t_L g829 ( .A1(n_720), .A2(n_167), .A3(n_169), .B(n_173), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_684), .B(n_624), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_651), .B(n_178), .Y(n_831) );
AOI221x1_ASAP7_75t_L g832 ( .A1(n_733), .A2(n_179), .B1(n_180), .B2(n_186), .C(n_187), .Y(n_832) );
OAI21xp5_ASAP7_75t_L g833 ( .A1(n_639), .A2(n_188), .B(n_190), .Y(n_833) );
AOI21xp5_ASAP7_75t_L g834 ( .A1(n_719), .A2(n_194), .B(n_196), .Y(n_834) );
OR2x2_ASAP7_75t_L g835 ( .A(n_648), .B(n_199), .Y(n_835) );
AOI21xp5_ASAP7_75t_L g836 ( .A1(n_724), .A2(n_208), .B(n_210), .Y(n_836) );
OA21x2_ASAP7_75t_L g837 ( .A1(n_724), .A2(n_213), .B(n_214), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_739), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_648), .B(n_217), .Y(n_839) );
INVx3_ASAP7_75t_L g840 ( .A(n_721), .Y(n_840) );
BUFx8_ASAP7_75t_L g841 ( .A(n_709), .Y(n_841) );
AO31x2_ASAP7_75t_L g842 ( .A1(n_723), .A2(n_218), .A3(n_219), .B(n_220), .Y(n_842) );
INVx1_ASAP7_75t_SL g843 ( .A(n_737), .Y(n_843) );
NAND2xp5_ASAP7_75t_SL g844 ( .A(n_653), .B(n_222), .Y(n_844) );
A2O1A1Ixp33_ASAP7_75t_L g845 ( .A1(n_665), .A2(n_224), .B(n_225), .C(n_228), .Y(n_845) );
OAI21xp5_ASAP7_75t_L g846 ( .A1(n_635), .A2(n_229), .B(n_230), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_651), .B(n_232), .Y(n_847) );
BUFx2_ASAP7_75t_SL g848 ( .A(n_660), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_657), .B(n_235), .Y(n_849) );
BUFx6f_ASAP7_75t_L g850 ( .A(n_623), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_657), .B(n_236), .Y(n_851) );
INVx3_ASAP7_75t_SL g852 ( .A(n_660), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_744), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_665), .A2(n_240), .B1(n_241), .B2(n_242), .Y(n_854) );
AOI221x1_ASAP7_75t_L g855 ( .A1(n_707), .A2(n_244), .B1(n_247), .B2(n_248), .C(n_249), .Y(n_855) );
BUFx10_ASAP7_75t_L g856 ( .A(n_692), .Y(n_856) );
OAI21xp5_ASAP7_75t_L g857 ( .A1(n_729), .A2(n_251), .B(n_252), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_703), .Y(n_858) );
CKINVDCx11_ASAP7_75t_R g859 ( .A(n_687), .Y(n_859) );
AO32x2_ASAP7_75t_L g860 ( .A1(n_641), .A2(n_722), .A3(n_728), .B1(n_718), .B2(n_736), .Y(n_860) );
NOR2xp33_ASAP7_75t_R g861 ( .A(n_679), .B(n_653), .Y(n_861) );
BUFx2_ASAP7_75t_SL g862 ( .A(n_660), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_708), .Y(n_863) );
AOI21xp5_ASAP7_75t_L g864 ( .A1(n_726), .A2(n_700), .B(n_711), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_716), .A2(n_734), .B(n_732), .Y(n_865) );
BUFx2_ASAP7_75t_L g866 ( .A(n_660), .Y(n_866) );
AO31x2_ASAP7_75t_L g867 ( .A1(n_725), .A2(n_722), .A3(n_641), .B(n_732), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_704), .A2(n_676), .B1(n_735), .B2(n_742), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_632), .B(n_638), .Y(n_869) );
BUFx2_ASAP7_75t_L g870 ( .A(n_704), .Y(n_870) );
AO31x2_ASAP7_75t_L g871 ( .A1(n_734), .A2(n_740), .A3(n_730), .B(n_695), .Y(n_871) );
AOI21xp33_ASAP7_75t_L g872 ( .A1(n_645), .A2(n_654), .B(n_663), .Y(n_872) );
A2O1A1Ixp33_ASAP7_75t_L g873 ( .A1(n_712), .A2(n_698), .B(n_713), .C(n_738), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_662), .Y(n_874) );
OAI21xp5_ASAP7_75t_L g875 ( .A1(n_743), .A2(n_731), .B(n_713), .Y(n_875) );
O2A1O1Ixp33_ASAP7_75t_SL g876 ( .A1(n_738), .A2(n_705), .B(n_629), .C(n_672), .Y(n_876) );
BUFx6f_ASAP7_75t_L g877 ( .A(n_738), .Y(n_877) );
INVx3_ASAP7_75t_L g878 ( .A(n_694), .Y(n_878) );
BUFx12f_ASAP7_75t_L g879 ( .A(n_619), .Y(n_879) );
AOI221xp5_ASAP7_75t_L g880 ( .A1(n_622), .A2(n_634), .B1(n_618), .B2(n_628), .C(n_616), .Y(n_880) );
A2O1A1Ixp33_ASAP7_75t_L g881 ( .A1(n_699), .A2(n_697), .B(n_693), .C(n_706), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_608), .B(n_574), .Y(n_882) );
INVx4_ASAP7_75t_L g883 ( .A(n_646), .Y(n_883) );
AND2x4_ASAP7_75t_L g884 ( .A(n_640), .B(n_646), .Y(n_884) );
BUFx10_ASAP7_75t_L g885 ( .A(n_640), .Y(n_885) );
AOI21xp33_ASAP7_75t_L g886 ( .A1(n_625), .A2(n_523), .B(n_553), .Y(n_886) );
AO31x2_ASAP7_75t_L g887 ( .A1(n_627), .A2(n_656), .A3(n_617), .B(n_720), .Y(n_887) );
BUFx2_ASAP7_75t_L g888 ( .A(n_606), .Y(n_888) );
OR2x2_ASAP7_75t_L g889 ( .A(n_606), .B(n_523), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_880), .A2(n_756), .B1(n_774), .B2(n_810), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_858), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_820), .B(n_801), .Y(n_892) );
AOI22xp33_ASAP7_75t_SL g893 ( .A1(n_813), .A2(n_853), .B1(n_841), .B2(n_764), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_863), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_753), .Y(n_895) );
BUFx2_ASAP7_75t_L g896 ( .A(n_841), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_795), .B(n_812), .Y(n_897) );
AND2x4_ASAP7_75t_L g898 ( .A(n_828), .B(n_793), .Y(n_898) );
BUFx6f_ASAP7_75t_L g899 ( .A(n_825), .Y(n_899) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_762), .A2(n_882), .B1(n_773), .B2(n_886), .C(n_781), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_843), .A2(n_797), .B1(n_764), .B2(n_794), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_789), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_816), .A2(n_835), .B1(n_787), .B2(n_830), .Y(n_903) );
INVx2_ASAP7_75t_L g904 ( .A(n_796), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_805), .B(n_792), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_805), .Y(n_906) );
INVx2_ASAP7_75t_SL g907 ( .A(n_771), .Y(n_907) );
OAI21xp5_ASAP7_75t_L g908 ( .A1(n_765), .A2(n_769), .B(n_849), .Y(n_908) );
AOI21xp5_ASAP7_75t_L g909 ( .A1(n_876), .A2(n_847), .B(n_831), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_815), .Y(n_910) );
OAI21x1_ASAP7_75t_L g911 ( .A1(n_785), .A2(n_837), .B(n_836), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_750), .B(n_748), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_838), .B(n_887), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g914 ( .A(n_820), .B(n_889), .Y(n_914) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_851), .A2(n_873), .B(n_768), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_887), .B(n_824), .Y(n_916) );
OR2x6_ASAP7_75t_L g917 ( .A(n_771), .B(n_793), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_887), .B(n_767), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_772), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_790), .B(n_819), .Y(n_920) );
OR2x2_ASAP7_75t_L g921 ( .A(n_888), .B(n_776), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_791), .Y(n_922) );
HB1xp67_ASAP7_75t_L g923 ( .A(n_752), .Y(n_923) );
HB1xp67_ASAP7_75t_L g924 ( .A(n_755), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_809), .Y(n_925) );
AO31x2_ASAP7_75t_L g926 ( .A1(n_760), .A2(n_845), .A3(n_854), .B(n_798), .Y(n_926) );
A2O1A1Ixp33_ASAP7_75t_L g927 ( .A1(n_759), .A2(n_777), .B(n_757), .C(n_808), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_784), .Y(n_928) );
AOI22xp33_ASAP7_75t_SL g929 ( .A1(n_763), .A2(n_755), .B1(n_827), .B2(n_839), .Y(n_929) );
OA21x2_ASAP7_75t_L g930 ( .A1(n_857), .A2(n_833), .B(n_846), .Y(n_930) );
NAND2xp5_ASAP7_75t_SL g931 ( .A(n_840), .B(n_878), .Y(n_931) );
OR2x6_ASAP7_75t_L g932 ( .A(n_780), .B(n_848), .Y(n_932) );
OA21x2_ASAP7_75t_L g933 ( .A1(n_766), .A2(n_806), .B(n_802), .Y(n_933) );
OA21x2_ASAP7_75t_L g934 ( .A1(n_746), .A2(n_874), .B(n_834), .Y(n_934) );
OA21x2_ASAP7_75t_L g935 ( .A1(n_821), .A2(n_822), .B(n_844), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_747), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_747), .Y(n_937) );
BUFx8_ASAP7_75t_L g938 ( .A(n_745), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_751), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_751), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_859), .A2(n_840), .B1(n_814), .B2(n_870), .Y(n_941) );
INVx4_ASAP7_75t_L g942 ( .A(n_780), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_871), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_800), .Y(n_944) );
OAI21x1_ASAP7_75t_L g945 ( .A1(n_878), .A2(n_825), .B(n_850), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_803), .B(n_884), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_804), .A2(n_782), .B1(n_818), .B2(n_786), .Y(n_947) );
O2A1O1Ixp33_ASAP7_75t_L g948 ( .A1(n_779), .A2(n_817), .B(n_807), .C(n_799), .Y(n_948) );
NOR2x1_ASAP7_75t_SL g949 ( .A(n_862), .B(n_883), .Y(n_949) );
AO31x2_ASAP7_75t_L g950 ( .A1(n_860), .A2(n_867), .A3(n_869), .B(n_866), .Y(n_950) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_788), .Y(n_951) );
AND2x4_ASAP7_75t_L g952 ( .A(n_883), .B(n_884), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_852), .B(n_872), .Y(n_953) );
INVx6_ASAP7_75t_L g954 ( .A(n_885), .Y(n_954) );
INVxp67_ASAP7_75t_L g955 ( .A(n_778), .Y(n_955) );
OAI22xp33_ASAP7_75t_L g956 ( .A1(n_823), .A2(n_775), .B1(n_749), .B2(n_761), .Y(n_956) );
A2O1A1Ixp33_ASAP7_75t_L g957 ( .A1(n_770), .A2(n_783), .B(n_877), .C(n_860), .Y(n_957) );
A2O1A1Ixp33_ASAP7_75t_L g958 ( .A1(n_877), .A2(n_860), .B(n_850), .C(n_811), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_800), .Y(n_959) );
OAI21x1_ASAP7_75t_L g960 ( .A1(n_829), .A2(n_842), .B(n_861), .Y(n_960) );
AOI221xp5_ASAP7_75t_L g961 ( .A1(n_811), .A2(n_754), .B1(n_879), .B2(n_856), .C(n_842), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_754), .B(n_829), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_858), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_858), .Y(n_964) );
A2O1A1Ixp33_ASAP7_75t_L g965 ( .A1(n_881), .A2(n_819), .B(n_794), .C(n_756), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_880), .A2(n_529), .B1(n_542), .B2(n_675), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_795), .B(n_812), .Y(n_967) );
NAND2xp5_ASAP7_75t_SL g968 ( .A(n_841), .B(n_569), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_820), .B(n_523), .Y(n_969) );
NOR2xp33_ASAP7_75t_SL g970 ( .A(n_827), .B(n_569), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_841), .Y(n_971) );
AO21x1_ASAP7_75t_L g972 ( .A1(n_826), .A2(n_758), .B(n_868), .Y(n_972) );
OR2x2_ASAP7_75t_L g973 ( .A(n_889), .B(n_523), .Y(n_973) );
OR2x6_ASAP7_75t_L g974 ( .A(n_771), .B(n_793), .Y(n_974) );
A2O1A1Ixp33_ASAP7_75t_L g975 ( .A1(n_881), .A2(n_819), .B(n_794), .C(n_756), .Y(n_975) );
INVx2_ASAP7_75t_L g976 ( .A(n_753), .Y(n_976) );
AO31x2_ASAP7_75t_L g977 ( .A1(n_832), .A2(n_855), .A3(n_881), .B(n_865), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_795), .B(n_812), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g979 ( .A1(n_881), .A2(n_864), .B(n_875), .Y(n_979) );
INVxp67_ASAP7_75t_SL g980 ( .A(n_841), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_858), .Y(n_981) );
AO31x2_ASAP7_75t_L g982 ( .A1(n_832), .A2(n_855), .A3(n_881), .B(n_865), .Y(n_982) );
INVx3_ASAP7_75t_L g983 ( .A(n_828), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_795), .A2(n_812), .B1(n_881), .B2(n_843), .Y(n_984) );
INVx4_ASAP7_75t_L g985 ( .A(n_771), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_858), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_820), .B(n_523), .Y(n_987) );
INVx3_ASAP7_75t_L g988 ( .A(n_828), .Y(n_988) );
A2O1A1Ixp33_ASAP7_75t_L g989 ( .A1(n_881), .A2(n_819), .B(n_794), .C(n_756), .Y(n_989) );
AOI21xp5_ASAP7_75t_L g990 ( .A1(n_881), .A2(n_864), .B(n_875), .Y(n_990) );
OR2x2_ASAP7_75t_L g991 ( .A(n_889), .B(n_523), .Y(n_991) );
A2O1A1Ixp33_ASAP7_75t_L g992 ( .A1(n_881), .A2(n_819), .B(n_794), .C(n_756), .Y(n_992) );
OAI22xp33_ASAP7_75t_L g993 ( .A1(n_755), .A2(n_494), .B1(n_510), .B2(n_560), .Y(n_993) );
NAND2xp5_ASAP7_75t_SL g994 ( .A(n_841), .B(n_569), .Y(n_994) );
INVxp67_ASAP7_75t_L g995 ( .A(n_889), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_795), .B(n_812), .Y(n_996) );
AO31x2_ASAP7_75t_L g997 ( .A1(n_832), .A2(n_855), .A3(n_881), .B(n_865), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_795), .B(n_812), .Y(n_998) );
CKINVDCx6p67_ASAP7_75t_R g999 ( .A(n_771), .Y(n_999) );
AOI21xp5_ASAP7_75t_L g1000 ( .A1(n_881), .A2(n_864), .B(n_875), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_880), .A2(n_529), .B1(n_542), .B2(n_675), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_820), .B(n_523), .Y(n_1002) );
INVx3_ASAP7_75t_L g1003 ( .A(n_828), .Y(n_1003) );
NOR2xp33_ASAP7_75t_L g1004 ( .A(n_756), .B(n_556), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_880), .A2(n_529), .B1(n_542), .B2(n_675), .Y(n_1005) );
INVx2_ASAP7_75t_L g1006 ( .A(n_753), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_820), .B(n_523), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_795), .B(n_812), .Y(n_1008) );
BUFx3_ASAP7_75t_L g1009 ( .A(n_841), .Y(n_1009) );
HB1xp67_ASAP7_75t_L g1010 ( .A(n_921), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_897), .B(n_967), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_906), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_900), .A2(n_993), .B1(n_1004), .B2(n_966), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_943), .Y(n_1014) );
INVxp67_ASAP7_75t_SL g1015 ( .A(n_897), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g1016 ( .A(n_923), .Y(n_1016) );
INVx3_ASAP7_75t_L g1017 ( .A(n_899), .Y(n_1017) );
OA21x2_ASAP7_75t_L g1018 ( .A1(n_979), .A2(n_1000), .B(n_990), .Y(n_1018) );
OR2x2_ASAP7_75t_L g1019 ( .A(n_913), .B(n_905), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_967), .B(n_978), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_913), .Y(n_1021) );
OR2x6_ASAP7_75t_L g1022 ( .A(n_917), .B(n_974), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_978), .B(n_996), .Y(n_1023) );
OAI21xp5_ASAP7_75t_L g1024 ( .A1(n_927), .A2(n_975), .B(n_965), .Y(n_1024) );
OAI211xp5_ASAP7_75t_L g1025 ( .A1(n_929), .A2(n_893), .B(n_890), .C(n_1001), .Y(n_1025) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_932), .Y(n_1026) );
OR2x6_ASAP7_75t_L g1027 ( .A(n_917), .B(n_974), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_936), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_891), .Y(n_1029) );
BUFx3_ASAP7_75t_L g1030 ( .A(n_999), .Y(n_1030) );
OR2x2_ASAP7_75t_L g1031 ( .A(n_905), .B(n_996), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_998), .B(n_1008), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_937), .Y(n_1033) );
AOI221xp5_ASAP7_75t_L g1034 ( .A1(n_1005), .A2(n_903), .B1(n_900), .B2(n_984), .C(n_928), .Y(n_1034) );
HB1xp67_ASAP7_75t_L g1035 ( .A(n_932), .Y(n_1035) );
AND2x4_ASAP7_75t_L g1036 ( .A(n_998), .B(n_1008), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_904), .B(n_910), .Y(n_1037) );
CKINVDCx20_ASAP7_75t_R g1038 ( .A(n_938), .Y(n_1038) );
OA21x2_ASAP7_75t_L g1039 ( .A1(n_958), .A2(n_962), .B(n_960), .Y(n_1039) );
OA21x2_ASAP7_75t_L g1040 ( .A1(n_911), .A2(n_939), .B(n_940), .Y(n_1040) );
INVx2_ASAP7_75t_SL g1041 ( .A(n_917), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_918), .Y(n_1042) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_950), .B(n_984), .Y(n_1043) );
HB1xp67_ASAP7_75t_L g1044 ( .A(n_932), .Y(n_1044) );
OA21x2_ASAP7_75t_L g1045 ( .A1(n_909), .A2(n_916), .B(n_961), .Y(n_1045) );
OA21x2_ASAP7_75t_L g1046 ( .A1(n_916), .A2(n_961), .B(n_918), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_976), .B(n_1006), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_894), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_902), .Y(n_1049) );
OA21x2_ASAP7_75t_L g1050 ( .A1(n_944), .A2(n_959), .B(n_915), .Y(n_1050) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_950), .B(n_922), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_963), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_964), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_995), .B(n_973), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_903), .A2(n_947), .B1(n_970), .B2(n_972), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_981), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_986), .Y(n_1057) );
OR2x2_ASAP7_75t_L g1058 ( .A(n_950), .B(n_991), .Y(n_1058) );
OR2x6_ASAP7_75t_L g1059 ( .A(n_974), .B(n_968), .Y(n_1059) );
INVx2_ASAP7_75t_L g1060 ( .A(n_895), .Y(n_1060) );
OAI221xp5_ASAP7_75t_SL g1061 ( .A1(n_955), .A2(n_956), .B1(n_957), .B2(n_989), .C(n_992), .Y(n_1061) );
AOI21xp5_ASAP7_75t_SL g1062 ( .A1(n_901), .A2(n_930), .B(n_933), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_912), .Y(n_1063) );
INVx3_ASAP7_75t_L g1064 ( .A(n_945), .Y(n_1064) );
INVx2_ASAP7_75t_L g1065 ( .A(n_919), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_925), .B(n_912), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_908), .B(n_920), .Y(n_1067) );
BUFx3_ASAP7_75t_L g1068 ( .A(n_898), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_908), .B(n_920), .Y(n_1069) );
AOI21xp33_ASAP7_75t_L g1070 ( .A1(n_948), .A2(n_947), .B(n_953), .Y(n_1070) );
BUFx3_ASAP7_75t_L g1071 ( .A(n_898), .Y(n_1071) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_914), .B(n_969), .Y(n_1072) );
AOI221xp5_ASAP7_75t_L g1073 ( .A1(n_924), .A2(n_994), .B1(n_892), .B2(n_1007), .C(n_1002), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_977), .Y(n_1074) );
OR2x2_ASAP7_75t_L g1075 ( .A(n_987), .B(n_953), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_982), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_946), .B(n_952), .Y(n_1077) );
OR2x2_ASAP7_75t_L g1078 ( .A(n_983), .B(n_988), .Y(n_1078) );
OAI221xp5_ASAP7_75t_L g1079 ( .A1(n_941), .A2(n_970), .B1(n_980), .B2(n_896), .C(n_971), .Y(n_1079) );
INVx4_ASAP7_75t_R g1080 ( .A(n_1009), .Y(n_1080) );
BUFx2_ASAP7_75t_L g1081 ( .A(n_983), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_985), .B(n_907), .Y(n_1082) );
INVx4_ASAP7_75t_L g1083 ( .A(n_985), .Y(n_1083) );
AND2x4_ASAP7_75t_L g1084 ( .A(n_949), .B(n_1003), .Y(n_1084) );
AOI222xp33_ASAP7_75t_L g1085 ( .A1(n_938), .A2(n_951), .B1(n_942), .B2(n_931), .C1(n_954), .C2(n_988), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_926), .B(n_1003), .Y(n_1086) );
OR2x6_ASAP7_75t_L g1087 ( .A(n_954), .B(n_942), .Y(n_1087) );
INVx2_ASAP7_75t_L g1088 ( .A(n_997), .Y(n_1088) );
AO21x2_ASAP7_75t_L g1089 ( .A1(n_926), .A2(n_934), .B(n_935), .Y(n_1089) );
OR2x2_ASAP7_75t_L g1090 ( .A(n_935), .B(n_934), .Y(n_1090) );
INVx3_ASAP7_75t_L g1091 ( .A(n_899), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_906), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1011), .B(n_1020), .Y(n_1093) );
AND2x4_ASAP7_75t_L g1094 ( .A(n_1086), .B(n_1028), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1011), .B(n_1020), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1023), .B(n_1032), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1023), .B(n_1032), .Y(n_1097) );
INVxp67_ASAP7_75t_SL g1098 ( .A(n_1015), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1028), .Y(n_1099) );
INVx3_ASAP7_75t_SL g1100 ( .A(n_1022), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_1067), .B(n_1069), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1086), .B(n_1036), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1033), .Y(n_1103) );
AND2x4_ASAP7_75t_L g1104 ( .A(n_1033), .B(n_1042), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1042), .B(n_1021), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1036), .B(n_1067), .Y(n_1106) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_1014), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1036), .B(n_1069), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1012), .B(n_1092), .Y(n_1109) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_1031), .A2(n_1055), .B1(n_1013), .B2(n_1034), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1012), .B(n_1092), .Y(n_1111) );
BUFx3_ASAP7_75t_L g1112 ( .A(n_1022), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_1019), .B(n_1058), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1051), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1051), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1047), .B(n_1060), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1047), .B(n_1060), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1063), .B(n_1031), .Y(n_1118) );
OR2x2_ASAP7_75t_L g1119 ( .A(n_1058), .B(n_1075), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1070), .B(n_1024), .Y(n_1120) );
INVx1_ASAP7_75t_SL g1121 ( .A(n_1081), .Y(n_1121) );
INVx2_ASAP7_75t_L g1122 ( .A(n_1040), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1052), .B(n_1056), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1052), .B(n_1056), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1046), .B(n_1050), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1046), .B(n_1050), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1046), .B(n_1050), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1057), .B(n_1066), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1129 ( .A(n_1064), .Y(n_1129) );
BUFx3_ASAP7_75t_L g1130 ( .A(n_1022), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1066), .B(n_1037), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1037), .B(n_1065), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_1073), .A2(n_1075), .B1(n_1059), .B2(n_1027), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1029), .B(n_1048), .Y(n_1134) );
BUFx3_ASAP7_75t_L g1135 ( .A(n_1022), .Y(n_1135) );
INVx4_ASAP7_75t_L g1136 ( .A(n_1027), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1046), .B(n_1049), .Y(n_1137) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_1064), .B(n_1088), .Y(n_1138) );
OR2x2_ASAP7_75t_L g1139 ( .A(n_1043), .B(n_1010), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1053), .B(n_1043), .Y(n_1140) );
OR2x2_ASAP7_75t_L g1141 ( .A(n_1016), .B(n_1081), .Y(n_1141) );
INVxp67_ASAP7_75t_SL g1142 ( .A(n_1090), .Y(n_1142) );
INVx1_ASAP7_75t_SL g1143 ( .A(n_1078), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1102), .B(n_1045), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1134), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_1131), .B(n_1054), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_1139), .B(n_1119), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1134), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_1131), .B(n_1068), .Y(n_1149) );
AND2x4_ASAP7_75t_L g1150 ( .A(n_1094), .B(n_1074), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1099), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1099), .Y(n_1152) );
INVx1_ASAP7_75t_SL g1153 ( .A(n_1116), .Y(n_1153) );
AND2x4_ASAP7_75t_L g1154 ( .A(n_1094), .B(n_1074), .Y(n_1154) );
HB1xp67_ASAP7_75t_L g1155 ( .A(n_1141), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1102), .B(n_1045), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1093), .B(n_1068), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1103), .Y(n_1158) );
INVxp67_ASAP7_75t_L g1159 ( .A(n_1141), .Y(n_1159) );
AND2x4_ASAP7_75t_SL g1160 ( .A(n_1136), .B(n_1027), .Y(n_1160) );
INVx4_ASAP7_75t_L g1161 ( .A(n_1100), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1106), .B(n_1045), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1103), .Y(n_1163) );
NAND2xp5_ASAP7_75t_SL g1164 ( .A(n_1121), .B(n_1084), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1106), .B(n_1045), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1108), .B(n_1089), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1108), .B(n_1137), .Y(n_1167) );
HB1xp67_ASAP7_75t_L g1168 ( .A(n_1143), .Y(n_1168) );
INVx1_ASAP7_75t_SL g1169 ( .A(n_1116), .Y(n_1169) );
NOR2xp33_ASAP7_75t_L g1170 ( .A(n_1128), .B(n_1079), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1137), .B(n_1089), .Y(n_1171) );
INVx1_ASAP7_75t_SL g1172 ( .A(n_1117), .Y(n_1172) );
AOI22xp5_ASAP7_75t_L g1173 ( .A1(n_1110), .A2(n_1025), .B1(n_1027), .B2(n_1059), .Y(n_1173) );
INVx2_ASAP7_75t_L g1174 ( .A(n_1122), .Y(n_1174) );
NOR4xp25_ASAP7_75t_SL g1175 ( .A(n_1098), .B(n_1061), .C(n_1080), .D(n_1076), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1109), .Y(n_1176) );
NAND4xp25_ASAP7_75t_L g1177 ( .A(n_1133), .B(n_1085), .C(n_1072), .D(n_1077), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1095), .B(n_1089), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1095), .B(n_1071), .Y(n_1179) );
AND2x4_ASAP7_75t_L g1180 ( .A(n_1094), .B(n_1076), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1113), .B(n_1018), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1096), .B(n_1039), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_1113), .B(n_1018), .Y(n_1183) );
INVx3_ASAP7_75t_L g1184 ( .A(n_1138), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1096), .B(n_1039), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1140), .B(n_1018), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1097), .B(n_1039), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1117), .B(n_1026), .Y(n_1188) );
INVx1_ASAP7_75t_SL g1189 ( .A(n_1132), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1094), .B(n_1039), .Y(n_1190) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1147), .B(n_1114), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1176), .B(n_1128), .Y(n_1192) );
NOR2x1_ASAP7_75t_L g1193 ( .A(n_1161), .B(n_1038), .Y(n_1193) );
INVx1_ASAP7_75t_SL g1194 ( .A(n_1153), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1147), .B(n_1114), .Y(n_1195) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1174), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1151), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1189), .B(n_1115), .Y(n_1198) );
INVx1_ASAP7_75t_SL g1199 ( .A(n_1169), .Y(n_1199) );
INVx3_ASAP7_75t_SL g1200 ( .A(n_1161), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1182), .B(n_1125), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1155), .B(n_1109), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1172), .B(n_1111), .Y(n_1203) );
OR2x2_ASAP7_75t_L g1204 ( .A(n_1178), .B(n_1115), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1151), .Y(n_1205) );
AND2x4_ASAP7_75t_L g1206 ( .A(n_1150), .B(n_1104), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1145), .B(n_1111), .Y(n_1207) );
HB1xp67_ASAP7_75t_L g1208 ( .A(n_1168), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1178), .B(n_1098), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1182), .B(n_1125), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1148), .B(n_1101), .Y(n_1211) );
HB1xp67_ASAP7_75t_L g1212 ( .A(n_1159), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1185), .B(n_1125), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1152), .Y(n_1214) );
INVx2_ASAP7_75t_L g1215 ( .A(n_1174), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1167), .B(n_1101), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1152), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1185), .B(n_1126), .Y(n_1218) );
INVx1_ASAP7_75t_SL g1219 ( .A(n_1149), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1187), .B(n_1126), .Y(n_1220) );
INVx2_ASAP7_75t_SL g1221 ( .A(n_1160), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1158), .Y(n_1222) );
OR2x2_ASAP7_75t_L g1223 ( .A(n_1181), .B(n_1142), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1224 ( .A(n_1181), .B(n_1142), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1187), .B(n_1126), .Y(n_1225) );
INVx1_ASAP7_75t_SL g1226 ( .A(n_1157), .Y(n_1226) );
OR2x2_ASAP7_75t_L g1227 ( .A(n_1183), .B(n_1107), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1163), .Y(n_1228) );
OR2x2_ASAP7_75t_L g1229 ( .A(n_1183), .B(n_1107), .Y(n_1229) );
NAND2x1p5_ASAP7_75t_L g1230 ( .A(n_1161), .B(n_1136), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1170), .B(n_1105), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1144), .B(n_1127), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1197), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1232), .B(n_1144), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1232), .B(n_1156), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1197), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1231), .B(n_1171), .Y(n_1237) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1196), .Y(n_1238) );
AOI22xp5_ASAP7_75t_L g1239 ( .A1(n_1193), .A2(n_1173), .B1(n_1110), .B2(n_1177), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1216), .B(n_1171), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1205), .Y(n_1241) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1196), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1205), .Y(n_1243) );
AND2x4_ASAP7_75t_L g1244 ( .A(n_1206), .B(n_1184), .Y(n_1244) );
AOI22xp33_ASAP7_75t_SL g1245 ( .A1(n_1221), .A2(n_1160), .B1(n_1136), .B2(n_1130), .Y(n_1245) );
INVx2_ASAP7_75t_L g1246 ( .A(n_1215), .Y(n_1246) );
HB1xp67_ASAP7_75t_L g1247 ( .A(n_1194), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1208), .B(n_1162), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1201), .B(n_1156), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1201), .B(n_1162), .Y(n_1250) );
OAI22xp33_ASAP7_75t_L g1251 ( .A1(n_1200), .A2(n_1136), .B1(n_1100), .B2(n_1059), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1214), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1210), .B(n_1165), .Y(n_1253) );
NOR2x1_ASAP7_75t_L g1254 ( .A(n_1223), .B(n_1164), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1210), .B(n_1165), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1214), .Y(n_1256) );
AND2x4_ASAP7_75t_L g1257 ( .A(n_1206), .B(n_1184), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1209), .B(n_1186), .Y(n_1258) );
AOI22xp5_ASAP7_75t_L g1259 ( .A1(n_1219), .A2(n_1120), .B1(n_1059), .B2(n_1179), .Y(n_1259) );
NOR2xp33_ASAP7_75t_L g1260 ( .A(n_1226), .B(n_1146), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1213), .B(n_1166), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1213), .B(n_1166), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1217), .Y(n_1263) );
AOI21xp33_ASAP7_75t_SL g1264 ( .A1(n_1251), .A2(n_1200), .B(n_1230), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1233), .Y(n_1265) );
XNOR2xp5_ASAP7_75t_L g1266 ( .A(n_1239), .B(n_1030), .Y(n_1266) );
NAND2x1_ASAP7_75t_L g1267 ( .A(n_1254), .B(n_1206), .Y(n_1267) );
INVx1_ASAP7_75t_SL g1268 ( .A(n_1247), .Y(n_1268) );
OR2x2_ASAP7_75t_L g1269 ( .A(n_1258), .B(n_1223), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1233), .Y(n_1270) );
O2A1O1Ixp33_ASAP7_75t_L g1271 ( .A1(n_1260), .A2(n_1120), .B(n_1212), .C(n_1044), .Y(n_1271) );
O2A1O1Ixp33_ASAP7_75t_SL g1272 ( .A1(n_1239), .A2(n_1221), .B(n_1199), .C(n_1035), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1236), .Y(n_1273) );
OAI21xp5_ASAP7_75t_SL g1274 ( .A1(n_1245), .A2(n_1230), .B(n_1084), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1234), .B(n_1218), .Y(n_1275) );
AND2x4_ASAP7_75t_L g1276 ( .A(n_1254), .B(n_1150), .Y(n_1276) );
O2A1O1Ixp5_ASAP7_75t_L g1277 ( .A1(n_1244), .A2(n_1211), .B(n_1202), .C(n_1084), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1234), .B(n_1218), .Y(n_1278) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1236), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1241), .Y(n_1280) );
NOR3xp33_ASAP7_75t_L g1281 ( .A(n_1259), .B(n_1082), .C(n_1083), .Y(n_1281) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_1244), .A2(n_1150), .B1(n_1154), .B2(n_1180), .Y(n_1282) );
INVxp67_ASAP7_75t_SL g1283 ( .A(n_1258), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1241), .Y(n_1284) );
AOI21xp33_ASAP7_75t_SL g1285 ( .A1(n_1266), .A2(n_1230), .B(n_1100), .Y(n_1285) );
OAI211xp5_ASAP7_75t_L g1286 ( .A1(n_1264), .A2(n_1083), .B(n_1175), .C(n_1030), .Y(n_1286) );
AOI221xp5_ASAP7_75t_L g1287 ( .A1(n_1272), .A2(n_1237), .B1(n_1248), .B2(n_1240), .C(n_1262), .Y(n_1287) );
AOI221xp5_ASAP7_75t_L g1288 ( .A1(n_1272), .A2(n_1261), .B1(n_1235), .B2(n_1250), .C(n_1249), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1269), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1265), .B(n_1243), .Y(n_1290) );
AOI22xp5_ASAP7_75t_L g1291 ( .A1(n_1266), .A2(n_1257), .B1(n_1191), .B2(n_1195), .Y(n_1291) );
NAND4xp25_ASAP7_75t_L g1292 ( .A(n_1281), .B(n_1112), .C(n_1135), .D(n_1130), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1269), .Y(n_1293) );
OAI322xp33_ASAP7_75t_L g1294 ( .A1(n_1268), .A2(n_1195), .A3(n_1191), .B1(n_1224), .B2(n_1255), .C1(n_1204), .C2(n_1198), .Y(n_1294) );
NOR2xp33_ASAP7_75t_L g1295 ( .A(n_1271), .B(n_1249), .Y(n_1295) );
AOI322xp5_ASAP7_75t_L g1296 ( .A1(n_1283), .A2(n_1250), .A3(n_1253), .B1(n_1225), .B2(n_1220), .C1(n_1257), .C2(n_1203), .Y(n_1296) );
OAI21xp5_ASAP7_75t_SL g1297 ( .A1(n_1285), .A2(n_1274), .B(n_1276), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1290), .Y(n_1298) );
NAND3xp33_ASAP7_75t_L g1299 ( .A(n_1287), .B(n_1277), .C(n_1267), .Y(n_1299) );
AOI322xp5_ASAP7_75t_L g1300 ( .A1(n_1295), .A2(n_1275), .A3(n_1278), .B1(n_1282), .B2(n_1253), .C1(n_1276), .C2(n_1225), .Y(n_1300) );
AND3x1_ASAP7_75t_L g1301 ( .A(n_1288), .B(n_1278), .C(n_1041), .Y(n_1301) );
AOI211xp5_ASAP7_75t_SL g1302 ( .A1(n_1286), .A2(n_1276), .B(n_1062), .C(n_1078), .Y(n_1302) );
OAI211xp5_ASAP7_75t_SL g1303 ( .A1(n_1296), .A2(n_1284), .B(n_1280), .C(n_1270), .Y(n_1303) );
AND4x1_ASAP7_75t_L g1304 ( .A(n_1291), .B(n_1083), .C(n_1273), .D(n_1279), .Y(n_1304) );
AOI222xp33_ASAP7_75t_L g1305 ( .A1(n_1289), .A2(n_1263), .B1(n_1256), .B2(n_1243), .C1(n_1252), .C2(n_1192), .Y(n_1305) );
AOI221xp5_ASAP7_75t_L g1306 ( .A1(n_1303), .A2(n_1294), .B1(n_1293), .B2(n_1290), .C(n_1292), .Y(n_1306) );
AOI22xp5_ASAP7_75t_L g1307 ( .A1(n_1299), .A2(n_1263), .B1(n_1256), .B2(n_1252), .Y(n_1307) );
NAND4xp25_ASAP7_75t_SL g1308 ( .A(n_1300), .B(n_1198), .C(n_1204), .D(n_1188), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_1301), .B(n_1190), .Y(n_1309) );
NAND4xp25_ASAP7_75t_SL g1310 ( .A(n_1305), .B(n_1207), .C(n_1229), .D(n_1227), .Y(n_1310) );
NAND2x1p5_ASAP7_75t_L g1311 ( .A(n_1304), .B(n_1041), .Y(n_1311) );
NAND4xp25_ASAP7_75t_L g1312 ( .A(n_1307), .B(n_1302), .C(n_1297), .D(n_1298), .Y(n_1312) );
NOR5xp2_ASAP7_75t_L g1313 ( .A(n_1308), .B(n_1298), .C(n_1129), .D(n_1217), .E(n_1222), .Y(n_1313) );
NAND2x1p5_ASAP7_75t_L g1314 ( .A(n_1309), .B(n_1087), .Y(n_1314) );
NOR3xp33_ASAP7_75t_SL g1315 ( .A(n_1310), .B(n_1087), .C(n_1118), .Y(n_1315) );
NOR2xp67_ASAP7_75t_L g1316 ( .A(n_1312), .B(n_1306), .Y(n_1316) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1314), .B(n_1311), .Y(n_1317) );
AO21x2_ASAP7_75t_L g1318 ( .A1(n_1315), .A2(n_1124), .B(n_1123), .Y(n_1318) );
AOI21xp33_ASAP7_75t_SL g1319 ( .A1(n_1317), .A2(n_1313), .B(n_1072), .Y(n_1319) );
OAI22xp5_ASAP7_75t_L g1320 ( .A1(n_1316), .A2(n_1135), .B1(n_1112), .B2(n_1227), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1319), .B(n_1318), .Y(n_1321) );
AOI211xp5_ASAP7_75t_L g1322 ( .A1(n_1320), .A2(n_1123), .B(n_1124), .C(n_1118), .Y(n_1322) );
XOR2xp5_ASAP7_75t_L g1323 ( .A(n_1321), .B(n_1229), .Y(n_1323) );
AOI221xp5_ASAP7_75t_L g1324 ( .A1(n_1322), .A2(n_1228), .B1(n_1246), .B2(n_1242), .C(n_1238), .Y(n_1324) );
OAI21xp5_ASAP7_75t_L g1325 ( .A1(n_1323), .A2(n_1091), .B(n_1017), .Y(n_1325) );
OAI21xp5_ASAP7_75t_L g1326 ( .A1(n_1324), .A2(n_1091), .B(n_1017), .Y(n_1326) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1325), .Y(n_1327) );
AOI21xp5_ASAP7_75t_L g1328 ( .A1(n_1327), .A2(n_1326), .B(n_1017), .Y(n_1328) );
endmodule