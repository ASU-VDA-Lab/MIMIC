module fake_netlist_6_1635_n_1154 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1154);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1154;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_465;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_161;
wire n_208;
wire n_462;
wire n_1033;
wire n_1052;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_168;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_840;
wire n_392;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_180;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1099;
wire n_1101;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_181;
wire n_1127;
wire n_182;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_963;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_872;
wire n_1139;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_901;
wire n_923;
wire n_504;
wire n_1078;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_167;
wire n_758;
wire n_174;
wire n_516;
wire n_720;
wire n_631;
wire n_525;
wire n_842;
wire n_1116;
wire n_611;
wire n_943;
wire n_156;
wire n_491;
wire n_843;
wire n_772;
wire n_656;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_343;
wire n_886;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_870;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_163;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_924;
wire n_475;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_936;
wire n_184;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_731;
wire n_570;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_159;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_973;
wire n_346;
wire n_1053;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_1153;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_612;
wire n_453;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_165;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_177;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_170;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_664;
wire n_171;
wire n_949;
wire n_678;
wire n_192;
wire n_169;
wire n_1007;
wire n_649;
wire n_855;
wire n_283;

INVx2_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_84),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_64),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_7),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_146),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_94),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_45),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_93),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_90),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_23),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_17),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_74),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_9),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_65),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_75),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_109),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_1),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_117),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_80),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_5),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_24),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_6),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_124),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_25),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_151),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_29),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_9),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_97),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_143),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_148),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_141),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_100),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_34),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_129),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_20),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_88),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_24),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_137),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_140),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_102),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_101),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_10),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_180),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_184),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_185),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_191),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_156),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_196),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_186),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_155),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_158),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_167),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_159),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_161),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_163),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_164),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_195),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_175),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_179),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_215),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_223),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_213),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_226),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_227),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_208),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_229),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_208),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_232),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_222),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_230),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_216),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_224),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_230),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_209),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_209),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_210),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_211),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_211),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_212),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_212),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_218),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_234),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_236),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_217),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_228),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_217),
.B(n_160),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_222),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_222),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_222),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_221),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_221),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_215),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_213),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_277),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_238),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_282),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_257),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_288),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

INVxp33_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_242),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_258),
.Y(n_300)
);

INVxp33_ASAP7_75t_SL g301 ( 
.A(n_266),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_263),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_249),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_256),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_253),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_284),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_244),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_262),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_263),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_248),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_285),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

INVxp33_ASAP7_75t_SL g317 ( 
.A(n_268),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_251),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_259),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_261),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_279),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_262),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_262),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_262),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_264),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_246),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_245),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_267),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_239),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_269),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_270),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_274),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_273),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_276),
.Y(n_336)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_265),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_328),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_255),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_289),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_294),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_306),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_291),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_312),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_292),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_335),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_328),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_313),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_336),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_331),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_298),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_325),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_307),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_R g358 ( 
.A(n_289),
.B(n_283),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_329),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_323),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_322),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_322),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_293),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_304),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_314),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_316),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_320),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_303),
.B(n_247),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_309),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_335),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_329),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_302),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_313),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_308),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_321),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_304),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_308),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_300),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_301),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_378),
.Y(n_382)
);

NAND2xp33_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_265),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_377),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_338),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_333),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_265),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_355),
.B(n_333),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_342),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_340),
.A2(n_332),
.B1(n_330),
.B2(n_334),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_339),
.B(n_301),
.Y(n_391)
);

AND2x6_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_330),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_365),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_367),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_368),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_352),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_364),
.Y(n_398)
);

BUFx8_ASAP7_75t_L g399 ( 
.A(n_372),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_356),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_352),
.Y(n_402)
);

OA21x2_ASAP7_75t_L g403 ( 
.A1(n_375),
.A2(n_305),
.B(n_295),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_351),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_332),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_350),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_354),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_359),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_348),
.B(n_273),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_381),
.Y(n_412)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_381),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_343),
.B(n_337),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_344),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_380),
.Y(n_418)
);

BUFx8_ASAP7_75t_L g419 ( 
.A(n_345),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_345),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_361),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_341),
.B(n_250),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_361),
.B(n_252),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_362),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_358),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_346),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_362),
.A2(n_272),
.B1(n_193),
.B2(n_206),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_376),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_376),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_379),
.B(n_254),
.Y(n_431)
);

OA21x2_ASAP7_75t_L g432 ( 
.A1(n_374),
.A2(n_295),
.B(n_324),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_379),
.A2(n_245),
.B1(n_287),
.B2(n_317),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_346),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_360),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_374),
.A2(n_326),
.B(n_299),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_360),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_378),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_370),
.B(n_265),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_370),
.B(n_271),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_378),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_378),
.A2(n_299),
.B(n_310),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_338),
.B(n_271),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_352),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_378),
.Y(n_445)
);

CKINVDCx11_ASAP7_75t_R g446 ( 
.A(n_345),
.Y(n_446)
);

OA22x2_ASAP7_75t_SL g447 ( 
.A1(n_375),
.A2(n_275),
.B1(n_186),
.B2(n_154),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_378),
.Y(n_448)
);

OAI22x1_ASAP7_75t_SL g449 ( 
.A1(n_341),
.A2(n_283),
.B1(n_317),
.B2(n_278),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_338),
.B(n_271),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_378),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_338),
.B(n_271),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_352),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_370),
.B(n_172),
.Y(n_454)
);

BUFx8_ASAP7_75t_L g455 ( 
.A(n_342),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_340),
.B(n_315),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_352),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_342),
.Y(n_458)
);

INVx5_ASAP7_75t_L g459 ( 
.A(n_372),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_352),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_338),
.B(n_327),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_370),
.A2(n_182),
.B1(n_192),
.B2(n_203),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_370),
.B(n_200),
.Y(n_463)
);

BUFx8_ASAP7_75t_SL g464 ( 
.A(n_345),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_378),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_378),
.Y(n_466)
);

OAI22x1_ASAP7_75t_L g467 ( 
.A1(n_341),
.A2(n_202),
.B1(n_205),
.B2(n_198),
.Y(n_467)
);

OA21x2_ASAP7_75t_L g468 ( 
.A1(n_378),
.A2(n_169),
.B(n_165),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_171),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_397),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_174),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_384),
.B(n_204),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_393),
.B(n_30),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_384),
.B(n_162),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_401),
.B(n_176),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_382),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_464),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_385),
.B(n_162),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_401),
.B(n_177),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_397),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_393),
.B(n_31),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_385),
.B(n_162),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_418),
.B(n_178),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_382),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_394),
.B(n_183),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_394),
.B(n_395),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_458),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_438),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_438),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_445),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_403),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_404),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_445),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_442),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_395),
.B(n_183),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_396),
.B(n_32),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_456),
.B(n_181),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_456),
.B(n_187),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_428),
.B(n_404),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_418),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_398),
.B(n_189),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_441),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_396),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_400),
.B(n_33),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_400),
.B(n_35),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_448),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_454),
.B(n_190),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_389),
.Y(n_508)
);

INVx6_ASAP7_75t_L g509 ( 
.A(n_397),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_397),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_451),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_386),
.B(n_183),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_466),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_477),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_500),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_500),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_R g517 ( 
.A(n_510),
.B(n_420),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_R g518 ( 
.A(n_510),
.B(n_420),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_493),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_492),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_487),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_502),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_508),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_499),
.A2(n_425),
.B1(n_429),
.B2(n_421),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_510),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_470),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_493),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_486),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_502),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_470),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_470),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_497),
.B(n_422),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_470),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_470),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_R g535 ( 
.A(n_480),
.B(n_426),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_509),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_480),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_509),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_480),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_480),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_486),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_480),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_509),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_509),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_476),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_483),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_506),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_506),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_R g549 ( 
.A(n_502),
.B(n_391),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_R g550 ( 
.A(n_502),
.B(n_446),
.Y(n_550)
);

INVxp33_ASAP7_75t_L g551 ( 
.A(n_483),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_514),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_545),
.Y(n_553)
);

INVxp33_ASAP7_75t_L g554 ( 
.A(n_517),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_548),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_551),
.B(n_532),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_545),
.Y(n_557)
);

BUFx6f_ASAP7_75t_SL g558 ( 
.A(n_528),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_520),
.B(n_498),
.C(n_462),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_541),
.B(n_424),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_519),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_540),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_519),
.Y(n_563)
);

AND3x2_ASAP7_75t_L g564 ( 
.A(n_537),
.B(n_417),
.C(n_427),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_527),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_527),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_521),
.B(n_435),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_524),
.B(n_496),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_523),
.Y(n_569)
);

NOR2x1p5_ASAP7_75t_L g570 ( 
.A(n_514),
.B(n_408),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_515),
.B(n_437),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_515),
.B(n_512),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_522),
.Y(n_573)
);

OAI22xp33_ASAP7_75t_L g574 ( 
.A1(n_546),
.A2(n_511),
.B1(n_513),
.B2(n_390),
.Y(n_574)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_522),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_516),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_516),
.B(n_417),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_549),
.B(n_410),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_518),
.A2(n_467),
.B1(n_478),
.B2(n_474),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_525),
.B(n_512),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_542),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_522),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_529),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_550),
.A2(n_478),
.B1(n_482),
.B2(n_474),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_SL g585 ( 
.A(n_535),
.B(n_406),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_544),
.B(n_482),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_540),
.B(n_496),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_529),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_536),
.A2(n_495),
.B1(n_485),
.B2(n_503),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_544),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_526),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_530),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_531),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_533),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_534),
.Y(n_595)
);

AOI21x1_ASAP7_75t_L g596 ( 
.A1(n_539),
.A2(n_494),
.B(n_491),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_538),
.B(n_485),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_543),
.Y(n_598)
);

BUFx6f_ASAP7_75t_SL g599 ( 
.A(n_547),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_519),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_514),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_519),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_540),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_520),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_519),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_547),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_532),
.A2(n_433),
.B1(n_431),
.B2(n_461),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_551),
.B(n_427),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_540),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_519),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_532),
.B(n_496),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_532),
.A2(n_495),
.B1(n_503),
.B2(n_463),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_532),
.B(n_496),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_523),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_514),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_532),
.B(n_504),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_520),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_551),
.B(n_434),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_532),
.B(n_416),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_536),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_540),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_545),
.Y(n_622)
);

BUFx4f_ASAP7_75t_L g623 ( 
.A(n_528),
.Y(n_623)
);

AND3x1_ASAP7_75t_L g624 ( 
.A(n_532),
.B(n_408),
.C(n_423),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_551),
.B(n_423),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_540),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_547),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_547),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_522),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_556),
.B(n_432),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_592),
.B(n_444),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_595),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_555),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_620),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_574),
.B(n_432),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_595),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_592),
.B(n_444),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_606),
.Y(n_638)
);

INVx4_ASAP7_75t_SL g639 ( 
.A(n_599),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_591),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_594),
.B(n_444),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_562),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_556),
.B(n_406),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_588),
.B(n_504),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_604),
.B(n_464),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_553),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_591),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_622),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_574),
.B(n_432),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_569),
.B(n_446),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_597),
.B(n_472),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_562),
.Y(n_652)
);

NAND3xp33_ASAP7_75t_L g653 ( 
.A(n_612),
.B(n_383),
.C(n_387),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_596),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_557),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_607),
.B(n_406),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_620),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_562),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_579),
.A2(n_388),
.B1(n_386),
.B2(n_443),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_572),
.B(n_590),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_594),
.B(n_444),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_627),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_611),
.B(n_476),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_591),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_591),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_568),
.A2(n_513),
.B1(n_511),
.B2(n_505),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_628),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_563),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_581),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_617),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_562),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_611),
.B(n_484),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_613),
.B(n_484),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_578),
.B(n_554),
.Y(n_674)
);

INVxp33_ASAP7_75t_L g675 ( 
.A(n_618),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_608),
.Y(n_676)
);

AND2x6_ASAP7_75t_L g677 ( 
.A(n_629),
.B(n_504),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_584),
.B(n_406),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_603),
.B(n_453),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_584),
.A2(n_449),
.B1(n_430),
.B2(n_383),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_563),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_SL g682 ( 
.A(n_621),
.B(n_413),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_613),
.B(n_488),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_603),
.B(n_453),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_616),
.B(n_488),
.Y(n_685)
);

NOR2x1p5_ASAP7_75t_L g686 ( 
.A(n_586),
.B(n_430),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_565),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_593),
.B(n_472),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_552),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_616),
.B(n_489),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_619),
.B(n_489),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_566),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_624),
.B(n_453),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_615),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_598),
.B(n_608),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_561),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_612),
.B(n_490),
.Y(n_697)
);

INVxp67_ASAP7_75t_SL g698 ( 
.A(n_600),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_602),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_585),
.B(n_409),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_580),
.B(n_402),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_605),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_603),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_614),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_560),
.B(n_402),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_623),
.B(n_453),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_603),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_571),
.B(n_407),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_676),
.B(n_625),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_633),
.Y(n_710)
);

INVx4_ASAP7_75t_SL g711 ( 
.A(n_640),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_676),
.B(n_618),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_647),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_638),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_675),
.B(n_576),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_667),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_662),
.Y(n_717)
);

INVx5_ASAP7_75t_L g718 ( 
.A(n_640),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_669),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_632),
.Y(n_720)
);

BUFx4_ASAP7_75t_L g721 ( 
.A(n_689),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_696),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_630),
.B(n_567),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_656),
.A2(n_568),
.B1(n_674),
.B2(n_678),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_630),
.B(n_567),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_655),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_682),
.B(n_623),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_698),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_640),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_698),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_639),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_695),
.B(n_589),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_699),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_705),
.B(n_589),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_691),
.B(n_577),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_680),
.A2(n_579),
.B1(n_558),
.B2(n_599),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_664),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_646),
.Y(n_738)
);

NAND2x1p5_ASAP7_75t_L g739 ( 
.A(n_647),
.B(n_587),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_654),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_703),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_660),
.B(n_577),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_648),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_682),
.B(n_609),
.Y(n_744)
);

OA22x2_ASAP7_75t_L g745 ( 
.A1(n_643),
.A2(n_564),
.B1(n_657),
.B2(n_706),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_668),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_681),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_687),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_654),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_691),
.B(n_636),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_664),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_703),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_704),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_663),
.B(n_573),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_651),
.B(n_609),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_692),
.Y(n_756)
);

INVx4_ASAP7_75t_SL g757 ( 
.A(n_664),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_659),
.A2(n_558),
.B1(n_559),
.B2(n_621),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_642),
.B(n_609),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_634),
.B(n_601),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_663),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_642),
.B(n_609),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_702),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_672),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_652),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_670),
.B(n_419),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_703),
.B(n_504),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_672),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_652),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_658),
.B(n_626),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_673),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_673),
.B(n_573),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_683),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_665),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_658),
.B(n_671),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_701),
.B(n_626),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_683),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_685),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_721),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_719),
.Y(n_780)
);

BUFx5_ASAP7_75t_L g781 ( 
.A(n_767),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_731),
.B(n_694),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_731),
.B(n_639),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_720),
.B(n_686),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_712),
.B(n_650),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_758),
.A2(n_700),
.B1(n_666),
.B2(n_653),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_709),
.B(n_708),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_761),
.B(n_635),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_L g789 ( 
.A(n_736),
.B(n_659),
.C(n_649),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_723),
.B(n_645),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_745),
.B(n_639),
.Y(n_791)
);

AND2x6_ASAP7_75t_SL g792 ( 
.A(n_766),
.B(n_419),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_740),
.B(n_635),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_714),
.Y(n_794)
);

OAI22xp33_ASAP7_75t_L g795 ( 
.A1(n_725),
.A2(n_649),
.B1(n_653),
.B2(n_666),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_750),
.B(n_685),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_724),
.B(n_665),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_715),
.B(n_665),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_727),
.A2(n_387),
.B1(n_688),
.B2(n_677),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_718),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_753),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_729),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_710),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_749),
.B(n_690),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_734),
.A2(n_677),
.B1(n_587),
.B2(n_693),
.Y(n_805)
);

AO22x1_ASAP7_75t_L g806 ( 
.A1(n_760),
.A2(n_644),
.B1(n_677),
.B2(n_455),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_716),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_732),
.A2(n_166),
.B1(n_677),
.B2(n_637),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_722),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_717),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_735),
.B(n_631),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_776),
.B(n_671),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_726),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_756),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_729),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_773),
.B(n_777),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_763),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_729),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_777),
.B(n_697),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_733),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_744),
.B(n_697),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_764),
.B(n_707),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_755),
.A2(n_166),
.B1(n_637),
.B2(n_631),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_742),
.B(n_707),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_775),
.B(n_641),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_768),
.B(n_605),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_737),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_775),
.B(n_641),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_771),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_759),
.B(n_661),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_739),
.B(n_661),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_767),
.A2(n_166),
.B1(n_644),
.B2(n_405),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_759),
.B(n_684),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_762),
.B(n_626),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_778),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_713),
.A2(n_505),
.B(n_570),
.C(n_679),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_737),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_728),
.B(n_730),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_746),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_SL g840 ( 
.A(n_718),
.B(n_626),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_754),
.B(n_610),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_737),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_767),
.A2(n_166),
.B1(n_644),
.B2(n_405),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_747),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_762),
.B(n_679),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_770),
.B(n_615),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_770),
.B(n_684),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_748),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_713),
.B(n_409),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_738),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_800),
.B(n_765),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_780),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_779),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_794),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_787),
.B(n_769),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_788),
.B(n_772),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_800),
.B(n_711),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_803),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_824),
.B(n_774),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_838),
.B(n_711),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_796),
.B(n_743),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_791),
.B(n_751),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_829),
.B(n_774),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_835),
.B(n_741),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_807),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_788),
.B(n_741),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_784),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_809),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_789),
.A2(n_752),
.B(n_436),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_810),
.B(n_812),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_801),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_815),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_820),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_816),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_837),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_813),
.B(n_752),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_816),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_814),
.B(n_751),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_785),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_817),
.B(n_718),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_850),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_822),
.B(n_757),
.Y(n_882)
);

INVxp33_ASAP7_75t_L g883 ( 
.A(n_846),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_839),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_821),
.B(n_757),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_789),
.A2(n_767),
.B(n_644),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_838),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_821),
.B(n_582),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_821),
.B(n_582),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_844),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_790),
.B(n_409),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_825),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_811),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_848),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_819),
.B(n_583),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_804),
.Y(n_896)
);

INVxp33_ASAP7_75t_L g897 ( 
.A(n_798),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_886),
.A2(n_786),
.B(n_795),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_883),
.B(n_879),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_857),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_875),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_869),
.A2(n_806),
.B(n_783),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_872),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_887),
.B(n_793),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_856),
.B(n_896),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_862),
.A2(n_836),
.B(n_797),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_897),
.A2(n_782),
.B(n_819),
.Y(n_907)
);

OAI21xp33_ASAP7_75t_L g908 ( 
.A1(n_856),
.A2(n_805),
.B(n_804),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_891),
.A2(n_831),
.B(n_799),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_882),
.A2(n_840),
.B(n_849),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_853),
.A2(n_834),
.B(n_845),
.C(n_826),
.Y(n_911)
);

INVx5_ASAP7_75t_L g912 ( 
.A(n_857),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_860),
.B(n_833),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_857),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_861),
.A2(n_840),
.B(n_808),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_885),
.A2(n_843),
.B(n_832),
.C(n_828),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_866),
.A2(n_841),
.B(n_826),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_855),
.B(n_847),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_885),
.A2(n_830),
.B(n_823),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_860),
.B(n_802),
.Y(n_920)
);

AOI21x1_ASAP7_75t_L g921 ( 
.A1(n_857),
.A2(n_827),
.B(n_818),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_863),
.A2(n_842),
.B(n_507),
.C(n_469),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_864),
.A2(n_468),
.B(n_575),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_860),
.B(n_781),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_895),
.A2(n_468),
.B(n_471),
.Y(n_925)
);

AO21x1_ASAP7_75t_L g926 ( 
.A1(n_860),
.A2(n_413),
.B(n_505),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_893),
.B(n_781),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_872),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_888),
.B(n_781),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_852),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_889),
.B(n_781),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_870),
.B(n_781),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_889),
.B(n_792),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_867),
.A2(n_409),
.B(n_411),
.C(n_412),
.Y(n_934)
);

BUFx4f_ASAP7_75t_L g935 ( 
.A(n_875),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_865),
.A2(n_873),
.B(n_890),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_876),
.B(n_166),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_872),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_859),
.B(n_411),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_874),
.A2(n_877),
.B(n_851),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_875),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_871),
.B(n_411),
.Y(n_942)
);

AOI21xp33_ASAP7_75t_L g943 ( 
.A1(n_851),
.A2(n_399),
.B(n_455),
.Y(n_943)
);

OR2x2_ASAP7_75t_SL g944 ( 
.A(n_875),
.B(n_411),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_898),
.A2(n_873),
.B(n_851),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_SL g946 ( 
.A(n_914),
.B(n_875),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_908),
.B(n_868),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_912),
.B(n_851),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_914),
.B(n_859),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_901),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_933),
.B(n_892),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_899),
.B(n_868),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_938),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_917),
.B(n_878),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_913),
.B(n_878),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_912),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_906),
.B(n_881),
.Y(n_957)
);

NAND2x1p5_ASAP7_75t_L g958 ( 
.A(n_912),
.B(n_858),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_935),
.B(n_852),
.Y(n_959)
);

AOI21x1_ASAP7_75t_L g960 ( 
.A1(n_937),
.A2(n_894),
.B(n_884),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_911),
.B(n_881),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_901),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_935),
.B(n_880),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_SL g964 ( 
.A1(n_934),
.A2(n_854),
.B(n_858),
.C(n_894),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_964),
.A2(n_957),
.B(n_961),
.C(n_948),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_945),
.A2(n_902),
.B1(n_900),
.B2(n_926),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_951),
.A2(n_924),
.B(n_907),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_953),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_956),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_951),
.A2(n_919),
.B(n_943),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_947),
.A2(n_909),
.B(n_923),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_952),
.B(n_905),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_959),
.A2(n_915),
.B(n_910),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_952),
.B(n_942),
.Y(n_974)
);

NAND3xp33_ASAP7_75t_SL g975 ( 
.A(n_946),
.B(n_916),
.C(n_941),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_954),
.A2(n_936),
.B(n_940),
.C(n_925),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_950),
.B(n_941),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_959),
.A2(n_927),
.B(n_922),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_956),
.B(n_901),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_962),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_963),
.A2(n_920),
.B1(n_928),
.B2(n_929),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_949),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_955),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_958),
.B(n_920),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_958),
.A2(n_931),
.B(n_904),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_SL g986 ( 
.A(n_960),
.B(n_903),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_947),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_956),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_956),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_984),
.B(n_921),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_966),
.A2(n_973),
.B1(n_981),
.B2(n_967),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_989),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_968),
.B(n_939),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_987),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_983),
.B(n_932),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_988),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_988),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_991),
.A2(n_975),
.B(n_970),
.Y(n_998)
);

AND2x6_ASAP7_75t_L g999 ( 
.A(n_997),
.B(n_412),
.Y(n_999)
);

O2A1O1Ixp5_ASAP7_75t_SL g1000 ( 
.A1(n_992),
.A2(n_969),
.B(n_979),
.C(n_977),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_998),
.A2(n_965),
.B(n_996),
.C(n_976),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_999),
.B(n_982),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_1002),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_1001),
.A2(n_1000),
.B(n_971),
.Y(n_1004)
);

AO21x2_ASAP7_75t_L g1005 ( 
.A1(n_1004),
.A2(n_994),
.B(n_990),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_1003),
.Y(n_1006)
);

AO22x2_ASAP7_75t_L g1007 ( 
.A1(n_1006),
.A2(n_969),
.B1(n_978),
.B2(n_990),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_SL g1008 ( 
.A1(n_1005),
.A2(n_986),
.B1(n_988),
.B2(n_980),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_1007),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1008),
.Y(n_1010)
);

NOR2xp67_ASAP7_75t_R g1011 ( 
.A(n_1010),
.B(n_412),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1009),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_1012),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_1011),
.A2(n_1005),
.B1(n_980),
.B2(n_995),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1012),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_1013),
.B(n_993),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_1015),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_1014),
.Y(n_1018)
);

OA21x2_ASAP7_75t_L g1019 ( 
.A1(n_1017),
.A2(n_974),
.B(n_993),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1016),
.B(n_980),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_1019),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_1020),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_1021),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_1022),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_1023),
.B(n_1019),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1024),
.B(n_1018),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_1026),
.B(n_972),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_1025),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_1027),
.B(n_412),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1028),
.B(n_985),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_1030),
.B(n_414),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_1029),
.B(n_414),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1030),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_1033),
.B(n_414),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1031),
.B(n_399),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1032),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_SL g1037 ( 
.A1(n_1035),
.A2(n_414),
.B(n_461),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1034),
.B(n_930),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1038),
.B(n_1036),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_1037),
.A2(n_415),
.B(n_416),
.Y(n_1040)
);

NOR2xp67_ASAP7_75t_L g1041 ( 
.A(n_1039),
.B(n_0),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_1040),
.B(n_0),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1041),
.B(n_1),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1042),
.B(n_918),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1043),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1044),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_L g1047 ( 
.A(n_1046),
.B(n_197),
.C(n_443),
.Y(n_1047)
);

NAND2x1_ASAP7_75t_L g1048 ( 
.A(n_1045),
.B(n_450),
.Y(n_1048)
);

OAI21xp33_ASAP7_75t_L g1049 ( 
.A1(n_1047),
.A2(n_452),
.B(n_450),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1048),
.B(n_2),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_1047),
.A2(n_452),
.B(n_388),
.C(n_459),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1050),
.A2(n_1051),
.B1(n_1049),
.B2(n_459),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1050),
.Y(n_1053)
);

AOI221xp5_ASAP7_75t_L g1054 ( 
.A1(n_1050),
.A2(n_457),
.B1(n_460),
.B2(n_501),
.C(n_459),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1053),
.B(n_2),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_1052),
.Y(n_1056)
);

INVxp67_ASAP7_75t_SL g1057 ( 
.A(n_1056),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_1055),
.Y(n_1058)
);

NOR3xp33_ASAP7_75t_L g1059 ( 
.A(n_1057),
.B(n_1054),
.C(n_3),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1058),
.A2(n_459),
.B1(n_457),
.B2(n_460),
.Y(n_1060)
);

NOR2x1_ASAP7_75t_L g1061 ( 
.A(n_1059),
.B(n_457),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1060),
.B(n_457),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1061),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1062),
.Y(n_1064)
);

NOR2x1_ASAP7_75t_L g1065 ( 
.A(n_1063),
.B(n_1064),
.Y(n_1065)
);

OAI211xp5_ASAP7_75t_L g1066 ( 
.A1(n_1064),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1065),
.A2(n_479),
.B(n_475),
.Y(n_1067)
);

OAI211xp5_ASAP7_75t_SL g1068 ( 
.A1(n_1066),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1065),
.A2(n_460),
.B(n_8),
.Y(n_1069)
);

NAND4xp75_ASAP7_75t_L g1070 ( 
.A(n_1067),
.B(n_1069),
.C(n_1068),
.D(n_11),
.Y(n_1070)
);

NAND4xp75_ASAP7_75t_L g1071 ( 
.A(n_1067),
.B(n_8),
.C(n_10),
.D(n_11),
.Y(n_1071)
);

OAI21xp33_ASAP7_75t_L g1072 ( 
.A1(n_1068),
.A2(n_460),
.B(n_12),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_1070),
.A2(n_12),
.B(n_13),
.Y(n_1073)
);

NOR4xp75_ASAP7_75t_L g1074 ( 
.A(n_1072),
.B(n_13),
.C(n_14),
.D(n_15),
.Y(n_1074)
);

AOI211xp5_ASAP7_75t_L g1075 ( 
.A1(n_1073),
.A2(n_1071),
.B(n_15),
.C(n_16),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_L g1076 ( 
.A(n_1074),
.B(n_14),
.C(n_16),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_1075),
.B(n_17),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_L g1078 ( 
.A(n_1076),
.B(n_18),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_SL g1079 ( 
.A1(n_1078),
.A2(n_18),
.B(n_19),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1077),
.Y(n_1080)
);

OAI22x1_ASAP7_75t_SL g1081 ( 
.A1(n_1080),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1079),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1082),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_1081),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1083),
.Y(n_1085)
);

XOR2x2_ASAP7_75t_L g1086 ( 
.A(n_1084),
.B(n_21),
.Y(n_1086)
);

NAND3x1_ASAP7_75t_L g1087 ( 
.A(n_1083),
.B(n_22),
.C(n_23),
.Y(n_1087)
);

NOR2x1_ASAP7_75t_R g1088 ( 
.A(n_1085),
.B(n_22),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_1086),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_1087),
.B(n_26),
.Y(n_1090)
);

NOR3xp33_ASAP7_75t_L g1091 ( 
.A(n_1090),
.B(n_27),
.C(n_28),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1088),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1092),
.B(n_1089),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1091),
.Y(n_1094)
);

AND2x2_ASAP7_75t_SL g1095 ( 
.A(n_1093),
.B(n_28),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_1094),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_SL g1097 ( 
.A(n_1096),
.B(n_447),
.C(n_36),
.Y(n_1097)
);

AND3x1_ASAP7_75t_L g1098 ( 
.A(n_1095),
.B(n_37),
.C(n_38),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1098),
.B(n_39),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1097),
.Y(n_1100)
);

XNOR2xp5_ASAP7_75t_L g1101 ( 
.A(n_1100),
.B(n_40),
.Y(n_1101)
);

AOI221xp5_ASAP7_75t_L g1102 ( 
.A1(n_1099),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.C(n_44),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1101),
.A2(n_405),
.B(n_473),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1102),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_1101),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1105),
.A2(n_944),
.B1(n_481),
.B2(n_473),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_SL g1107 ( 
.A1(n_1104),
.A2(n_481),
.B1(n_473),
.B2(n_48),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1103),
.A2(n_405),
.B1(n_392),
.B2(n_473),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1104),
.A2(n_405),
.B(n_481),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1107),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1108),
.A2(n_1106),
.B1(n_1109),
.B2(n_481),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1108),
.A2(n_505),
.B1(n_465),
.B2(n_49),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1110),
.A2(n_392),
.B1(n_47),
.B2(n_50),
.Y(n_1113)
);

OAI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_1111),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1112),
.A2(n_53),
.B(n_54),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1115),
.A2(n_1114),
.B(n_1113),
.Y(n_1116)
);

AOI221xp5_ASAP7_75t_L g1117 ( 
.A1(n_1115),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.C(n_58),
.Y(n_1117)
);

AOI222xp33_ASAP7_75t_L g1118 ( 
.A1(n_1114),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.C1(n_62),
.C2(n_63),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1115),
.Y(n_1119)
);

AO221x1_ASAP7_75t_L g1120 ( 
.A1(n_1114),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.C(n_69),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_1115),
.B(n_70),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1115),
.A2(n_71),
.B(n_72),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1115),
.B(n_73),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1115),
.A2(n_76),
.B(n_77),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1115),
.A2(n_78),
.B(n_79),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1115),
.A2(n_81),
.B(n_82),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1115),
.B(n_83),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1119),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1116),
.A2(n_85),
.B(n_86),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1121),
.Y(n_1130)
);

INVxp33_ASAP7_75t_SL g1131 ( 
.A(n_1123),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_1127),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1125),
.A2(n_87),
.B1(n_89),
.B2(n_91),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1126),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1120),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1122),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_SL g1137 ( 
.A1(n_1128),
.A2(n_1124),
.B1(n_1118),
.B2(n_1117),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1136),
.Y(n_1138)
);

AOI222xp33_ASAP7_75t_SL g1139 ( 
.A1(n_1135),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.C1(n_98),
.C2(n_99),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1131),
.A2(n_392),
.B1(n_104),
.B2(n_105),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1134),
.A2(n_392),
.B1(n_106),
.B2(n_108),
.Y(n_1141)
);

AOI21xp33_ASAP7_75t_L g1142 ( 
.A1(n_1132),
.A2(n_103),
.B(n_111),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1138),
.A2(n_1137),
.B(n_1130),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1141),
.A2(n_1133),
.B(n_1129),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1139),
.A2(n_1140),
.B(n_1142),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1138),
.A2(n_112),
.B(n_113),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1143),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1147),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1148),
.A2(n_1145),
.B1(n_1144),
.B2(n_1146),
.Y(n_1149)
);

OAI221xp5_ASAP7_75t_R g1150 ( 
.A1(n_1149),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.C(n_121),
.Y(n_1150)
);

AOI221xp5_ASAP7_75t_L g1151 ( 
.A1(n_1150),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.C(n_127),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1151),
.A2(n_128),
.B(n_131),
.Y(n_1152)
);

AOI211xp5_ASAP7_75t_L g1153 ( 
.A1(n_1152),
.A2(n_132),
.B(n_133),
.C(n_134),
.Y(n_1153)
);

AOI211xp5_ASAP7_75t_L g1154 ( 
.A1(n_1153),
.A2(n_135),
.B(n_136),
.C(n_139),
.Y(n_1154)
);


endmodule