module fake_ibex_1486_n_875 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_875);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_875;

wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_698;
wire n_187;
wire n_667;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_723;
wire n_270;
wire n_170;
wire n_383;
wire n_346;
wire n_840;
wire n_561;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_158;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_798;
wire n_832;
wire n_732;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_617;
wire n_496;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_651;
wire n_581;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_729;
wire n_807;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_820;
wire n_805;
wire n_670;
wire n_728;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_202;
wire n_159;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx2_ASAP7_75t_L g157 ( 
.A(n_37),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_14),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_0),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_22),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_48),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_62),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_41),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_80),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_83),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_64),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_33),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_7),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_90),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_104),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_153),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_31),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_88),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_17),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_26),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_50),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_135),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_1),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_128),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_18),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_13),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_109),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_148),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_127),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_69),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_87),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_30),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_14),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_16),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_137),
.Y(n_200)
);

BUFx2_ASAP7_75t_SL g201 ( 
.A(n_3),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_29),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_46),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_96),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_45),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_91),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_75),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_134),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_84),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_55),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_136),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_141),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_58),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_60),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_82),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_L g218 ( 
.A(n_92),
.B(n_11),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_13),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_40),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_73),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_33),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_114),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_100),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_26),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_93),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_156),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_86),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_66),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_76),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_132),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_106),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_120),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_95),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_21),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_43),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_151),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_152),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_107),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_81),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_97),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_117),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_L g244 ( 
.A(n_111),
.B(n_28),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_63),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_35),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_74),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_68),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_130),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_49),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_4),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_32),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_178),
.Y(n_256)
);

AOI22x1_ASAP7_75t_SL g257 ( 
.A1(n_173),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_248),
.Y(n_258)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_175),
.B(n_3),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_174),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_193),
.B(n_6),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_178),
.B(n_7),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

CKINVDCx11_ASAP7_75t_R g268 ( 
.A(n_190),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_8),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_235),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_182),
.B(n_8),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_227),
.B(n_9),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_173),
.B(n_202),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_183),
.B(n_9),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_235),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_183),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_202),
.B(n_10),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g280 ( 
.A(n_186),
.B(n_160),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_222),
.B(n_10),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

BUFx8_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_157),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_163),
.Y(n_288)
);

CKINVDCx11_ASAP7_75t_R g289 ( 
.A(n_190),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_197),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_222),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_291)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_199),
.B(n_12),
.Y(n_292)
);

OA21x2_ASAP7_75t_L g293 ( 
.A1(n_157),
.A2(n_89),
.B(n_150),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g294 ( 
.A(n_167),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_236),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_236),
.B(n_19),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_225),
.B(n_20),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_211),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_246),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_159),
.Y(n_300)
);

AND2x4_ASAP7_75t_L g301 ( 
.A(n_251),
.B(n_23),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_211),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_195),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_188),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_235),
.Y(n_306)
);

OA22x2_ASAP7_75t_SL g307 ( 
.A1(n_195),
.A2(n_238),
.B1(n_212),
.B2(n_221),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g308 ( 
.A1(n_232),
.A2(n_94),
.B(n_149),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_212),
.Y(n_309)
);

INVxp33_ASAP7_75t_SL g310 ( 
.A(n_167),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_237),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_234),
.B(n_24),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_232),
.B(n_25),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_189),
.B(n_27),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_158),
.B(n_27),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_161),
.B(n_164),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_221),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_165),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_201),
.B(n_29),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_166),
.B(n_30),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_198),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_266),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_285),
.B(n_168),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_285),
.B(n_312),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_262),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_292),
.A2(n_219),
.B1(n_249),
.B2(n_247),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

OAI22x1_ASAP7_75t_L g328 ( 
.A1(n_303),
.A2(n_207),
.B1(n_176),
.B2(n_181),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_267),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_258),
.B(n_176),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_312),
.B(n_169),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_315),
.B(n_171),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_258),
.B(n_181),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_253),
.B(n_209),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_300),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_281),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_292),
.A2(n_250),
.B1(n_180),
.B2(n_184),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_281),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_266),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_261),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_261),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_269),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_284),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_315),
.B(n_187),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_275),
.B(n_204),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_R g349 ( 
.A(n_311),
.B(n_294),
.Y(n_349)
);

AND2x6_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_191),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_273),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_273),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_261),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_276),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_255),
.B(n_196),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_261),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_284),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_271),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_316),
.B(n_218),
.Y(n_359)
);

OR2x6_ASAP7_75t_L g360 ( 
.A(n_295),
.B(n_244),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_276),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_310),
.B(n_207),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_271),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_301),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_320),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_310),
.B(n_224),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_271),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_316),
.B(n_318),
.Y(n_368)
);

BUFx10_ASAP7_75t_L g369 ( 
.A(n_311),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_280),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_280),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_318),
.B(n_200),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_277),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_277),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_277),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_254),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_290),
.A2(n_216),
.B1(n_213),
.B2(n_208),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_287),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_286),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_287),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_294),
.B(n_238),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_287),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_279),
.B(n_231),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g384 ( 
.A(n_274),
.B(n_231),
.C(n_203),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_286),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_299),
.A2(n_230),
.B1(n_215),
.B2(n_205),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_288),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_306),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_293),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_306),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_288),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_304),
.B(n_162),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_304),
.Y(n_393)
);

NAND2xp33_ASAP7_75t_SL g394 ( 
.A(n_263),
.B(n_179),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_265),
.B(n_206),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_274),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_298),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_298),
.Y(n_398)
);

AND3x2_ASAP7_75t_L g399 ( 
.A(n_307),
.B(n_170),
.C(n_229),
.Y(n_399)
);

INVx4_ASAP7_75t_SL g400 ( 
.A(n_259),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_256),
.B(n_185),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_306),
.Y(n_402)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_259),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_302),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_302),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_259),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_272),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_254),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_254),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_278),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_254),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_313),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_412),
.B(n_348),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_341),
.A2(n_297),
.B1(n_282),
.B2(n_296),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_348),
.B(n_314),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_391),
.Y(n_416)
);

BUFx6f_ASAP7_75t_SL g417 ( 
.A(n_369),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_336),
.B(n_317),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_341),
.B(n_291),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_404),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_383),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_405),
.Y(n_422)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_350),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_383),
.B(n_192),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_332),
.A2(n_309),
.B1(n_289),
.B2(n_268),
.Y(n_425)
);

BUFx12f_ASAP7_75t_L g426 ( 
.A(n_369),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_330),
.B(n_214),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_334),
.B(n_194),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_332),
.B(n_319),
.Y(n_429)
);

O2A1O1Ixp33_ASAP7_75t_L g430 ( 
.A1(n_322),
.A2(n_321),
.B(n_240),
.C(n_220),
.Y(n_430)
);

O2A1O1Ixp5_ASAP7_75t_L g431 ( 
.A1(n_389),
.A2(n_241),
.B(n_223),
.C(n_226),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_324),
.B(n_264),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_387),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_362),
.B(n_245),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_351),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_361),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_326),
.A2(n_228),
.B1(n_233),
.B2(n_242),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_366),
.B(n_177),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_333),
.B(n_347),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_335),
.B(n_239),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_345),
.B(n_268),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_392),
.B(n_293),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_324),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_333),
.B(n_308),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_364),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_350),
.A2(n_257),
.B1(n_289),
.B2(n_260),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_339),
.A2(n_260),
.B1(n_35),
.B2(n_36),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_401),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_347),
.B(n_260),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_365),
.B(n_260),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_349),
.Y(n_452)
);

OAI22x1_ASAP7_75t_SL g453 ( 
.A1(n_399),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_453)
);

AND2x6_ASAP7_75t_SL g454 ( 
.A(n_360),
.B(n_39),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_396),
.B(n_42),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_395),
.B(n_44),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_L g457 ( 
.A(n_328),
.B(n_47),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_395),
.B(n_51),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_323),
.B(n_52),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_368),
.B(n_331),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_368),
.B(n_331),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_361),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_361),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_323),
.B(n_53),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_370),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_379),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_371),
.B(n_54),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_407),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_350),
.A2(n_352),
.B1(n_354),
.B2(n_389),
.Y(n_469)
);

NAND3xp33_ASAP7_75t_SL g470 ( 
.A(n_381),
.B(n_56),
.C(n_57),
.Y(n_470)
);

OAI221xp5_ASAP7_75t_L g471 ( 
.A1(n_377),
.A2(n_59),
.B1(n_61),
.B2(n_65),
.C(n_67),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_410),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_359),
.B(n_71),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_359),
.B(n_72),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_369),
.B(n_355),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_384),
.B(n_77),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_359),
.B(n_78),
.Y(n_478)
);

NAND2xp33_ASAP7_75t_L g479 ( 
.A(n_350),
.B(n_79),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_350),
.B(n_386),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_372),
.B(n_98),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_394),
.B(n_99),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_397),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_397),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_397),
.B(n_398),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_360),
.A2(n_101),
.B1(n_103),
.B2(n_105),
.Y(n_488)
);

NOR3xp33_ASAP7_75t_L g489 ( 
.A(n_398),
.B(n_108),
.C(n_110),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_398),
.B(n_112),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_419),
.A2(n_328),
.B1(n_360),
.B2(n_357),
.Y(n_491)
);

O2A1O1Ixp33_ASAP7_75t_SL g492 ( 
.A1(n_443),
.A2(n_338),
.B(n_357),
.C(n_346),
.Y(n_492)
);

O2A1O1Ixp33_ASAP7_75t_L g493 ( 
.A1(n_413),
.A2(n_360),
.B(n_337),
.C(n_343),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_426),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_420),
.Y(n_495)
);

A2O1A1Ixp33_ASAP7_75t_L g496 ( 
.A1(n_415),
.A2(n_445),
.B(n_427),
.C(n_440),
.Y(n_496)
);

NOR2xp67_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_113),
.Y(n_497)
);

NOR2x1p5_ASAP7_75t_L g498 ( 
.A(n_418),
.B(n_376),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_421),
.B(n_329),
.Y(n_499)
);

O2A1O1Ixp33_ASAP7_75t_L g500 ( 
.A1(n_430),
.A2(n_325),
.B(n_327),
.C(n_340),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_437),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_462),
.Y(n_502)
);

AND2x4_ASAP7_75t_SL g503 ( 
.A(n_442),
.B(n_411),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_449),
.B(n_376),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_449),
.B(n_411),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_422),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_452),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_463),
.Y(n_508)
);

AND2x2_ASAP7_75t_SL g509 ( 
.A(n_423),
.B(n_409),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_423),
.B(n_408),
.Y(n_510)
);

NAND2x1p5_ASAP7_75t_L g511 ( 
.A(n_485),
.B(n_408),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_444),
.B(n_115),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_436),
.B(n_406),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_417),
.B(n_406),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_468),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_417),
.B(n_374),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_446),
.B(n_403),
.Y(n_517)
);

BUFx4f_ASAP7_75t_L g518 ( 
.A(n_419),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_485),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_471),
.B(n_374),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_475),
.B(n_400),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_429),
.B(n_424),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_432),
.B(n_400),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_472),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_483),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_465),
.B(n_403),
.Y(n_526)
);

A2O1A1Ixp33_ASAP7_75t_L g527 ( 
.A1(n_427),
.A2(n_373),
.B(n_363),
.C(n_390),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_439),
.B(n_118),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_473),
.Y(n_529)
);

AO22x1_ASAP7_75t_L g530 ( 
.A1(n_419),
.A2(n_403),
.B1(n_122),
.B2(n_123),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_457),
.B(n_121),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_469),
.B(n_403),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_431),
.A2(n_373),
.B(n_388),
.Y(n_533)
);

OR2x6_ASAP7_75t_SL g534 ( 
.A(n_425),
.B(n_124),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_481),
.A2(n_367),
.B1(n_388),
.B2(n_382),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_434),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_431),
.A2(n_380),
.B(n_378),
.Y(n_537)
);

AO21x1_ASAP7_75t_L g538 ( 
.A1(n_489),
.A2(n_378),
.B(n_126),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_466),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_414),
.B(n_402),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_488),
.B(n_402),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_460),
.A2(n_353),
.B1(n_344),
.B2(n_342),
.Y(n_542)
);

A2O1A1Ixp33_ASAP7_75t_L g543 ( 
.A1(n_460),
.A2(n_402),
.B(n_353),
.C(n_344),
.Y(n_543)
);

AOI21x1_ASAP7_75t_L g544 ( 
.A1(n_456),
.A2(n_402),
.B(n_353),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_483),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_419),
.A2(n_353),
.B1(n_344),
.B2(n_342),
.Y(n_546)
);

NOR2x1_ASAP7_75t_L g547 ( 
.A(n_435),
.B(n_344),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_458),
.A2(n_375),
.B(n_358),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_486),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_486),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_461),
.B(n_419),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_487),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_482),
.B(n_342),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_482),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_428),
.B(n_342),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_438),
.B(n_133),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_476),
.Y(n_557)
);

A2O1A1Ixp33_ASAP7_75t_L g558 ( 
.A1(n_467),
.A2(n_356),
.B(n_138),
.C(n_140),
.Y(n_558)
);

OA22x2_ASAP7_75t_L g559 ( 
.A1(n_454),
.A2(n_448),
.B1(n_453),
.B2(n_459),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_474),
.B(n_478),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_416),
.Y(n_561)
);

OR2x6_ASAP7_75t_SL g562 ( 
.A(n_441),
.B(n_484),
.Y(n_562)
);

AOI21x1_ASAP7_75t_L g563 ( 
.A1(n_490),
.A2(n_356),
.B(n_142),
.Y(n_563)
);

INVx3_ASAP7_75t_SL g564 ( 
.A(n_464),
.Y(n_564)
);

AND2x4_ASAP7_75t_SL g565 ( 
.A(n_433),
.B(n_480),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_467),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_451),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_455),
.A2(n_479),
.B(n_450),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_477),
.B(n_489),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_549),
.B(n_551),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_519),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_522),
.A2(n_470),
.B1(n_549),
.B2(n_506),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_548),
.A2(n_544),
.B(n_563),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_494),
.Y(n_574)
);

AO32x2_ASAP7_75t_L g575 ( 
.A1(n_542),
.A2(n_535),
.A3(n_567),
.B1(n_529),
.B2(n_538),
.Y(n_575)
);

BUFx12f_ASAP7_75t_L g576 ( 
.A(n_494),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_515),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_511),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_524),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_491),
.A2(n_518),
.B1(n_554),
.B2(n_559),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_499),
.B(n_498),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_534),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_523),
.B(n_536),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_552),
.Y(n_584)
);

OA21x2_ASAP7_75t_L g585 ( 
.A1(n_543),
.A2(n_537),
.B(n_533),
.Y(n_585)
);

NAND3x1_ASAP7_75t_L g586 ( 
.A(n_559),
.B(n_518),
.C(n_562),
.Y(n_586)
);

O2A1O1Ixp5_ASAP7_75t_SL g587 ( 
.A1(n_540),
.A2(n_542),
.B(n_555),
.C(n_553),
.Y(n_587)
);

AOI21x1_ASAP7_75t_L g588 ( 
.A1(n_569),
.A2(n_568),
.B(n_530),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_525),
.B(n_550),
.Y(n_589)
);

NOR4xp25_ASAP7_75t_L g590 ( 
.A(n_493),
.B(n_500),
.C(n_527),
.D(n_554),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_503),
.Y(n_591)
);

OA21x2_ASAP7_75t_L g592 ( 
.A1(n_533),
.A2(n_537),
.B(n_558),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_545),
.Y(n_593)
);

O2A1O1Ixp33_ASAP7_75t_L g594 ( 
.A1(n_566),
.A2(n_505),
.B(n_556),
.C(n_504),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_561),
.B(n_495),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_497),
.A2(n_541),
.B1(n_507),
.B2(n_528),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_501),
.Y(n_597)
);

INVx6_ASAP7_75t_SL g598 ( 
.A(n_526),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_508),
.A2(n_502),
.B1(n_557),
.B2(n_539),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_514),
.Y(n_600)
);

NOR2x1_ASAP7_75t_L g601 ( 
.A(n_531),
.B(n_547),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_513),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_511),
.Y(n_603)
);

AO32x2_ASAP7_75t_L g604 ( 
.A1(n_520),
.A2(n_516),
.A3(n_514),
.B1(n_564),
.B2(n_532),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_565),
.B(n_509),
.Y(n_605)
);

AOI221xp5_ASAP7_75t_L g606 ( 
.A1(n_512),
.A2(n_521),
.B1(n_526),
.B2(n_510),
.C(n_517),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_520),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_522),
.B(n_429),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_523),
.B(n_421),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_551),
.B(n_317),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_492),
.A2(n_443),
.B(n_560),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_492),
.A2(n_443),
.B(n_560),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_549),
.B(n_413),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_549),
.B(n_413),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_499),
.B(n_413),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_499),
.B(n_413),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_499),
.B(n_413),
.Y(n_617)
);

NAND3xp33_ASAP7_75t_SL g618 ( 
.A(n_491),
.B(n_309),
.C(n_336),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_499),
.B(n_413),
.Y(n_619)
);

NOR2xp67_ASAP7_75t_L g620 ( 
.A(n_494),
.B(n_426),
.Y(n_620)
);

OAI21x1_ASAP7_75t_SL g621 ( 
.A1(n_551),
.A2(n_423),
.B(n_493),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_548),
.A2(n_544),
.B(n_563),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_519),
.Y(n_623)
);

BUFx8_ASAP7_75t_L g624 ( 
.A(n_507),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_506),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_522),
.B(n_429),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_515),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_494),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_494),
.B(n_426),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_515),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_549),
.B(n_413),
.Y(n_631)
);

AO31x2_ASAP7_75t_L g632 ( 
.A1(n_538),
.A2(n_543),
.A3(n_542),
.B(n_445),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_549),
.B(n_413),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_523),
.B(n_421),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_549),
.B(n_413),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_506),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_506),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_523),
.B(n_421),
.Y(n_638)
);

AO32x2_ASAP7_75t_L g639 ( 
.A1(n_542),
.A2(n_535),
.A3(n_389),
.B1(n_488),
.B2(n_448),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_549),
.B(n_413),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_519),
.Y(n_641)
);

NAND2x1p5_ASAP7_75t_L g642 ( 
.A(n_506),
.B(n_494),
.Y(n_642)
);

AOI21xp33_ASAP7_75t_L g643 ( 
.A1(n_522),
.A2(n_332),
.B(n_413),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_548),
.A2(n_544),
.B(n_563),
.Y(n_644)
);

OAI22x1_ASAP7_75t_L g645 ( 
.A1(n_498),
.A2(n_309),
.B1(n_307),
.B2(n_447),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_519),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_R g647 ( 
.A(n_494),
.B(n_426),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_515),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_494),
.B(n_426),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_519),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_492),
.A2(n_443),
.B(n_560),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_515),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_577),
.Y(n_653)
);

NAND3xp33_ASAP7_75t_L g654 ( 
.A(n_572),
.B(n_580),
.C(n_587),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_608),
.B(n_626),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_577),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_648),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_584),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_573),
.A2(n_622),
.B(n_644),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_641),
.Y(n_660)
);

AND2x4_ASAP7_75t_SL g661 ( 
.A(n_629),
.B(n_649),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_648),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_641),
.B(n_571),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_615),
.B(n_616),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_584),
.B(n_602),
.Y(n_665)
);

A2O1A1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_594),
.A2(n_602),
.B(n_640),
.C(n_635),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_579),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_617),
.B(n_619),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_630),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_643),
.B(n_613),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_586),
.A2(n_614),
.B1(n_633),
.B2(n_631),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_652),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_627),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_593),
.Y(n_674)
);

OA21x2_ASAP7_75t_L g675 ( 
.A1(n_611),
.A2(n_651),
.B(n_612),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_625),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_597),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_590),
.A2(n_607),
.B(n_588),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_570),
.A2(n_585),
.B(n_592),
.Y(n_679)
);

OA21x2_ASAP7_75t_L g680 ( 
.A1(n_606),
.A2(n_575),
.B(n_596),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_595),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_578),
.B(n_641),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_589),
.Y(n_683)
);

OA21x2_ASAP7_75t_L g684 ( 
.A1(n_575),
.A2(n_632),
.B(n_600),
.Y(n_684)
);

CKINVDCx16_ASAP7_75t_R g685 ( 
.A(n_647),
.Y(n_685)
);

BUFx12f_ASAP7_75t_L g686 ( 
.A(n_576),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_636),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_585),
.A2(n_599),
.B(n_601),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_574),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_646),
.A2(n_642),
.B(n_632),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_583),
.A2(n_618),
.B(n_638),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_581),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_591),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_637),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_605),
.A2(n_639),
.B(n_604),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_609),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_639),
.A2(n_604),
.B(n_610),
.Y(n_697)
);

NOR2x1_ASAP7_75t_SL g698 ( 
.A(n_571),
.B(n_650),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_609),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_583),
.A2(n_634),
.B(n_638),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_634),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_582),
.A2(n_628),
.B(n_620),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_571),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_623),
.B(n_645),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_598),
.Y(n_705)
);

AO21x2_ASAP7_75t_L g706 ( 
.A1(n_591),
.A2(n_624),
.B(n_629),
.Y(n_706)
);

NAND2x1p5_ASAP7_75t_L g707 ( 
.A(n_624),
.B(n_649),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_647),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_629),
.B(n_649),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_584),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_603),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_608),
.B(n_626),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_572),
.B(n_546),
.C(n_489),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_577),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_584),
.B(n_496),
.Y(n_715)
);

OAI21x1_ASAP7_75t_SL g716 ( 
.A1(n_580),
.A2(n_594),
.B(n_621),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_653),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_665),
.B(n_658),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_655),
.B(n_712),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_656),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_657),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_665),
.B(n_710),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_662),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_677),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_685),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_714),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_659),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_663),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_655),
.B(n_712),
.C(n_671),
.Y(n_729)
);

BUFx2_ASAP7_75t_SL g730 ( 
.A(n_708),
.Y(n_730)
);

BUFx10_ASAP7_75t_L g731 ( 
.A(n_661),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_663),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_670),
.A2(n_671),
.B1(n_715),
.B2(n_664),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_668),
.B(n_681),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_715),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_676),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_676),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_683),
.B(n_673),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_674),
.B(n_667),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_690),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_669),
.B(n_672),
.Y(n_741)
);

INVx3_ASAP7_75t_SL g742 ( 
.A(n_709),
.Y(n_742)
);

AO21x2_ASAP7_75t_L g743 ( 
.A1(n_678),
.A2(n_679),
.B(n_654),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_708),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_703),
.B(n_700),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_666),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_683),
.B(n_692),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_675),
.A2(n_688),
.B(n_716),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_697),
.Y(n_749)
);

OR2x6_ASAP7_75t_L g750 ( 
.A(n_691),
.B(n_704),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_695),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_698),
.B(n_682),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_687),
.B(n_694),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_660),
.Y(n_754)
);

AO21x2_ASAP7_75t_L g755 ( 
.A1(n_713),
.A2(n_704),
.B(n_691),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_736),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_749),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_740),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_719),
.B(n_689),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_718),
.B(n_684),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_718),
.B(n_684),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_729),
.A2(n_709),
.B1(n_680),
.B2(n_701),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_722),
.B(n_711),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_733),
.A2(n_745),
.B1(n_742),
.B2(n_709),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_745),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_717),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_754),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_735),
.B(n_699),
.Y(n_768)
);

AND2x4_ASAP7_75t_SL g769 ( 
.A(n_752),
.B(n_682),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_735),
.B(n_660),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_720),
.Y(n_771)
);

AND2x4_ASAP7_75t_SL g772 ( 
.A(n_752),
.B(n_696),
.Y(n_772)
);

NOR2x1_ASAP7_75t_L g773 ( 
.A(n_754),
.B(n_706),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_750),
.B(n_748),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_721),
.B(n_705),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_740),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_746),
.B(n_702),
.Y(n_777)
);

AO31x2_ASAP7_75t_L g778 ( 
.A1(n_746),
.A2(n_702),
.A3(n_706),
.B(n_693),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_727),
.A2(n_707),
.B(n_686),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_723),
.B(n_707),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_750),
.B(n_751),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_773),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_765),
.B(n_743),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_757),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_760),
.B(n_743),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_781),
.B(n_774),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_766),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_756),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_773),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_760),
.B(n_743),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_765),
.B(n_750),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_761),
.B(n_755),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_767),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_761),
.B(n_755),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_767),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_763),
.B(n_755),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_763),
.B(n_755),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_756),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_785),
.B(n_781),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_788),
.B(n_775),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_798),
.B(n_775),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_785),
.B(n_771),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_790),
.B(n_758),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_793),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_784),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_790),
.B(n_758),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_796),
.B(n_776),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_792),
.B(n_771),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_798),
.B(n_768),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_787),
.B(n_768),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_797),
.B(n_774),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_797),
.B(n_774),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_802),
.B(n_792),
.Y(n_813)
);

AND2x2_ASAP7_75t_SL g814 ( 
.A(n_804),
.B(n_793),
.Y(n_814)
);

AND2x2_ASAP7_75t_SL g815 ( 
.A(n_804),
.B(n_795),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_804),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_808),
.B(n_783),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_802),
.B(n_808),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_799),
.B(n_794),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_803),
.B(n_794),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_809),
.B(n_783),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_804),
.B(n_786),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_800),
.A2(n_779),
.B(n_759),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_807),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_805),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_801),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_819),
.B(n_799),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_818),
.B(n_803),
.Y(n_828)
);

AOI221xp5_ASAP7_75t_L g829 ( 
.A1(n_823),
.A2(n_812),
.B1(n_811),
.B2(n_810),
.C(n_806),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_826),
.A2(n_811),
.B1(n_812),
.B2(n_814),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_824),
.Y(n_831)
);

OAI221xp5_ASAP7_75t_L g832 ( 
.A1(n_816),
.A2(n_764),
.B1(n_779),
.B2(n_762),
.C(n_742),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_825),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_821),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_814),
.A2(n_742),
.B1(n_786),
.B2(n_795),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_815),
.A2(n_762),
.B1(n_791),
.B2(n_780),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_SL g837 ( 
.A1(n_815),
.A2(n_744),
.B(n_782),
.C(n_791),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_834),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_831),
.Y(n_839)
);

NOR3xp33_ASAP7_75t_L g840 ( 
.A(n_832),
.B(n_725),
.C(n_738),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_828),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_829),
.A2(n_822),
.B1(n_821),
.B2(n_813),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_833),
.Y(n_843)
);

NAND4xp25_ASAP7_75t_L g844 ( 
.A(n_840),
.B(n_836),
.C(n_830),
.D(n_835),
.Y(n_844)
);

NOR3x1_ASAP7_75t_L g845 ( 
.A(n_839),
.B(n_836),
.C(n_789),
.Y(n_845)
);

AOI221xp5_ASAP7_75t_L g846 ( 
.A1(n_841),
.A2(n_837),
.B1(n_819),
.B2(n_820),
.C(n_817),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_844),
.A2(n_846),
.B(n_840),
.Y(n_847)
);

NAND3xp33_ASAP7_75t_L g848 ( 
.A(n_845),
.B(n_842),
.C(n_838),
.Y(n_848)
);

NOR2x1_ASAP7_75t_L g849 ( 
.A(n_847),
.B(n_730),
.Y(n_849)
);

NAND3xp33_ASAP7_75t_L g850 ( 
.A(n_848),
.B(n_843),
.C(n_737),
.Y(n_850)
);

XNOR2x1_ASAP7_75t_L g851 ( 
.A(n_849),
.B(n_730),
.Y(n_851)
);

NOR2x1_ASAP7_75t_L g852 ( 
.A(n_850),
.B(n_780),
.Y(n_852)
);

AND4x1_ASAP7_75t_L g853 ( 
.A(n_852),
.B(n_731),
.C(n_747),
.D(n_827),
.Y(n_853)
);

NAND4xp75_ASAP7_75t_L g854 ( 
.A(n_851),
.B(n_731),
.C(n_777),
.D(n_734),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_854),
.A2(n_822),
.B(n_753),
.C(n_777),
.Y(n_855)
);

XNOR2xp5_ASAP7_75t_L g856 ( 
.A(n_853),
.B(n_753),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_854),
.B(n_731),
.Y(n_857)
);

INVxp33_ASAP7_75t_SL g858 ( 
.A(n_857),
.Y(n_858)
);

AOI22x1_ASAP7_75t_L g859 ( 
.A1(n_856),
.A2(n_731),
.B1(n_822),
.B2(n_789),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_855),
.Y(n_860)
);

OAI31xp33_ASAP7_75t_L g861 ( 
.A1(n_857),
.A2(n_732),
.A3(n_728),
.B(n_769),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_856),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_862),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_858),
.A2(n_817),
.B1(n_782),
.B2(n_770),
.Y(n_864)
);

OAI22x1_ASAP7_75t_L g865 ( 
.A1(n_860),
.A2(n_782),
.B1(n_724),
.B2(n_726),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_858),
.B(n_778),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_SL g867 ( 
.A1(n_861),
.A2(n_769),
.B(n_772),
.Y(n_867)
);

AOI21x1_ASAP7_75t_L g868 ( 
.A1(n_859),
.A2(n_741),
.B(n_726),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_863),
.A2(n_741),
.B(n_739),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_868),
.Y(n_870)
);

NOR2x2_ASAP7_75t_L g871 ( 
.A(n_867),
.B(n_825),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_865),
.B(n_778),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_870),
.B(n_866),
.Y(n_873)
);

AO21x2_ASAP7_75t_L g874 ( 
.A1(n_873),
.A2(n_869),
.B(n_872),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_874),
.A2(n_864),
.B1(n_871),
.B2(n_767),
.Y(n_875)
);


endmodule