module fake_jpeg_25418_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_45),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_50),
.B(n_72),
.Y(n_111)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_52),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_26),
.B1(n_31),
.B2(n_28),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_62),
.B1(n_74),
.B2(n_33),
.Y(n_95)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_28),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_54),
.B(n_25),
.Y(n_113)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_26),
.B1(n_31),
.B2(n_28),
.Y(n_62)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_26),
.B1(n_31),
.B2(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_77),
.B(n_86),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_54),
.C(n_61),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_103),
.C(n_113),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_30),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_51),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_64),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_88),
.Y(n_135)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_92),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_35),
.B1(n_24),
.B2(n_27),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_57),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_98),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_51),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_102),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_54),
.B(n_41),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_24),
.B1(n_27),
.B2(n_22),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_22),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_33),
.B1(n_22),
.B2(n_32),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_43),
.Y(n_116)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_115),
.A2(n_44),
.B(n_34),
.C(n_23),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_144),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_146),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_39),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_129),
.B(n_140),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_44),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_94),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_23),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_0),
.B(n_1),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_0),
.B(n_1),
.Y(n_157)
);

FAx1_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_35),
.CI(n_21),
.CON(n_144),
.SN(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_32),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_35),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_157),
.B(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_150),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_125),
.B(n_93),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_128),
.C(n_137),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_160),
.C(n_142),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_32),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_161),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_96),
.B1(n_100),
.B2(n_81),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_153),
.A2(n_164),
.B1(n_171),
.B2(n_177),
.Y(n_201)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_158),
.Y(n_209)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_141),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_34),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_101),
.C(n_90),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_163),
.B(n_168),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_130),
.A2(n_80),
.B1(n_81),
.B2(n_89),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_97),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_167),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_83),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_172),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_136),
.B(n_79),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_170),
.B(n_178),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_80),
.B1(n_109),
.B2(n_115),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_79),
.B1(n_92),
.B2(n_110),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_132),
.B1(n_119),
.B2(n_134),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_116),
.A2(n_129),
.B(n_140),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_119),
.A2(n_108),
.B1(n_90),
.B2(n_112),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_129),
.B(n_145),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_181),
.A2(n_205),
.B(n_213),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_182),
.A2(n_195),
.B1(n_198),
.B2(n_204),
.Y(n_225)
);

NAND2xp33_ASAP7_75t_R g188 ( 
.A(n_176),
.B(n_129),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_SL g215 ( 
.A(n_188),
.B(n_156),
.C(n_180),
.Y(n_215)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_191),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_210),
.C(n_20),
.Y(n_228)
);

AO22x2_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_122),
.B1(n_106),
.B2(n_99),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_18),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_175),
.A2(n_155),
.B1(n_151),
.B2(n_154),
.Y(n_198)
);

OAI22x1_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_84),
.B1(n_122),
.B2(n_35),
.Y(n_199)
);

OAI22x1_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_173),
.B1(n_165),
.B2(n_20),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_118),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_154),
.A2(n_121),
.B1(n_120),
.B2(n_21),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_159),
.A2(n_120),
.B1(n_23),
.B2(n_21),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_18),
.B1(n_16),
.B2(n_3),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_34),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_20),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_34),
.C(n_23),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_147),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_211),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_157),
.B(n_21),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_168),
.B(n_158),
.Y(n_214)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_215),
.A2(n_216),
.B1(n_224),
.B2(n_231),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_148),
.B(n_2),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_220),
.Y(n_250)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_20),
.Y(n_221)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_230),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_10),
.B(n_15),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_240),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_186),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_229),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_194),
.C(n_185),
.Y(n_254)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_18),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_204),
.A2(n_182),
.B1(n_199),
.B2(n_195),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_235),
.B1(n_205),
.B2(n_195),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_234),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_1),
.B(n_2),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_181),
.A2(n_18),
.B(n_16),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_201),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_16),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_207),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_239),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_200),
.B(n_10),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_16),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_244),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_243),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_187),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_201),
.B1(n_195),
.B2(n_210),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_253),
.B1(n_258),
.B2(n_260),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_256),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_213),
.B1(n_203),
.B2(n_183),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_257),
.C(n_238),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_203),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_222),
.B(n_11),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_197),
.B1(n_190),
.B2(n_4),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_216),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_221),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_252),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_255),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_265),
.B(n_267),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_251),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_262),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_225),
.B1(n_215),
.B2(n_230),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_282),
.B1(n_253),
.B2(n_249),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_228),
.C(n_241),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_272),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_246),
.A2(n_223),
.B(n_219),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_264),
.B(n_242),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_223),
.C(n_237),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_262),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_275),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_217),
.Y(n_274)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_250),
.B(n_234),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_278),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_235),
.C(n_233),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_232),
.Y(n_281)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_236),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_286),
.A2(n_269),
.B1(n_4),
.B2(n_6),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_290),
.B(n_292),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_268),
.B(n_257),
.CI(n_244),
.CON(n_291),
.SN(n_291)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_295),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_256),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_259),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_9),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_2),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_299),
.Y(n_310)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_270),
.C(n_266),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_303),
.C(n_304),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_278),
.B(n_279),
.Y(n_301)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_280),
.C(n_272),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_280),
.C(n_279),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_305),
.A2(n_311),
.B1(n_297),
.B2(n_288),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_291),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_293),
.B(n_9),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_309),
.B(n_285),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_294),
.A2(n_13),
.B1(n_14),
.B2(n_6),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_289),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_316),
.B(n_321),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_296),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_320),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_290),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_300),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_304),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_319),
.B(n_306),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_302),
.C(n_307),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_308),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_323),
.B(n_321),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_331),
.B(n_332),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_316),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_329),
.A2(n_328),
.B(n_322),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_330),
.B(n_313),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_334),
.C(n_302),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_308),
.B(n_291),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_14),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_3),
.B(n_4),
.Y(n_340)
);


endmodule