module fake_jpeg_15764_n_288 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_29),
.B(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_32),
.C(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_37),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_24),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_14),
.B1(n_15),
.B2(n_13),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_50),
.B1(n_14),
.B2(n_15),
.Y(n_55)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_14),
.B1(n_15),
.B2(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_20),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_27),
.B(n_44),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_41),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_70),
.B1(n_44),
.B2(n_48),
.Y(n_84)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_76)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_37),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_25),
.B(n_16),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_80),
.B(n_16),
.Y(n_94)
);

NOR2x1_ASAP7_75t_R g80 ( 
.A(n_52),
.B(n_50),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_32),
.C(n_50),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

AO22x2_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_43),
.B1(n_28),
.B2(n_33),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_70),
.B1(n_61),
.B2(n_64),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_57),
.B1(n_44),
.B2(n_38),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_27),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_42),
.C(n_28),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_99),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_101),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_38),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_108),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_60),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_98),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_80),
.B1(n_77),
.B2(n_88),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_38),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_63),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_57),
.B1(n_59),
.B2(n_65),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_85),
.B1(n_83),
.B2(n_81),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_83),
.B1(n_90),
.B2(n_73),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_107),
.A2(n_110),
.B1(n_85),
.B2(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_71),
.B(n_25),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_26),
.B(n_18),
.C(n_24),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_53),
.B1(n_58),
.B2(n_21),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_115),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_116),
.B(n_119),
.Y(n_148)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_133),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_84),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_121),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_84),
.B1(n_73),
.B2(n_89),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_124),
.A2(n_103),
.B1(n_107),
.B2(n_93),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_86),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_108),
.C(n_106),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_76),
.B(n_56),
.Y(n_129)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_94),
.B(n_101),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_113),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_24),
.B(n_17),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_19),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_87),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_87),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_139),
.Y(n_166)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_48),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_149),
.Y(n_170)
);

AOI22x1_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_109),
.B1(n_93),
.B2(n_63),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_117),
.B1(n_119),
.B2(n_131),
.Y(n_164)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_19),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_155),
.Y(n_172)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_130),
.B(n_17),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_127),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_154),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_62),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_62),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_151),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_120),
.B(n_121),
.C(n_124),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_139),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_134),
.B(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_126),
.B(n_129),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_178),
.B1(n_180),
.B2(n_153),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_126),
.B1(n_121),
.B2(n_111),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_163),
.A2(n_176),
.B1(n_181),
.B2(n_158),
.Y(n_201)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_152),
.B(n_125),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_175),
.Y(n_184)
);

NAND2x1_ASAP7_75t_SL g191 ( 
.A(n_168),
.B(n_180),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_173),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_136),
.A2(n_125),
.B1(n_91),
.B2(n_69),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_148),
.A2(n_17),
.B(n_26),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_179),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_134),
.B(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_56),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_18),
.B(n_67),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_68),
.B1(n_67),
.B2(n_21),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_135),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_144),
.C(n_143),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_192),
.C(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_158),
.B1(n_154),
.B2(n_148),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_159),
.B1(n_136),
.B2(n_169),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_191),
.A2(n_201),
.B1(n_204),
.B2(n_13),
.Y(n_220)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_149),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_195),
.A2(n_200),
.B(n_174),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_160),
.C(n_172),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_156),
.C(n_153),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_199),
.C(n_163),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_150),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_149),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_173),
.B1(n_172),
.B2(n_183),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_155),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_208),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_211),
.B1(n_213),
.B2(n_223),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_159),
.B1(n_169),
.B2(n_171),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_175),
.B1(n_174),
.B2(n_140),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_141),
.C(n_142),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_216),
.B(n_217),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_182),
.C(n_181),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_187),
.A2(n_165),
.B(n_72),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_48),
.C(n_33),
.Y(n_221)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_13),
.B1(n_49),
.B2(n_2),
.Y(n_223)
);

BUFx12_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_222),
.A2(n_203),
.B1(n_217),
.B2(n_212),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_214),
.A2(n_204),
.B1(n_201),
.B2(n_184),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_234),
.B1(n_216),
.B2(n_221),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_202),
.B1(n_191),
.B2(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_23),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_202),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_0),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_240),
.B(n_241),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_207),
.B(n_49),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_252),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_207),
.C(n_30),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_228),
.C(n_227),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_230),
.B(n_11),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_247),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_248),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_232),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_11),
.B(n_23),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_250),
.B(n_251),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_23),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_0),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_224),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_256),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_239),
.B(n_236),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_257),
.B(n_259),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_229),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_224),
.B(n_23),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_262),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_22),
.Y(n_262)
);

AOI21x1_ASAP7_75t_L g265 ( 
.A1(n_261),
.A2(n_0),
.B(n_1),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_265),
.A2(n_6),
.B(n_7),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_30),
.C(n_3),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_268),
.B(n_253),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_2),
.C(n_3),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_271),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_4),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_274),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_258),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_5),
.Y(n_276)
);

A2O1A1O1Ixp25_ASAP7_75t_L g281 ( 
.A1(n_276),
.A2(n_277),
.B(n_268),
.C(n_7),
.D(n_8),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_6),
.B(n_7),
.Y(n_277)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g279 ( 
.A1(n_278),
.A2(n_6),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_281),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_267),
.C(n_270),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_283),
.A2(n_275),
.B(n_8),
.Y(n_284)
);

AO21x1_ASAP7_75t_SL g285 ( 
.A1(n_284),
.A2(n_282),
.B(n_9),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_10),
.B(n_6),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_286),
.Y(n_287)
);

OA22x2_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_9),
.B1(n_10),
.B2(n_264),
.Y(n_288)
);


endmodule