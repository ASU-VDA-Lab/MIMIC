module fake_ariane_2633_n_1722 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1722);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1722;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_552;
wire n_348;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_9),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_8),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_1),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_5),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_20),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_23),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_83),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_23),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_5),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_1),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_21),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_108),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_115),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_91),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_34),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_54),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_93),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_13),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_32),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_58),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_3),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_79),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_103),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_7),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_29),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_138),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_101),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_35),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_32),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_16),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_54),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_114),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_86),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_65),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_31),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_25),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_88),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_156),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_2),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_16),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_136),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_133),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_21),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_2),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_99),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_87),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_48),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_35),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_121),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_13),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_137),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_130),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_4),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_89),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_127),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_24),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_37),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_25),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_125),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_45),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_105),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_117),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_26),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_77),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_147),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_109),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_43),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_151),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_6),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_38),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_122),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_56),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_149),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_92),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_40),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_43),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_140),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_85),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_27),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_10),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_62),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_40),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_143),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_3),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_33),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_78),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_59),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_61),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_135),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_55),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_73),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_76),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_41),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_0),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_128),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_148),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_102),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_59),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_45),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_7),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_146),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_26),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_70),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_104),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_15),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_111),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_119),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_157),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_31),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_41),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_6),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_39),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_153),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_47),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_27),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_20),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_30),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_69),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_56),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_134),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_80),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_90),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_36),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_96),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_74),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_22),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_154),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_95),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_19),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_63),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_44),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_4),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_132),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_9),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_49),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_12),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_68),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_42),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_18),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_72),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_50),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_0),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_112),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_18),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_34),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_30),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_39),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_107),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_150),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_139),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_52),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_22),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_216),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_187),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_162),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_158),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_166),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_166),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_267),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_172),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_165),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_159),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_167),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_172),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_175),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_162),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_224),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_168),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_160),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_164),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_175),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_216),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_185),
.Y(n_336)
);

INVxp33_ASAP7_75t_SL g337 ( 
.A(n_163),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_169),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_291),
.B(n_8),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_202),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_176),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_182),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_186),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_274),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_192),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_207),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_210),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_193),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_253),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_183),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_197),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_291),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_183),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_310),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_199),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_199),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_198),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_203),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_205),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_205),
.B(n_10),
.Y(n_361)
);

INVxp33_ASAP7_75t_SL g362 ( 
.A(n_211),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_209),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_219),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_209),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_215),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_215),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_217),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_223),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_217),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_225),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_225),
.B(n_11),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_228),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_220),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_184),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_228),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_226),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_208),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_234),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_234),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_230),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_232),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_240),
.B(n_11),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_223),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_224),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_224),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_238),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_161),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_161),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_240),
.B(n_12),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_204),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_241),
.Y(n_392)
);

BUFx2_ASAP7_75t_SL g393 ( 
.A(n_260),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_177),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_239),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_241),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_264),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_180),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_204),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_245),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_247),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_369),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_320),
.B(n_251),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_322),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_264),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_384),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_317),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_266),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_319),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_320),
.Y(n_411)
);

NAND2xp33_ASAP7_75t_L g412 ( 
.A(n_324),
.B(n_326),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_321),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_321),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_323),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_325),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_322),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_350),
.B(n_179),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_331),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_323),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_350),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_322),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_338),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_322),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_327),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_328),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_341),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_342),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_332),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_344),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_346),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_328),
.B(n_266),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_333),
.B(n_260),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_334),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_349),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_336),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_352),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_358),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_334),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_351),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_351),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_354),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_316),
.B(n_335),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_359),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_356),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_375),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_356),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_394),
.B(n_294),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_357),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_378),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_357),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_364),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_360),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_360),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_374),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_R g458 ( 
.A(n_330),
.B(n_170),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_363),
.B(n_177),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_377),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_340),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_363),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_365),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_365),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_366),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_381),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_382),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_366),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_387),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_401),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_367),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_367),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_368),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_395),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_370),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_411),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_418),
.B(n_329),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_411),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_402),
.B(n_370),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_402),
.B(n_362),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_413),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_441),
.B(n_400),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_405),
.B(n_353),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_408),
.B(n_339),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_441),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_441),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_413),
.B(n_414),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_414),
.Y(n_488)
);

AND2x4_ASAP7_75t_SL g489 ( 
.A(n_470),
.B(n_385),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_445),
.B(n_455),
.Y(n_490)
);

AND2x2_ASAP7_75t_SL g491 ( 
.A(n_412),
.B(n_361),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_441),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_415),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_445),
.B(n_343),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_441),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_455),
.B(n_371),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_441),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_421),
.B(n_422),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_442),
.Y(n_499)
);

INVxp33_ASAP7_75t_L g500 ( 
.A(n_418),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_442),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_442),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_442),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_442),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_442),
.B(n_449),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_427),
.B(n_373),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_428),
.Y(n_507)
);

BUFx4f_ASAP7_75t_L g508 ( 
.A(n_449),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_449),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_449),
.B(n_269),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_448),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_449),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_470),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_450),
.A2(n_337),
.B1(n_383),
.B2(n_372),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_436),
.B(n_376),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_423),
.B(n_318),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_471),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_450),
.B(n_345),
.Y(n_518)
);

AND2x2_ASAP7_75t_SL g519 ( 
.A(n_434),
.B(n_390),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_435),
.A2(n_301),
.B1(n_399),
.B2(n_391),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_444),
.B(n_379),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_416),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_444),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_471),
.Y(n_524)
);

AND2x2_ASAP7_75t_SL g525 ( 
.A(n_434),
.B(n_265),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_403),
.A2(n_309),
.B1(n_248),
.B2(n_250),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_451),
.B(n_379),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_451),
.B(n_380),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_462),
.B(n_380),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_471),
.B(n_269),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_471),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_471),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_462),
.B(n_285),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_448),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_463),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_471),
.B(n_285),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_452),
.B(n_394),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_464),
.B(n_392),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_475),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_475),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_470),
.B(n_386),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_465),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_465),
.B(n_392),
.Y(n_543)
);

BUFx10_ASAP7_75t_L g544 ( 
.A(n_410),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_472),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_475),
.B(n_288),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_420),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_475),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_475),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_475),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_472),
.B(n_396),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_470),
.B(n_398),
.Y(n_552)
);

INVx4_ASAP7_75t_SL g553 ( 
.A(n_404),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_404),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_403),
.A2(n_397),
.B1(n_396),
.B2(n_265),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_459),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_473),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_406),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_473),
.Y(n_559)
);

NAND2x1p5_ASAP7_75t_L g560 ( 
.A(n_459),
.B(n_397),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_425),
.B(n_294),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_406),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_429),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_431),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_443),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_443),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_438),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_461),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_430),
.B(n_288),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_407),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_432),
.Y(n_571)
);

NAND2x1_ASAP7_75t_L g572 ( 
.A(n_443),
.B(n_283),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_433),
.B(n_300),
.Y(n_573)
);

OAI22xp33_ASAP7_75t_L g574 ( 
.A1(n_437),
.A2(n_257),
.B1(n_261),
.B2(n_262),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_447),
.B(n_388),
.Y(n_575)
);

OR2x6_ASAP7_75t_L g576 ( 
.A(n_460),
.B(n_389),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_SL g577 ( 
.A(n_439),
.B(n_223),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_459),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_459),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_447),
.A2(n_221),
.B1(n_315),
.B2(n_314),
.Y(n_580)
);

AO22x2_ASAP7_75t_L g581 ( 
.A1(n_447),
.A2(n_221),
.B1(n_315),
.B2(n_314),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_440),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_452),
.B(n_275),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_453),
.Y(n_584)
);

AND2x2_ASAP7_75t_SL g585 ( 
.A(n_453),
.B(n_249),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_453),
.B(n_456),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_446),
.B(n_454),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_456),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_456),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_457),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_466),
.A2(n_263),
.B1(n_272),
.B2(n_273),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_468),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_467),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_468),
.B(n_300),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_468),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_469),
.Y(n_596)
);

AND2x6_ASAP7_75t_L g597 ( 
.A(n_409),
.B(n_311),
.Y(n_597)
);

OAI22xp33_ASAP7_75t_L g598 ( 
.A1(n_474),
.A2(n_277),
.B1(n_282),
.B2(n_286),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_409),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_404),
.A2(n_299),
.B1(n_292),
.B2(n_295),
.Y(n_600)
);

INVxp67_ASAP7_75t_SL g601 ( 
.A(n_419),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_417),
.A2(n_289),
.B1(n_298),
.B2(n_302),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_417),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_458),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_417),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_417),
.B(n_201),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_L g607 ( 
.A(n_424),
.B(n_171),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_419),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_419),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_424),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_424),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_426),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_595),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_491),
.B(n_190),
.Y(n_614)
);

INVxp33_ASAP7_75t_L g615 ( 
.A(n_537),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_560),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_484),
.B(n_244),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_491),
.B(n_311),
.Y(n_618)
);

NOR2x1p5_ASAP7_75t_L g619 ( 
.A(n_563),
.B(n_593),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_484),
.B(n_276),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_490),
.B(n_293),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_490),
.B(n_180),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_525),
.B(n_483),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_477),
.B(n_516),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_581),
.A2(n_206),
.B1(n_181),
.B2(n_189),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_525),
.B(n_181),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_483),
.B(n_189),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_563),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_519),
.B(n_494),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_519),
.A2(n_258),
.B1(n_283),
.B2(n_255),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_569),
.B(n_304),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_494),
.B(n_191),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_570),
.B(n_347),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_560),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_514),
.A2(n_305),
.B1(n_307),
.B2(n_191),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_552),
.B(n_513),
.Y(n_636)
);

NAND2x1_ASAP7_75t_L g637 ( 
.A(n_487),
.B(n_426),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_524),
.B(n_249),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_595),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_480),
.B(n_506),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_518),
.B(n_348),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_581),
.A2(n_268),
.B1(n_233),
.B2(n_235),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_480),
.B(n_206),
.Y(n_643)
);

NOR2xp67_ASAP7_75t_SL g644 ( 
.A(n_593),
.B(n_213),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_506),
.B(n_213),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_569),
.B(n_294),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_524),
.B(n_171),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_596),
.B(n_233),
.Y(n_648)
);

INVxp33_ASAP7_75t_SL g649 ( 
.A(n_590),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_521),
.B(n_235),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_521),
.B(n_242),
.Y(n_651)
);

BUFx6f_ASAP7_75t_SL g652 ( 
.A(n_596),
.Y(n_652)
);

NOR2xp67_ASAP7_75t_SL g653 ( 
.A(n_571),
.B(n_242),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_581),
.A2(n_278),
.B1(n_243),
.B2(n_256),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_476),
.Y(n_655)
);

OAI22xp33_ASAP7_75t_L g656 ( 
.A1(n_561),
.A2(n_576),
.B1(n_578),
.B2(n_556),
.Y(n_656)
);

NOR2xp67_ASAP7_75t_L g657 ( 
.A(n_604),
.B(n_173),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_528),
.B(n_243),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_528),
.B(n_256),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_595),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_522),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_500),
.B(n_355),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_500),
.B(n_564),
.Y(n_663)
);

O2A1O1Ixp5_ASAP7_75t_L g664 ( 
.A1(n_505),
.A2(n_279),
.B(n_308),
.C(n_297),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_529),
.B(n_268),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_529),
.B(n_556),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_556),
.B(n_278),
.Y(n_667)
);

AOI221x1_ASAP7_75t_L g668 ( 
.A1(n_594),
.A2(n_426),
.B1(n_312),
.B2(n_267),
.C(n_306),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_SL g669 ( 
.A(n_571),
.B(n_279),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_567),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_573),
.B(n_280),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_591),
.B(n_280),
.C(n_308),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_478),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_573),
.B(n_297),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_578),
.B(n_14),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_578),
.B(n_174),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_576),
.B(n_214),
.Y(n_677)
);

AND2x4_ASAP7_75t_SL g678 ( 
.A(n_544),
.B(n_547),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_481),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_487),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_558),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_579),
.B(n_178),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_585),
.A2(n_214),
.B1(n_252),
.B2(n_223),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_579),
.B(n_14),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_544),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_585),
.A2(n_252),
.B1(n_312),
.B2(n_306),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_579),
.B(n_15),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_487),
.A2(n_313),
.B1(n_188),
.B2(n_194),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_488),
.B(n_493),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_558),
.Y(n_690)
);

O2A1O1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_496),
.A2(n_17),
.B(n_19),
.C(n_24),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_L g692 ( 
.A1(n_576),
.A2(n_254),
.B1(n_196),
.B2(n_303),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_562),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_487),
.A2(n_246),
.B1(n_195),
.B2(n_296),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_568),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_562),
.Y(n_696)
);

AOI22x1_ASAP7_75t_L g697 ( 
.A1(n_507),
.A2(n_259),
.B1(n_200),
.B2(n_290),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_511),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_523),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_544),
.B(n_28),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_524),
.B(n_171),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_524),
.B(n_531),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_531),
.B(n_171),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_547),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_531),
.B(n_171),
.Y(n_705)
);

NOR2xp67_ASAP7_75t_L g706 ( 
.A(n_582),
.B(n_212),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_482),
.B(n_28),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_535),
.Y(n_708)
);

NOR2xp67_ASAP7_75t_L g709 ( 
.A(n_520),
.B(n_218),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_547),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_540),
.B(n_508),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_542),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_599),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_545),
.B(n_222),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_SL g715 ( 
.A(n_587),
.B(n_227),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_487),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_540),
.B(n_171),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_557),
.B(n_29),
.Y(n_718)
);

INVx8_ASAP7_75t_L g719 ( 
.A(n_498),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_540),
.B(n_171),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_559),
.Y(n_721)
);

NOR2xp67_ASAP7_75t_L g722 ( 
.A(n_587),
.B(n_229),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_599),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_566),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_485),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_489),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_575),
.B(n_231),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_485),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_575),
.B(n_479),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_486),
.Y(n_730)
);

NAND2x1p5_ASAP7_75t_L g731 ( 
.A(n_503),
.B(n_312),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_584),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_498),
.A2(n_271),
.B1(n_237),
.B2(n_287),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_503),
.B(n_36),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_565),
.B(n_236),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_588),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_489),
.B(n_37),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_589),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_533),
.A2(n_312),
.B1(n_306),
.B2(n_267),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_515),
.B(n_270),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_533),
.A2(n_312),
.B1(n_306),
.B2(n_267),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_527),
.B(n_284),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_592),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_495),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_549),
.B(n_281),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_495),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_497),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_583),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_549),
.B(n_38),
.Y(n_749)
);

BUFx5_ASAP7_75t_L g750 ( 
.A(n_498),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_538),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_498),
.Y(n_752)
);

OAI22xp33_ASAP7_75t_SL g753 ( 
.A1(n_526),
.A2(n_534),
.B1(n_600),
.B2(n_602),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_543),
.B(n_551),
.Y(n_754)
);

INVx8_ASAP7_75t_L g755 ( 
.A(n_498),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_586),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_555),
.B(n_42),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_533),
.B(n_44),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_533),
.B(n_46),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_492),
.B(n_46),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_603),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_603),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_624),
.B(n_541),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_729),
.A2(n_509),
.B(n_505),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_640),
.A2(n_580),
.B1(n_574),
.B2(n_598),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_617),
.B(n_597),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_641),
.B(n_510),
.Y(n_767)
);

AOI21x1_ASAP7_75t_L g768 ( 
.A1(n_702),
.A2(n_501),
.B(n_499),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_649),
.B(n_606),
.Y(n_769)
);

OAI21xp33_ASAP7_75t_L g770 ( 
.A1(n_620),
.A2(n_510),
.B(n_530),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_754),
.A2(n_601),
.B(n_492),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_655),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_752),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_752),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_629),
.B(n_597),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_618),
.A2(n_614),
.B(n_643),
.C(n_666),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_702),
.A2(n_548),
.B(n_504),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_689),
.A2(n_548),
.B(n_504),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_662),
.B(n_546),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_623),
.B(n_621),
.Y(n_780)
);

OAI21x1_ASAP7_75t_L g781 ( 
.A1(n_731),
.A2(n_497),
.B(n_499),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_618),
.A2(n_536),
.B(n_546),
.C(n_530),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_752),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_707),
.A2(n_577),
.B(n_539),
.C(n_548),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_751),
.B(n_597),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_615),
.B(n_504),
.Y(n_786)
);

O2A1O1Ixp5_ASAP7_75t_L g787 ( 
.A1(n_745),
.A2(n_572),
.B(n_512),
.C(n_539),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_671),
.B(n_597),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_671),
.B(n_597),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_656),
.B(n_554),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_756),
.A2(n_512),
.B(n_539),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_673),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_674),
.B(n_608),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_674),
.B(n_608),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_752),
.B(n_608),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_631),
.A2(n_532),
.B1(n_517),
.B2(n_502),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_693),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_627),
.B(n_554),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_632),
.B(n_532),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_614),
.A2(n_550),
.B(n_605),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_613),
.A2(n_605),
.B(n_609),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_639),
.A2(n_607),
.B(n_612),
.Y(n_802)
);

NOR2x1p5_ASAP7_75t_SL g803 ( 
.A(n_750),
.B(n_611),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_660),
.A2(n_607),
.B(n_610),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_680),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_646),
.B(n_553),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_716),
.A2(n_686),
.B1(n_719),
.B2(n_755),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_663),
.B(n_553),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_716),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_679),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_719),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_SL g812 ( 
.A(n_719),
.B(n_553),
.Y(n_812)
);

OR2x6_ASAP7_75t_L g813 ( 
.A(n_755),
.B(n_51),
.Y(n_813)
);

OAI21xp33_ASAP7_75t_L g814 ( 
.A1(n_630),
.A2(n_53),
.B(n_55),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_646),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_676),
.A2(n_100),
.B(n_64),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_635),
.A2(n_60),
.B(n_66),
.C(n_71),
.Y(n_817)
);

NAND3xp33_ASAP7_75t_L g818 ( 
.A(n_698),
.B(n_75),
.C(n_81),
.Y(n_818)
);

INVx11_ASAP7_75t_L g819 ( 
.A(n_652),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_636),
.A2(n_82),
.B1(n_84),
.B2(n_94),
.Y(n_820)
);

NOR2x1_ASAP7_75t_L g821 ( 
.A(n_628),
.B(n_97),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_628),
.B(n_98),
.Y(n_822)
);

O2A1O1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_753),
.A2(n_760),
.B(n_622),
.C(n_636),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_748),
.B(n_633),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_661),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_699),
.Y(n_826)
);

CKINVDCx10_ASAP7_75t_R g827 ( 
.A(n_652),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_SL g828 ( 
.A1(n_637),
.A2(n_106),
.B(n_110),
.C(n_113),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_760),
.A2(n_116),
.B(n_120),
.C(n_123),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_616),
.A2(n_124),
.B1(n_126),
.B2(n_141),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_686),
.A2(n_142),
.B1(n_144),
.B2(n_152),
.Y(n_831)
);

INVx4_ASAP7_75t_L g832 ( 
.A(n_755),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_667),
.A2(n_659),
.B(n_645),
.C(n_651),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_625),
.A2(n_654),
.B1(n_642),
.B2(n_683),
.Y(n_834)
);

NOR2x1p5_ASAP7_75t_SL g835 ( 
.A(n_750),
.B(n_761),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_708),
.Y(n_836)
);

OR2x6_ASAP7_75t_L g837 ( 
.A(n_677),
.B(n_695),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_650),
.A2(n_665),
.B(n_658),
.C(n_721),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_634),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_682),
.A2(n_735),
.B(n_711),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_712),
.B(n_626),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_675),
.B(n_684),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_SL g843 ( 
.A(n_669),
.B(n_700),
.C(n_672),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_685),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_675),
.A2(n_687),
.B1(n_684),
.B2(n_619),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_648),
.B(n_670),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_687),
.B(n_718),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_683),
.A2(n_727),
.B1(n_740),
.B2(n_742),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_696),
.Y(n_849)
);

AOI21xp33_ASAP7_75t_L g850 ( 
.A1(n_692),
.A2(n_757),
.B(n_714),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_762),
.A2(n_724),
.B(n_732),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_736),
.A2(n_738),
.B(n_743),
.Y(n_852)
);

CKINVDCx8_ASAP7_75t_R g853 ( 
.A(n_726),
.Y(n_853)
);

CKINVDCx10_ASAP7_75t_R g854 ( 
.A(n_677),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_750),
.B(n_685),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_718),
.B(n_648),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_664),
.A2(n_734),
.B(n_749),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_725),
.A2(n_744),
.B(n_730),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_750),
.B(n_704),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_678),
.B(n_677),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_723),
.B(n_706),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_728),
.A2(n_746),
.B(n_747),
.Y(n_862)
);

BUFx12f_ASAP7_75t_L g863 ( 
.A(n_737),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_696),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_734),
.A2(n_749),
.B(n_759),
.C(n_758),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_625),
.B(n_642),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_654),
.B(n_690),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_750),
.B(n_710),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_681),
.B(n_713),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_722),
.B(n_657),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_691),
.A2(n_737),
.B(n_720),
.C(n_647),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_678),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_731),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_715),
.A2(n_688),
.B(n_733),
.C(n_694),
.Y(n_874)
);

AOI21xp33_ASAP7_75t_L g875 ( 
.A1(n_709),
.A2(n_741),
.B(n_739),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_703),
.A2(n_705),
.B(n_717),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_638),
.B(n_739),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_668),
.A2(n_638),
.B(n_697),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_653),
.B(n_644),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_750),
.B(n_741),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_624),
.B(n_522),
.Y(n_881)
);

BUFx12f_ASAP7_75t_L g882 ( 
.A(n_726),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_729),
.A2(n_754),
.B(n_666),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_640),
.B(n_617),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_655),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_640),
.B(n_617),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_640),
.B(n_617),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_729),
.A2(n_754),
.B(n_666),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_640),
.A2(n_629),
.B1(n_617),
.B2(n_620),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_640),
.B(n_617),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_662),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_640),
.B(n_617),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_655),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_640),
.B(n_617),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_707),
.A2(n_640),
.B(n_617),
.C(n_620),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_695),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_656),
.B(n_563),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_640),
.A2(n_620),
.B(n_617),
.C(n_629),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_640),
.B(n_617),
.Y(n_899)
);

AO32x1_ASAP7_75t_L g900 ( 
.A1(n_723),
.A2(n_595),
.A3(n_696),
.B1(n_693),
.B2(n_724),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_640),
.A2(n_629),
.B1(n_617),
.B2(n_620),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_640),
.A2(n_629),
.B1(n_617),
.B2(n_620),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_729),
.A2(n_754),
.B(n_666),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_640),
.A2(n_629),
.B1(n_617),
.B2(n_620),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_629),
.A2(n_618),
.B(n_623),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_695),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_R g907 ( 
.A(n_726),
.B(n_590),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_729),
.A2(n_754),
.B(n_666),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_695),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_640),
.B(n_617),
.Y(n_910)
);

AOI21x1_ASAP7_75t_L g911 ( 
.A1(n_702),
.A2(n_701),
.B(n_647),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_649),
.B(n_317),
.Y(n_912)
);

CKINVDCx6p67_ASAP7_75t_R g913 ( 
.A(n_652),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_629),
.A2(n_618),
.B(n_623),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_640),
.A2(n_620),
.B1(n_617),
.B2(n_629),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_640),
.B(n_617),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_649),
.B(n_317),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_640),
.B(n_617),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_649),
.B(n_317),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_707),
.A2(n_640),
.B(n_617),
.C(n_620),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_640),
.B(n_617),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_649),
.B(n_317),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_729),
.A2(n_754),
.B(n_666),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_640),
.A2(n_620),
.B(n_617),
.C(n_629),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_649),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_663),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_649),
.B(n_317),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_640),
.A2(n_629),
.B1(n_617),
.B2(n_620),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_752),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_640),
.B(n_617),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_729),
.A2(n_754),
.B(n_666),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_628),
.B(n_619),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_729),
.A2(n_754),
.B(n_666),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_662),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_884),
.B(n_886),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_895),
.A2(n_920),
.B(n_898),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_763),
.B(n_846),
.Y(n_937)
);

NAND3xp33_ASAP7_75t_L g938 ( 
.A(n_847),
.B(n_842),
.C(n_845),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_883),
.A2(n_903),
.B(n_888),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_781),
.A2(n_768),
.B(n_911),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_825),
.Y(n_941)
);

INVxp67_ASAP7_75t_SL g942 ( 
.A(n_834),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_905),
.B(n_914),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_908),
.A2(n_931),
.B(n_923),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_887),
.B(n_890),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_892),
.B(n_894),
.Y(n_946)
);

AO221x1_ASAP7_75t_L g947 ( 
.A1(n_834),
.A2(n_831),
.B1(n_928),
.B2(n_889),
.C(n_904),
.Y(n_947)
);

AOI221x1_ASAP7_75t_L g948 ( 
.A1(n_865),
.A2(n_814),
.B1(n_889),
.B2(n_901),
.C(n_928),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_933),
.A2(n_840),
.B(n_899),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_772),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_910),
.B(n_916),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_918),
.A2(n_930),
.B(n_921),
.Y(n_952)
);

AOI21xp33_ASAP7_75t_L g953 ( 
.A1(n_765),
.A2(n_866),
.B(n_823),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_915),
.B(n_901),
.Y(n_954)
);

AOI21xp33_ASAP7_75t_L g955 ( 
.A1(n_765),
.A2(n_881),
.B(n_902),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_891),
.B(n_934),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_902),
.B(n_904),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_926),
.Y(n_958)
);

INVxp67_ASAP7_75t_SL g959 ( 
.A(n_867),
.Y(n_959)
);

AO31x2_ASAP7_75t_L g960 ( 
.A1(n_784),
.A2(n_880),
.A3(n_780),
.B(n_876),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_926),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_776),
.A2(n_815),
.B(n_905),
.C(n_914),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_800),
.A2(n_777),
.B(n_858),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_856),
.A2(n_857),
.B1(n_897),
.B2(n_769),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_800),
.A2(n_862),
.B(n_787),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_841),
.B(n_767),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_907),
.Y(n_967)
);

BUFx4f_ASAP7_75t_L g968 ( 
.A(n_913),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_774),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_851),
.A2(n_801),
.B(n_791),
.Y(n_970)
);

NAND2x1_ASAP7_75t_L g971 ( 
.A(n_832),
.B(n_811),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_852),
.A2(n_764),
.B(n_778),
.Y(n_972)
);

AOI21xp33_ASAP7_75t_L g973 ( 
.A1(n_912),
.A2(n_917),
.B(n_927),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_798),
.A2(n_771),
.B(n_833),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_766),
.A2(n_838),
.B(n_799),
.Y(n_975)
);

NAND2x1p5_ASAP7_75t_L g976 ( 
.A(n_774),
.B(n_783),
.Y(n_976)
);

OA21x2_ASAP7_75t_L g977 ( 
.A1(n_878),
.A2(n_816),
.B(n_804),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_824),
.B(n_919),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_850),
.A2(n_817),
.B(n_770),
.C(n_874),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_775),
.A2(n_794),
.B(n_793),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_925),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_779),
.B(n_792),
.Y(n_982)
);

O2A1O1Ixp5_ASAP7_75t_L g983 ( 
.A1(n_822),
.A2(n_795),
.B(n_861),
.C(n_859),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_802),
.A2(n_855),
.B(n_871),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_922),
.A2(n_843),
.B1(n_932),
.B2(n_786),
.Y(n_985)
);

AO21x1_ASAP7_75t_L g986 ( 
.A1(n_831),
.A2(n_788),
.B(n_789),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_829),
.A2(n_782),
.B(n_785),
.C(n_820),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_810),
.B(n_893),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_826),
.B(n_885),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_837),
.B(n_860),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_875),
.A2(n_836),
.B(n_805),
.C(n_809),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_SL g992 ( 
.A(n_853),
.B(n_882),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_863),
.B(n_932),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_807),
.B(n_929),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_796),
.A2(n_869),
.B(n_868),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_849),
.A2(n_864),
.B(n_806),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_818),
.A2(n_877),
.B(n_870),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_877),
.A2(n_773),
.B(n_821),
.Y(n_998)
);

O2A1O1Ixp5_ASAP7_75t_L g999 ( 
.A1(n_879),
.A2(n_773),
.B(n_900),
.C(n_811),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_830),
.A2(n_828),
.B(n_812),
.Y(n_1000)
);

AO31x2_ASAP7_75t_L g1001 ( 
.A1(n_900),
.A2(n_808),
.A3(n_835),
.B(n_803),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_783),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_783),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_900),
.A2(n_813),
.B(n_929),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_813),
.A2(n_837),
.B(n_872),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_813),
.A2(n_896),
.B(n_909),
.Y(n_1006)
);

NAND2x1p5_ASAP7_75t_L g1007 ( 
.A(n_929),
.B(n_839),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_SL g1008 ( 
.A1(n_844),
.A2(n_906),
.B(n_854),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_837),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_873),
.A2(n_844),
.B(n_839),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_819),
.B(n_873),
.Y(n_1011)
);

INVx8_ASAP7_75t_L g1012 ( 
.A(n_827),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_932),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_781),
.A2(n_768),
.B(n_911),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_781),
.A2(n_768),
.B(n_911),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_774),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_763),
.B(n_500),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_774),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_768),
.A2(n_781),
.B(n_840),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_842),
.B(n_905),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_883),
.A2(n_903),
.B(n_888),
.Y(n_1021)
);

AND2x6_ASAP7_75t_L g1022 ( 
.A(n_774),
.B(n_716),
.Y(n_1022)
);

AO21x1_ASAP7_75t_L g1023 ( 
.A1(n_842),
.A2(n_847),
.B(n_848),
.Y(n_1023)
);

BUFx5_ASAP7_75t_L g1024 ( 
.A(n_772),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_781),
.A2(n_768),
.B(n_911),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_883),
.A2(n_903),
.B(n_888),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_883),
.A2(n_903),
.B(n_888),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_895),
.A2(n_920),
.B(n_898),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_SL g1029 ( 
.A1(n_905),
.A2(n_914),
.B(n_823),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_825),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_883),
.A2(n_903),
.B(n_888),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_895),
.A2(n_920),
.B(n_924),
.C(n_898),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_883),
.A2(n_903),
.B(n_888),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_768),
.A2(n_840),
.B(n_790),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_772),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_842),
.B(n_905),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_932),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_895),
.A2(n_920),
.B(n_924),
.C(n_898),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_797),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_819),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_832),
.B(n_932),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_884),
.B(n_886),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_772),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_SL g1044 ( 
.A1(n_842),
.A2(n_847),
.B(n_884),
.Y(n_1044)
);

O2A1O1Ixp5_ASAP7_75t_L g1045 ( 
.A1(n_842),
.A2(n_847),
.B(n_857),
.C(n_865),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_895),
.A2(n_920),
.B(n_898),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_884),
.B(n_886),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_883),
.A2(n_903),
.B(n_888),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_884),
.B(n_886),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_884),
.B(n_886),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_884),
.B(n_886),
.Y(n_1051)
);

OAI21xp33_ASAP7_75t_L g1052 ( 
.A1(n_847),
.A2(n_842),
.B(n_895),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_895),
.A2(n_920),
.B(n_898),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_883),
.A2(n_903),
.B(n_888),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_895),
.A2(n_920),
.B(n_898),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_763),
.B(n_500),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_884),
.B(n_886),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_895),
.A2(n_920),
.B(n_898),
.Y(n_1058)
);

AO21x1_ASAP7_75t_L g1059 ( 
.A1(n_842),
.A2(n_847),
.B(n_848),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_772),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_819),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_895),
.A2(n_920),
.B(n_924),
.C(n_898),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_884),
.B(n_886),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_883),
.A2(n_903),
.B(n_888),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_842),
.A2(n_847),
.B1(n_640),
.B2(n_845),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_884),
.B(n_886),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_881),
.B(n_624),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_884),
.B(n_886),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_SL g1069 ( 
.A1(n_905),
.A2(n_914),
.B(n_823),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_763),
.B(n_500),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_895),
.A2(n_920),
.B(n_924),
.C(n_898),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_895),
.A2(n_920),
.B(n_898),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_884),
.B(n_886),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_774),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_781),
.A2(n_768),
.B(n_911),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_950),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1035),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_937),
.B(n_1017),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_1041),
.Y(n_1079)
);

AO32x1_ASAP7_75t_L g1080 ( 
.A1(n_1065),
.A2(n_964),
.A3(n_947),
.B1(n_1059),
.B2(n_1023),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1043),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1060),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_973),
.B(n_1068),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1056),
.B(n_1070),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_988),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_1041),
.Y(n_1086)
);

OAI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_957),
.A2(n_954),
.B1(n_948),
.B2(n_978),
.Y(n_1087)
);

OR2x6_ASAP7_75t_L g1088 ( 
.A(n_1008),
.B(n_1013),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_968),
.Y(n_1089)
);

INVxp67_ASAP7_75t_SL g1090 ( 
.A(n_958),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1068),
.B(n_952),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_1012),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_968),
.Y(n_1093)
);

BUFx4f_ASAP7_75t_SL g1094 ( 
.A(n_967),
.Y(n_1094)
);

NAND2xp33_ASAP7_75t_L g1095 ( 
.A(n_1052),
.B(n_935),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_942),
.B(n_945),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_1037),
.B(n_990),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1037),
.B(n_1005),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_R g1099 ( 
.A(n_1040),
.B(n_1061),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_1011),
.B(n_1006),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_955),
.A2(n_938),
.B(n_953),
.C(n_1045),
.Y(n_1101)
);

AO21x1_ASAP7_75t_L g1102 ( 
.A1(n_936),
.A2(n_1055),
.B(n_1028),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_942),
.B(n_946),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_989),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1011),
.B(n_1009),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_966),
.A2(n_1042),
.B1(n_1073),
.B2(n_1057),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1067),
.B(n_956),
.Y(n_1107)
);

AND2x6_ASAP7_75t_L g1108 ( 
.A(n_969),
.B(n_1016),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_982),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_941),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_1012),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_993),
.B(n_985),
.Y(n_1112)
);

O2A1O1Ixp5_ASAP7_75t_L g1113 ( 
.A1(n_1046),
.A2(n_1072),
.B(n_1058),
.C(n_1053),
.Y(n_1113)
);

NAND2xp33_ASAP7_75t_L g1114 ( 
.A(n_951),
.B(n_1047),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_1022),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1039),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1032),
.A2(n_1062),
.B(n_1071),
.C(n_1038),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1039),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_969),
.Y(n_1119)
);

BUFx4_ASAP7_75t_SL g1120 ( 
.A(n_981),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_939),
.A2(n_1031),
.B(n_1033),
.Y(n_1121)
);

BUFx2_ASAP7_75t_R g1122 ( 
.A(n_1030),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1022),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_1022),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_958),
.B(n_961),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_944),
.A2(n_1048),
.B(n_1021),
.Y(n_1126)
);

AND2x2_ASAP7_75t_SL g1127 ( 
.A(n_961),
.B(n_993),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_1002),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1049),
.B(n_1050),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_969),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1026),
.A2(n_1064),
.B(n_1054),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_1002),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_1007),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_1051),
.B(n_1063),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1027),
.A2(n_949),
.B(n_974),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1066),
.B(n_959),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_SL g1137 ( 
.A(n_992),
.B(n_1022),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1016),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1016),
.Y(n_1139)
);

INVxp67_ASAP7_75t_SL g1140 ( 
.A(n_976),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1024),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_1007),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1024),
.Y(n_1143)
);

INVx3_ASAP7_75t_SL g1144 ( 
.A(n_1012),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_986),
.A2(n_1024),
.B1(n_991),
.B2(n_979),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_959),
.B(n_1036),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1016),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1020),
.B(n_943),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1024),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1018),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_1003),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_975),
.A2(n_1032),
.B(n_1038),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_943),
.B(n_1062),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1071),
.B(n_1010),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1029),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_962),
.A2(n_991),
.B1(n_979),
.B2(n_987),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1018),
.B(n_1074),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1018),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1018),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_962),
.B(n_1069),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_1074),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1074),
.B(n_998),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1074),
.B(n_976),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_997),
.B(n_1004),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_996),
.A2(n_994),
.B1(n_980),
.B2(n_995),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_994),
.B(n_960),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_971),
.B(n_1001),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_960),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_960),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_960),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1000),
.A2(n_977),
.B1(n_965),
.B2(n_963),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_983),
.B(n_999),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_977),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_984),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_977),
.A2(n_972),
.B(n_970),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1001),
.B(n_999),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1001),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1034),
.B(n_940),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1001),
.Y(n_1179)
);

BUFx12f_ASAP7_75t_L g1180 ( 
.A(n_1044),
.Y(n_1180)
);

BUFx12f_ASAP7_75t_L g1181 ( 
.A(n_1044),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1014),
.Y(n_1182)
);

CKINVDCx11_ASAP7_75t_R g1183 ( 
.A(n_1015),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1025),
.B(n_1075),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1019),
.A2(n_1014),
.B(n_940),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1019),
.A2(n_1014),
.B(n_940),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_968),
.Y(n_1187)
);

BUFx2_ASAP7_75t_SL g1188 ( 
.A(n_1040),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_968),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1068),
.B(n_1065),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1068),
.B(n_1065),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1065),
.B(n_656),
.Y(n_1192)
);

AND2x2_ASAP7_75t_SL g1193 ( 
.A(n_957),
.B(n_625),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_941),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_947),
.A2(n_834),
.B1(n_641),
.B2(n_662),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1041),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_941),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_937),
.B(n_1017),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_957),
.A2(n_954),
.B(n_973),
.C(n_1065),
.Y(n_1199)
);

NOR2x1_ASAP7_75t_L g1200 ( 
.A(n_967),
.B(n_628),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1067),
.B(n_941),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_936),
.A2(n_715),
.B(n_1046),
.C(n_1028),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1065),
.B(n_656),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1067),
.B(n_941),
.Y(n_1204)
);

AOI21xp33_ASAP7_75t_SL g1205 ( 
.A1(n_973),
.A2(n_649),
.B(n_582),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_973),
.B(n_649),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1068),
.B(n_1065),
.Y(n_1207)
);

INVx6_ASAP7_75t_SL g1208 ( 
.A(n_1041),
.Y(n_1208)
);

AND2x6_ASAP7_75t_L g1209 ( 
.A(n_1041),
.B(n_774),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_957),
.A2(n_954),
.B1(n_1065),
.B2(n_847),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1022),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1068),
.B(n_1065),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1065),
.B(n_656),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_973),
.B(n_649),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1146),
.Y(n_1215)
);

CKINVDCx11_ASAP7_75t_R g1216 ( 
.A(n_1111),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1083),
.B(n_1206),
.Y(n_1217)
);

CKINVDCx14_ASAP7_75t_R g1218 ( 
.A(n_1092),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1076),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1193),
.A2(n_1192),
.B1(n_1213),
.B2(n_1203),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_1121),
.A2(n_1131),
.B(n_1126),
.Y(n_1221)
);

BUFx12f_ASAP7_75t_L g1222 ( 
.A(n_1187),
.Y(n_1222)
);

OAI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1190),
.A2(n_1191),
.B1(n_1212),
.B2(n_1207),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1077),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1167),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1110),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1160),
.B(n_1190),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1125),
.B(n_1166),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1195),
.A2(n_1102),
.B1(n_1212),
.B2(n_1191),
.Y(n_1229)
);

BUFx12f_ASAP7_75t_L g1230 ( 
.A(n_1088),
.Y(n_1230)
);

BUFx8_ASAP7_75t_SL g1231 ( 
.A(n_1089),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1081),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1082),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1175),
.A2(n_1172),
.B(n_1135),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1116),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1194),
.Y(n_1236)
);

CKINVDCx16_ASAP7_75t_R g1237 ( 
.A(n_1099),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1166),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1118),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1094),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1160),
.B(n_1090),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1170),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1167),
.Y(n_1243)
);

INVx4_ASAP7_75t_L g1244 ( 
.A(n_1108),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1164),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1164),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1085),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1162),
.B(n_1115),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1104),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1113),
.A2(n_1210),
.B(n_1199),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1207),
.B(n_1153),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1108),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1112),
.A2(n_1156),
.B1(n_1114),
.B2(n_1095),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1168),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1156),
.A2(n_1112),
.B1(n_1210),
.B2(n_1127),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1214),
.B(n_1134),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1145),
.A2(n_1117),
.B1(n_1101),
.B2(n_1106),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_1144),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1136),
.A2(n_1084),
.B1(n_1198),
.B2(n_1078),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1169),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1136),
.A2(n_1103),
.B1(n_1096),
.B2(n_1129),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1120),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1109),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_SL g1264 ( 
.A1(n_1137),
.A2(n_1091),
.B1(n_1164),
.B2(n_1096),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1132),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1103),
.B(n_1153),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1129),
.B(n_1107),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1177),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1202),
.A2(n_1152),
.B(n_1091),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1148),
.Y(n_1270)
);

INVx8_ASAP7_75t_L g1271 ( 
.A(n_1209),
.Y(n_1271)
);

INVx5_ASAP7_75t_L g1272 ( 
.A(n_1123),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1177),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1179),
.Y(n_1274)
);

OAI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1137),
.A2(n_1088),
.B1(n_1201),
.B2(n_1204),
.Y(n_1275)
);

BUFx12f_ASAP7_75t_L g1276 ( 
.A(n_1147),
.Y(n_1276)
);

OAI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1197),
.A2(n_1087),
.B1(n_1208),
.B2(n_1086),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1128),
.Y(n_1278)
);

INVxp67_ASAP7_75t_SL g1279 ( 
.A(n_1154),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1122),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1155),
.B(n_1176),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1093),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1100),
.A2(n_1098),
.B1(n_1124),
.B2(n_1211),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1162),
.B(n_1211),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1179),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1128),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1189),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1139),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1098),
.A2(n_1100),
.B1(n_1097),
.B2(n_1208),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1173),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1183),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1148),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1171),
.A2(n_1185),
.B(n_1186),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1182),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1138),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1163),
.B(n_1165),
.Y(n_1296)
);

AO21x2_ASAP7_75t_L g1297 ( 
.A1(n_1178),
.A2(n_1174),
.B(n_1141),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1108),
.Y(n_1298)
);

AO21x1_ASAP7_75t_L g1299 ( 
.A1(n_1080),
.A2(n_1143),
.B(n_1149),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1108),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1157),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1122),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1105),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_1188),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1209),
.A2(n_1181),
.B1(n_1180),
.B2(n_1086),
.Y(n_1305)
);

INVx4_ASAP7_75t_L g1306 ( 
.A(n_1209),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1158),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1161),
.B(n_1158),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1079),
.A2(n_1196),
.B1(n_1086),
.B2(n_1205),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1184),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1161),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1119),
.Y(n_1312)
);

NAND2x1p5_ASAP7_75t_L g1313 ( 
.A(n_1133),
.B(n_1142),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1119),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1119),
.Y(n_1315)
);

CKINVDCx16_ASAP7_75t_R g1316 ( 
.A(n_1151),
.Y(n_1316)
);

AO21x2_ASAP7_75t_L g1317 ( 
.A1(n_1184),
.A2(n_1080),
.B(n_1140),
.Y(n_1317)
);

BUFx2_ASAP7_75t_R g1318 ( 
.A(n_1080),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1130),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1200),
.A2(n_1130),
.B(n_1150),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1150),
.Y(n_1321)
);

CKINVDCx11_ASAP7_75t_R g1322 ( 
.A(n_1159),
.Y(n_1322)
);

BUFx12f_ASAP7_75t_L g1323 ( 
.A(n_1092),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1076),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1164),
.Y(n_1325)
);

AO31x2_ASAP7_75t_L g1326 ( 
.A1(n_1299),
.A2(n_1260),
.A3(n_1254),
.B(n_1242),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1254),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1223),
.B(n_1227),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_1216),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1215),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_1304),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1225),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1226),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1281),
.B(n_1227),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1281),
.B(n_1251),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1267),
.B(n_1251),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1236),
.Y(n_1337)
);

OAI21xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1253),
.A2(n_1229),
.B(n_1250),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1225),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1217),
.A2(n_1257),
.B(n_1255),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1294),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1238),
.Y(n_1342)
);

BUFx4f_ASAP7_75t_SL g1343 ( 
.A(n_1258),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1238),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1270),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1270),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1292),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1261),
.B(n_1256),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1259),
.B(n_1247),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1279),
.B(n_1310),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1225),
.B(n_1243),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1228),
.B(n_1241),
.Y(n_1352)
);

OR2x6_ASAP7_75t_L g1353 ( 
.A(n_1271),
.B(n_1244),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1235),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1243),
.B(n_1245),
.Y(n_1355)
);

AO21x1_ASAP7_75t_SL g1356 ( 
.A1(n_1269),
.A2(n_1241),
.B(n_1266),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1316),
.B(n_1237),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1239),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1266),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1246),
.B(n_1325),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1228),
.B(n_1290),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1294),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_SL g1363 ( 
.A(n_1262),
.Y(n_1363)
);

BUFx10_ASAP7_75t_L g1364 ( 
.A(n_1262),
.Y(n_1364)
);

OR2x6_ASAP7_75t_L g1365 ( 
.A(n_1271),
.B(n_1244),
.Y(n_1365)
);

AOI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1299),
.A2(n_1221),
.B(n_1293),
.Y(n_1366)
);

OR2x6_ASAP7_75t_L g1367 ( 
.A(n_1271),
.B(n_1244),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1278),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1282),
.B(n_1216),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1265),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1296),
.B(n_1219),
.Y(n_1371)
);

NAND2x1p5_ASAP7_75t_L g1372 ( 
.A(n_1306),
.B(n_1272),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1224),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1232),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1233),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1286),
.B(n_1273),
.Y(n_1376)
);

AO21x2_ASAP7_75t_L g1377 ( 
.A1(n_1277),
.A2(n_1317),
.B(n_1297),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1324),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1268),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1296),
.B(n_1273),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1249),
.B(n_1301),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1274),
.B(n_1308),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1304),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1303),
.Y(n_1384)
);

AO21x1_ASAP7_75t_SL g1385 ( 
.A1(n_1220),
.A2(n_1295),
.B(n_1307),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1285),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1274),
.B(n_1308),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1303),
.Y(n_1388)
);

CKINVDCx6p67_ASAP7_75t_R g1389 ( 
.A(n_1258),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1287),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1248),
.B(n_1284),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1297),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1297),
.Y(n_1393)
);

INVx4_ASAP7_75t_L g1394 ( 
.A(n_1252),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1263),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1317),
.B(n_1264),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1326),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1341),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1327),
.Y(n_1399)
);

INVxp67_ASAP7_75t_L g1400 ( 
.A(n_1356),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1352),
.B(n_1234),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1334),
.B(n_1234),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1359),
.B(n_1234),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1341),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1334),
.B(n_1318),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1330),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1335),
.B(n_1288),
.Y(n_1407)
);

INVxp67_ASAP7_75t_L g1408 ( 
.A(n_1356),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1352),
.B(n_1311),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1359),
.B(n_1313),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1335),
.B(n_1291),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1380),
.B(n_1291),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1362),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1330),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1351),
.B(n_1300),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1380),
.B(n_1248),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1362),
.Y(n_1417)
);

NOR2x1_ASAP7_75t_L g1418 ( 
.A(n_1394),
.B(n_1328),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1382),
.B(n_1248),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1340),
.B(n_1309),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1387),
.B(n_1350),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1361),
.B(n_1280),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1338),
.B(n_1322),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1350),
.B(n_1284),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1345),
.B(n_1313),
.Y(n_1425)
);

AO31x2_ASAP7_75t_L g1426 ( 
.A1(n_1392),
.A2(n_1393),
.A3(n_1379),
.B(n_1386),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1354),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1361),
.B(n_1302),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1376),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1333),
.Y(n_1430)
);

NAND3xp33_ASAP7_75t_L g1431 ( 
.A(n_1423),
.B(n_1348),
.C(n_1370),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1430),
.B(n_1337),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1429),
.B(n_1371),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1421),
.B(n_1360),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1430),
.B(n_1336),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1429),
.B(n_1371),
.Y(n_1436)
);

NAND4xp25_ASAP7_75t_L g1437 ( 
.A(n_1412),
.B(n_1369),
.C(n_1383),
.D(n_1331),
.Y(n_1437)
);

OAI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1420),
.A2(n_1349),
.B1(n_1396),
.B2(n_1381),
.C(n_1395),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1423),
.A2(n_1396),
.B(n_1357),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1421),
.B(n_1402),
.Y(n_1440)
);

OAI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_1420),
.A2(n_1395),
.B1(n_1289),
.B2(n_1373),
.C(n_1374),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1405),
.A2(n_1373),
.B1(n_1374),
.B2(n_1375),
.C(n_1378),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1421),
.B(n_1402),
.Y(n_1443)
);

NOR3xp33_ASAP7_75t_L g1444 ( 
.A(n_1418),
.B(n_1390),
.C(n_1368),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1407),
.B(n_1368),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1400),
.A2(n_1353),
.B(n_1367),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1407),
.B(n_1347),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1400),
.A2(n_1305),
.B1(n_1389),
.B2(n_1329),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1405),
.A2(n_1275),
.B1(n_1385),
.B2(n_1230),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1402),
.B(n_1346),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1398),
.B(n_1346),
.Y(n_1451)
);

OAI221xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1405),
.A2(n_1378),
.B1(n_1375),
.B2(n_1360),
.C(n_1342),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1408),
.A2(n_1365),
.B(n_1353),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1398),
.B(n_1342),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1413),
.B(n_1344),
.Y(n_1455)
);

OAI211xp5_ASAP7_75t_L g1456 ( 
.A1(n_1408),
.A2(n_1418),
.B(n_1413),
.C(n_1417),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1417),
.B(n_1344),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1409),
.B(n_1358),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1424),
.B(n_1355),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_L g1460 ( 
.A(n_1403),
.B(n_1314),
.C(n_1319),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1399),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1425),
.A2(n_1366),
.B(n_1320),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1411),
.A2(n_1389),
.B1(n_1394),
.B2(n_1283),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1412),
.A2(n_1218),
.B(n_1366),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1426),
.Y(n_1465)
);

NAND4xp25_ASAP7_75t_L g1466 ( 
.A(n_1412),
.B(n_1240),
.C(n_1287),
.D(n_1394),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1411),
.A2(n_1372),
.B(n_1298),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1416),
.B(n_1332),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1416),
.B(n_1332),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1415),
.B(n_1391),
.Y(n_1470)
);

NAND3xp33_ASAP7_75t_L g1471 ( 
.A(n_1425),
.B(n_1321),
.C(n_1312),
.Y(n_1471)
);

OAI221xp5_ASAP7_75t_SL g1472 ( 
.A1(n_1401),
.A2(n_1353),
.B1(n_1365),
.B2(n_1367),
.C(n_1315),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1419),
.B(n_1339),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1461),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1440),
.B(n_1443),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1444),
.B(n_1440),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1462),
.Y(n_1477)
);

OAI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1431),
.A2(n_1422),
.B1(n_1428),
.B2(n_1410),
.C(n_1397),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1433),
.B(n_1401),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1450),
.B(n_1406),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1432),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1461),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1455),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1457),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1470),
.B(n_1404),
.Y(n_1485)
);

INVxp67_ASAP7_75t_SL g1486 ( 
.A(n_1460),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1465),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1433),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1435),
.B(n_1406),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1436),
.B(n_1409),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1458),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1451),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1454),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1434),
.B(n_1415),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1447),
.Y(n_1495)
);

AND2x2_ASAP7_75t_SL g1496 ( 
.A(n_1442),
.B(n_1411),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1439),
.B(n_1414),
.Y(n_1497)
);

AND2x2_ASAP7_75t_SL g1498 ( 
.A(n_1449),
.B(n_1415),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1437),
.B(n_1343),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1471),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1459),
.B(n_1419),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1471),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1465),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1460),
.Y(n_1504)
);

OR2x6_ASAP7_75t_L g1505 ( 
.A(n_1477),
.B(n_1446),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1474),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1474),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1500),
.B(n_1502),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1482),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1496),
.A2(n_1438),
.B1(n_1431),
.B2(n_1463),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1500),
.B(n_1445),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1502),
.B(n_1422),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1504),
.B(n_1459),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1479),
.B(n_1422),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1504),
.B(n_1427),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1475),
.B(n_1468),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1486),
.B(n_1427),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1482),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1479),
.B(n_1428),
.Y(n_1519)
);

AND3x1_ASAP7_75t_L g1520 ( 
.A(n_1499),
.B(n_1464),
.C(n_1467),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1487),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1489),
.Y(n_1522)
);

NAND2x2_ASAP7_75t_L g1523 ( 
.A(n_1481),
.B(n_1240),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1475),
.B(n_1469),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1494),
.B(n_1415),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1489),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1483),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1475),
.B(n_1494),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1494),
.B(n_1469),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1497),
.B(n_1488),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1494),
.B(n_1473),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1476),
.B(n_1473),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1488),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1497),
.B(n_1428),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1493),
.Y(n_1535)
);

INVxp67_ASAP7_75t_SL g1536 ( 
.A(n_1486),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1483),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1484),
.Y(n_1538)
);

NAND3xp33_ASAP7_75t_SL g1539 ( 
.A(n_1477),
.B(n_1456),
.C(n_1448),
.Y(n_1539)
);

NOR3xp33_ASAP7_75t_L g1540 ( 
.A(n_1478),
.B(n_1441),
.C(n_1452),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1487),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1484),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1481),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1528),
.B(n_1476),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1536),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1521),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1521),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1507),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1508),
.B(n_1492),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1540),
.B(n_1496),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1543),
.B(n_1323),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1512),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1507),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1506),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1509),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1541),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1541),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1512),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1518),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1514),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1514),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1533),
.Y(n_1562)
);

NAND2x1p5_ASAP7_75t_L g1563 ( 
.A(n_1520),
.B(n_1496),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1539),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1533),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1528),
.B(n_1476),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1515),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1525),
.B(n_1476),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1525),
.B(n_1501),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1535),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1535),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1510),
.A2(n_1498),
.B1(n_1478),
.B2(n_1377),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1527),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1537),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1511),
.B(n_1492),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1523),
.Y(n_1576)
);

INVx2_ASAP7_75t_SL g1577 ( 
.A(n_1523),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1530),
.B(n_1490),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1522),
.B(n_1491),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_1534),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1534),
.B(n_1485),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1519),
.Y(n_1582)
);

OAI31xp33_ASAP7_75t_L g1583 ( 
.A1(n_1530),
.A2(n_1517),
.A3(n_1519),
.B(n_1526),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1525),
.B(n_1501),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1538),
.B(n_1491),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1542),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1569),
.B(n_1532),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1558),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1548),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1548),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1563),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1563),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1566),
.B(n_1505),
.Y(n_1593)
);

AO21x2_ASAP7_75t_L g1594 ( 
.A1(n_1550),
.A2(n_1513),
.B(n_1493),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1564),
.B(n_1516),
.Y(n_1595)
);

CKINVDCx16_ASAP7_75t_R g1596 ( 
.A(n_1551),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1563),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1578),
.B(n_1490),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1566),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1553),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1572),
.B(n_1485),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_L g1602 ( 
.A(n_1549),
.B(n_1505),
.Y(n_1602)
);

NOR2xp67_ASAP7_75t_L g1603 ( 
.A(n_1572),
.B(n_1532),
.Y(n_1603)
);

OAI21x1_ASAP7_75t_L g1604 ( 
.A1(n_1546),
.A2(n_1503),
.B(n_1487),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1553),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1562),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1545),
.B(n_1516),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1549),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1562),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1578),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1580),
.B(n_1524),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1565),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1569),
.B(n_1584),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1575),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1565),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1554),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1552),
.B(n_1323),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1573),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1566),
.A2(n_1505),
.B1(n_1498),
.B2(n_1481),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1582),
.B(n_1480),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1582),
.B(n_1480),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1546),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1603),
.A2(n_1601),
.B1(n_1610),
.B2(n_1599),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1608),
.B(n_1583),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1614),
.B(n_1560),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1592),
.A2(n_1561),
.B1(n_1560),
.B2(n_1505),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1594),
.A2(n_1581),
.B(n_1577),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1596),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1617),
.B(n_1597),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1618),
.Y(n_1630)
);

AO21x1_ASAP7_75t_L g1631 ( 
.A1(n_1616),
.A2(n_1571),
.B(n_1570),
.Y(n_1631)
);

OAI21xp33_ASAP7_75t_L g1632 ( 
.A1(n_1595),
.A2(n_1567),
.B(n_1579),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1591),
.A2(n_1560),
.B1(n_1561),
.B2(n_1498),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1599),
.A2(n_1593),
.B1(n_1598),
.B2(n_1566),
.Y(n_1634)
);

INVxp67_ASAP7_75t_L g1635 ( 
.A(n_1588),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1594),
.B(n_1561),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1591),
.A2(n_1576),
.B1(n_1577),
.B2(n_1567),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1594),
.A2(n_1576),
.B(n_1585),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1613),
.B(n_1544),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1602),
.A2(n_1544),
.B(n_1573),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1593),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1589),
.Y(n_1642)
);

BUFx6f_ASAP7_75t_L g1643 ( 
.A(n_1593),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1619),
.A2(n_1586),
.B(n_1574),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1589),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1611),
.B(n_1574),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1598),
.B(n_1607),
.Y(n_1647)
);

OAI32xp33_ASAP7_75t_L g1648 ( 
.A1(n_1620),
.A2(n_1568),
.A3(n_1571),
.B1(n_1570),
.B2(n_1586),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1613),
.B(n_1584),
.Y(n_1649)
);

NAND2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1628),
.B(n_1384),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1628),
.B(n_1587),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1635),
.B(n_1587),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1641),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1641),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1643),
.B(n_1363),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1643),
.B(n_1620),
.Y(n_1656)
);

NAND2x1_ASAP7_75t_L g1657 ( 
.A(n_1639),
.B(n_1568),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1647),
.B(n_1621),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1642),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1649),
.B(n_1529),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1646),
.B(n_1621),
.Y(n_1661)
);

NOR2xp67_ASAP7_75t_SL g1662 ( 
.A(n_1643),
.B(n_1276),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1625),
.Y(n_1663)
);

AND2x2_ASAP7_75t_SL g1664 ( 
.A(n_1624),
.B(n_1630),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1632),
.B(n_1590),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1623),
.A2(n_1622),
.B1(n_1557),
.B2(n_1546),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1636),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1634),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1664),
.B(n_1645),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1651),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1653),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1664),
.A2(n_1631),
.B(n_1638),
.Y(n_1672)
);

NOR3xp33_ASAP7_75t_L g1673 ( 
.A(n_1654),
.B(n_1629),
.C(n_1640),
.Y(n_1673)
);

NAND4xp25_ASAP7_75t_SL g1674 ( 
.A(n_1668),
.B(n_1627),
.C(n_1637),
.D(n_1644),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_L g1675 ( 
.A(n_1659),
.B(n_1590),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1663),
.A2(n_1648),
.B1(n_1633),
.B2(n_1626),
.C(n_1605),
.Y(n_1676)
);

NOR3xp33_ASAP7_75t_SL g1677 ( 
.A(n_1652),
.B(n_1605),
.C(n_1600),
.Y(n_1677)
);

AOI21xp33_ASAP7_75t_L g1678 ( 
.A1(n_1656),
.A2(n_1622),
.B(n_1606),
.Y(n_1678)
);

NOR4xp25_ASAP7_75t_L g1679 ( 
.A(n_1667),
.B(n_1615),
.C(n_1612),
.D(n_1609),
.Y(n_1679)
);

NOR2xp67_ASAP7_75t_L g1680 ( 
.A(n_1674),
.B(n_1655),
.Y(n_1680)
);

AOI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1672),
.A2(n_1656),
.B1(n_1667),
.B2(n_1650),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1677),
.A2(n_1666),
.B(n_1650),
.Y(n_1682)
);

NAND4xp75_ASAP7_75t_L g1683 ( 
.A(n_1671),
.B(n_1658),
.C(n_1665),
.D(n_1655),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1670),
.B(n_1661),
.Y(n_1684)
);

AOI211xp5_ASAP7_75t_L g1685 ( 
.A1(n_1679),
.A2(n_1662),
.B(n_1606),
.C(n_1609),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1673),
.B(n_1660),
.Y(n_1686)
);

O2A1O1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1669),
.A2(n_1678),
.B(n_1676),
.C(n_1675),
.Y(n_1687)
);

AOI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1672),
.A2(n_1615),
.B1(n_1612),
.B2(n_1600),
.C(n_1657),
.Y(n_1688)
);

XNOR2x1_ASAP7_75t_SL g1689 ( 
.A(n_1671),
.B(n_1231),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1681),
.B(n_1554),
.Y(n_1690)
);

NAND3xp33_ASAP7_75t_L g1691 ( 
.A(n_1687),
.B(n_1680),
.C(n_1688),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1686),
.B(n_1555),
.Y(n_1692)
);

NAND5xp2_ASAP7_75t_SL g1693 ( 
.A(n_1682),
.B(n_1364),
.C(n_1529),
.D(n_1531),
.E(n_1524),
.Y(n_1693)
);

NOR3xp33_ASAP7_75t_L g1694 ( 
.A(n_1683),
.B(n_1557),
.C(n_1556),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1684),
.B(n_1364),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1691),
.A2(n_1685),
.B1(n_1689),
.B2(n_1557),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1694),
.B(n_1555),
.Y(n_1697)
);

AO22x2_ASAP7_75t_L g1698 ( 
.A1(n_1690),
.A2(n_1695),
.B1(n_1692),
.B2(n_1547),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1693),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1690),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1692),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1692),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1698),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1696),
.A2(n_1559),
.B1(n_1547),
.B2(n_1556),
.Y(n_1704)
);

AND3x1_ASAP7_75t_L g1705 ( 
.A(n_1701),
.B(n_1559),
.C(n_1231),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1702),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1698),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1705),
.B(n_1699),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1703),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1706),
.B(n_1700),
.Y(n_1710)
);

XNOR2x1_ASAP7_75t_L g1711 ( 
.A(n_1708),
.B(n_1705),
.Y(n_1711)
);

NAND3xp33_ASAP7_75t_SL g1712 ( 
.A(n_1711),
.B(n_1707),
.C(n_1710),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1712),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1712),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1714),
.B(n_1713),
.Y(n_1715)
);

OAI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1714),
.A2(n_1709),
.B1(n_1704),
.B2(n_1697),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1715),
.A2(n_1604),
.B1(n_1282),
.B2(n_1222),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1716),
.B(n_1604),
.Y(n_1718)
);

NAND3xp33_ASAP7_75t_L g1719 ( 
.A(n_1718),
.B(n_1388),
.C(n_1384),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1719),
.A2(n_1717),
.B1(n_1276),
.B2(n_1222),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1720),
.A2(n_1388),
.B1(n_1364),
.B2(n_1466),
.C(n_1495),
.Y(n_1721)
);

AOI211xp5_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1446),
.B(n_1453),
.C(n_1472),
.Y(n_1722)
);


endmodule