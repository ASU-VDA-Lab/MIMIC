module fake_netlist_6_3910_n_3857 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_440, n_587, n_695, n_507, n_580, n_762, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_783, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_805, n_396, n_495, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_442, n_480, n_142, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_807, n_739, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_768, n_38, n_471, n_289, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_727, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_797, n_666, n_371, n_795, n_770, n_567, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_752, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_803, n_290, n_220, n_809, n_118, n_224, n_48, n_25, n_93, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_779, n_9, n_800, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_777, n_407, n_450, n_103, n_808, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_745, n_654, n_323, n_606, n_393, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_731, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_792, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_788, n_325, n_767, n_804, n_329, n_464, n_600, n_802, n_561, n_33, n_477, n_549, n_533, n_408, n_806, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_743, n_766, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_728, n_681, n_729, n_110, n_151, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_722, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_736, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_778, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_3857);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_762;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_783;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_805;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_807;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_727;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_567;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_800;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_777;
input n_407;
input n_450;
input n_103;
input n_808;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_745;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_731;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_792;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_788;
input n_325;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_802;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_806;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_722;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_778;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_3857;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_2576;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_1674;
wire n_1199;
wire n_3392;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_3152;
wire n_3579;
wire n_1212;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_3844;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_3741;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_3465;
wire n_1975;
wire n_1743;
wire n_1930;
wire n_1009;
wire n_2405;
wire n_3706;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_1371;
wire n_873;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_836;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_2356;
wire n_1143;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_2480;
wire n_2739;
wire n_1300;
wire n_3023;
wire n_822;
wire n_3232;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3316;
wire n_2212;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_943;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_940;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_3765;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_1088;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3368;
wire n_917;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_1446;
wire n_2591;
wire n_3507;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_913;
wire n_1658;
wire n_2593;
wire n_867;
wire n_3506;
wire n_3568;
wire n_3269;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_1967;
wire n_1193;
wire n_1054;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_824;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_3732;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_3446;
wire n_3317;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_3716;
wire n_1873;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_1866;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3842;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1605;
wire n_1330;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_1014;
wire n_3734;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_1265;
wire n_2711;
wire n_3490;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_3247;
wire n_871;
wire n_3069;
wire n_922;
wire n_1760;
wire n_1335;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_1801;
wire n_928;
wire n_835;
wire n_2347;
wire n_850;
wire n_1214;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_825;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_1588;
wire n_3785;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_1515;
wire n_961;
wire n_3510;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_890;
wire n_2377;
wire n_3271;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_3545;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_3073;
wire n_2431;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_3253;
wire n_1779;
wire n_1465;
wire n_3337;
wire n_3431;
wire n_3450;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_1627;
wire n_1164;
wire n_1295;
wire n_2954;
wire n_3477;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1565;
wire n_1067;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_3616;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_2535;
wire n_1880;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_963;
wire n_2767;
wire n_3793;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1714;
wire n_872;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_2897;
wire n_847;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_1913;
wire n_3608;
wire n_837;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_3491;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3426;
wire n_3158;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2643;
wire n_2590;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_3470;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_1432;
wire n_2208;
wire n_843;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_2134;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_947;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_1049;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2896;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_998;
wire n_3200;
wire n_1665;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_3390;
wire n_3656;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_1178;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1048;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_1021;
wire n_931;
wire n_3393;
wire n_811;
wire n_2442;
wire n_1207;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_3641;
wire n_1837;
wire n_1314;
wire n_2218;
wire n_831;
wire n_964;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_2748;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2323;
wire n_1220;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_1775;
wire n_1286;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_3364;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_3425;
wire n_2384;
wire n_1745;
wire n_914;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_3547;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_2249;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3284;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3205;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_906;
wire n_2315;
wire n_1733;
wire n_1077;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_3016;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1129;
wire n_2829;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_3338;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3276;
wire n_1934;
wire n_3250;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_845;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_892;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1037;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_901;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_1108;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_3819;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_3501;
wire n_1840;
wire n_1152;
wire n_1705;
wire n_3262;
wire n_3544;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_2376;
wire n_972;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_1637;
wire n_934;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_3712;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_2154;
wire n_2727;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3469;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_3156;
wire n_1931;
wire n_2083;
wire n_1269;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_2128;
wire n_1650;
wire n_1794;
wire n_1962;
wire n_1236;
wire n_1045;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_834;
wire n_2695;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1746;
wire n_1002;
wire n_1325;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_3524;
wire n_2671;
wire n_2888;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_3711;
wire n_3776;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_3511;
wire n_2054;
wire n_876;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_841;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1882;
wire n_1023;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1929;
wire n_1007;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_3806;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_933;
wire n_3343;
wire n_3303;
wire n_978;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_823;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1120;
wire n_1583;
wire n_832;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_1848;
wire n_1785;
wire n_1147;
wire n_1114;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_957;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3336;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_3584;
wire n_1414;
wire n_3486;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_3556;
wire n_2034;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_2444;
wire n_839;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3697;
wire n_3643;
wire n_1584;
wire n_2425;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_829;
wire n_1156;
wire n_3123;
wire n_2600;
wire n_984;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_859;
wire n_3086;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_3285;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_3478;
wire n_1349;
wire n_2071;
wire n_1144;
wire n_3669;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_3344;
wire n_2334;
wire n_3295;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1133;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1629;
wire n_2221;
wire n_1170;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_2553;
wire n_1040;
wire n_915;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_3815;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_3274;
wire n_2899;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_3504;
wire n_1449;
wire n_827;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_434),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_169),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_68),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_664),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_533),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_502),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_170),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_480),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_387),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_263),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_484),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_223),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_791),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_109),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_11),
.Y(n_825)
);

BUFx10_ASAP7_75t_L g826 ( 
.A(n_580),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_220),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_681),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_581),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_258),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_89),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_75),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_694),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_739),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_723),
.Y(n_835)
);

BUFx5_ASAP7_75t_L g836 ( 
.A(n_44),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_194),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_112),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_778),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_357),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_716),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_36),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_185),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_648),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_87),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_192),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_310),
.Y(n_847)
);

BUFx5_ASAP7_75t_L g848 ( 
.A(n_191),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_734),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_249),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_692),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_495),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_502),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_341),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_752),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_466),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_109),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_126),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_529),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_55),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_210),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_416),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_544),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_31),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_383),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_203),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_404),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_414),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_672),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_732),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_593),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_164),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_114),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_290),
.Y(n_874)
);

INVx1_ASAP7_75t_SL g875 ( 
.A(n_705),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_129),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_431),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_115),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_528),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_351),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_436),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_21),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_240),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_232),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_568),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_529),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_720),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_553),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_752),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_687),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_785),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_170),
.Y(n_892)
);

CKINVDCx14_ASAP7_75t_R g893 ( 
.A(n_469),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_352),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_432),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_253),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_635),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_749),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_37),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_738),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_505),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_521),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_693),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_601),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_236),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_697),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_5),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_371),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_425),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_669),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_561),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_61),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_724),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_571),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_652),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_136),
.Y(n_916)
);

INVxp67_ASAP7_75t_SL g917 ( 
.A(n_755),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_246),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_80),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_750),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_726),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_419),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_568),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_53),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_375),
.Y(n_925)
);

INVxp67_ASAP7_75t_SL g926 ( 
.A(n_421),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_252),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_501),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_29),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_48),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_771),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_73),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_286),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_668),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_256),
.Y(n_935)
);

BUFx10_ASAP7_75t_L g936 ( 
.A(n_39),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_730),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_60),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_606),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_18),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_496),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_665),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_585),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_744),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_189),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_458),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_151),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_387),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_736),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_747),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_145),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_227),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_148),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_447),
.Y(n_954)
);

BUFx5_ASAP7_75t_L g955 ( 
.A(n_457),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_666),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_295),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_706),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_229),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_271),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_757),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_240),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_376),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_204),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_722),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_467),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_505),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_534),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_372),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_741),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_672),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_689),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_487),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_464),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_755),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_277),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_115),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_110),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_574),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_144),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_226),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_760),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_534),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_749),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_793),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_392),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_378),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_90),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_528),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_718),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_737),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_594),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_649),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_457),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_532),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_443),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_595),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_609),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_25),
.Y(n_999)
);

BUFx10_ASAP7_75t_L g1000 ( 
.A(n_268),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_270),
.Y(n_1001)
);

CKINVDCx16_ASAP7_75t_R g1002 ( 
.A(n_786),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_372),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_623),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_725),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_711),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_288),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_543),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_335),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_579),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_674),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_31),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_268),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_456),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_130),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_751),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_292),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_256),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_254),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_221),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_207),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_364),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_8),
.Y(n_1023)
);

CKINVDCx14_ASAP7_75t_R g1024 ( 
.A(n_180),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_545),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_29),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_337),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_5),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_214),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_759),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_780),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_317),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_124),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_521),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_801),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_276),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_558),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_775),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_3),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_208),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_714),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_293),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_547),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_39),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_72),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_728),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_380),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_3),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_643),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_756),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_435),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_537),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_471),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_682),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_712),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_299),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_788),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_743),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_726),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_27),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_355),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_285),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_512),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_608),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_747),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_538),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_703),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_127),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_101),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_373),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_51),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_681),
.Y(n_1072)
);

BUFx5_ASAP7_75t_L g1073 ( 
.A(n_52),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_77),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_97),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_402),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_696),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_471),
.Y(n_1078)
);

CKINVDCx16_ASAP7_75t_R g1079 ( 
.A(n_147),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_179),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_715),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_185),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_150),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_323),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_66),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_657),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_77),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_139),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_253),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_404),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_421),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_255),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_56),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_757),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_249),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_180),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_283),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_501),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_95),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_86),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_292),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_9),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_200),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_724),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_607),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_83),
.Y(n_1106)
);

CKINVDCx16_ASAP7_75t_R g1107 ( 
.A(n_371),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_308),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_408),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_37),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_299),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_671),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_75),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_592),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_794),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_516),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_735),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_616),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_710),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_716),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_327),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_748),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_343),
.Y(n_1123)
);

BUFx10_ASAP7_75t_L g1124 ( 
.A(n_687),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_308),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_758),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_334),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_442),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_803),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_413),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_38),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_213),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_153),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_727),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_583),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_36),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_219),
.Y(n_1137)
);

CKINVDCx16_ASAP7_75t_R g1138 ( 
.A(n_710),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_641),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_206),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_178),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_754),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_286),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_348),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_99),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_290),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_386),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_210),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_157),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_375),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_116),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_607),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_30),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_460),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_436),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_47),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_686),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_333),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_288),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_745),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_141),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_458),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_35),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_725),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_661),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_142),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_753),
.Y(n_1167)
);

BUFx10_ASAP7_75t_L g1168 ( 
.A(n_622),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_362),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_201),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_370),
.Y(n_1171)
);

BUFx10_ASAP7_75t_L g1172 ( 
.A(n_216),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_615),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_696),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_169),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_767),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_448),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_260),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_270),
.Y(n_1179)
);

BUFx8_ASAP7_75t_SL g1180 ( 
.A(n_322),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_390),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_717),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_278),
.Y(n_1183)
);

BUFx10_ASAP7_75t_L g1184 ( 
.A(n_282),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_276),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_516),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_506),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_445),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_732),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_118),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_150),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_368),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_357),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_478),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_769),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_656),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_514),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_417),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_767),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_54),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_808),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_134),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_578),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_273),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_333),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_614),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_98),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_650),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_280),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_476),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_809),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_400),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_140),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_145),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_798),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_729),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_158),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_112),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_713),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_156),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_783),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_691),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_467),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_714),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_388),
.Y(n_1225)
);

BUFx5_ASAP7_75t_L g1226 ( 
.A(n_517),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_729),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_296),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_302),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_94),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_139),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_430),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_119),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_213),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_360),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_593),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_682),
.Y(n_1237)
);

BUFx10_ASAP7_75t_L g1238 ( 
.A(n_733),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_396),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_34),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_343),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_799),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_10),
.Y(n_1243)
);

CKINVDCx16_ASAP7_75t_R g1244 ( 
.A(n_737),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_57),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_294),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_167),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_205),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_385),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_706),
.Y(n_1250)
);

BUFx10_ASAP7_75t_L g1251 ( 
.A(n_499),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_741),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_94),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_461),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_187),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_692),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_487),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_481),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_773),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_148),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_373),
.Y(n_1261)
);

CKINVDCx16_ASAP7_75t_R g1262 ( 
.A(n_376),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_464),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_241),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_472),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_23),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_344),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_14),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_141),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_418),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_691),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_805),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_498),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_707),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_282),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_35),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_225),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_348),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_26),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_756),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_271),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_742),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_784),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_597),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_773),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_466),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_355),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_153),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_750),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_537),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_452),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_731),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_797),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_550),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_746),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_667),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_126),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_184),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_475),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_83),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_195),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_332),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_701),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_359),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_134),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_554),
.Y(n_1306)
);

CKINVDCx16_ASAP7_75t_R g1307 ( 
.A(n_411),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_182),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_264),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_353),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_721),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_740),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_235),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_647),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_588),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_763),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_162),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_219),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_472),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_488),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_306),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_636),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_191),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_549),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_121),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_209),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_580),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_350),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_262),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_312),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_11),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_483),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_33),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_731),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_405),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_680),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_227),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_667),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_454),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_688),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_248),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_20),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_492),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_285),
.Y(n_1344)
);

BUFx10_ASAP7_75t_L g1345 ( 
.A(n_719),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_629),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_923),
.Y(n_1347)
);

INVxp33_ASAP7_75t_L g1348 ( 
.A(n_1054),
.Y(n_1348)
);

CKINVDCx16_ASAP7_75t_R g1349 ( 
.A(n_1002),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_836),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_893),
.B(n_0),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1180),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_836),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_836),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_836),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_836),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_836),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_836),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_985),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_848),
.Y(n_1360)
);

INVxp67_ASAP7_75t_SL g1361 ( 
.A(n_1242),
.Y(n_1361)
);

INVxp67_ASAP7_75t_L g1362 ( 
.A(n_942),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1035),
.Y(n_1363)
);

INVxp33_ASAP7_75t_SL g1364 ( 
.A(n_1291),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1115),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_848),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_848),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_848),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_848),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_857),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_848),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_848),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_955),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_955),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_955),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_955),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_1024),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1201),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_954),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1211),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1215),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_857),
.B(n_0),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_955),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_955),
.Y(n_1384)
);

INVxp67_ASAP7_75t_SL g1385 ( 
.A(n_1242),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_955),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1073),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1079),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1073),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_1107),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1272),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1073),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1073),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1138),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1272),
.Y(n_1395)
);

INVxp33_ASAP7_75t_SL g1396 ( 
.A(n_811),
.Y(n_1396)
);

CKINVDCx16_ASAP7_75t_R g1397 ( 
.A(n_1244),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1073),
.Y(n_1398)
);

INVxp33_ASAP7_75t_L g1399 ( 
.A(n_1020),
.Y(n_1399)
);

INVxp33_ASAP7_75t_SL g1400 ( 
.A(n_811),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1073),
.Y(n_1401)
);

CKINVDCx16_ASAP7_75t_R g1402 ( 
.A(n_1262),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1307),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_838),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_821),
.Y(n_1405)
);

INVxp67_ASAP7_75t_SL g1406 ( 
.A(n_857),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1073),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1226),
.Y(n_1408)
);

CKINVDCx16_ASAP7_75t_R g1409 ( 
.A(n_826),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1226),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1226),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1226),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1226),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_812),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1226),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1226),
.Y(n_1416)
);

CKINVDCx14_ASAP7_75t_R g1417 ( 
.A(n_1050),
.Y(n_1417)
);

INVxp33_ASAP7_75t_L g1418 ( 
.A(n_1276),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_902),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_821),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_857),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_885),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_902),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_905),
.Y(n_1424)
);

INVxp33_ASAP7_75t_L g1425 ( 
.A(n_1297),
.Y(n_1425)
);

INVxp33_ASAP7_75t_L g1426 ( 
.A(n_827),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_905),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_916),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1293),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_916),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_918),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_918),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_916),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_814),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_885),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_935),
.Y(n_1436)
);

INVxp67_ASAP7_75t_SL g1437 ( 
.A(n_916),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_949),
.B(n_1),
.Y(n_1438)
);

INVxp67_ASAP7_75t_SL g1439 ( 
.A(n_949),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_826),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_949),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_819),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_935),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_938),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_938),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1006),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1006),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1089),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_826),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1089),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1105),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1105),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1185),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_949),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1185),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1188),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_896),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_822),
.Y(n_1458)
);

INVxp33_ASAP7_75t_SL g1459 ( 
.A(n_824),
.Y(n_1459)
);

INVxp33_ASAP7_75t_L g1460 ( 
.A(n_827),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_959),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1188),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1209),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1209),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1255),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1255),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_828),
.Y(n_1467)
);

INVxp33_ASAP7_75t_SL g1468 ( 
.A(n_824),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_830),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1260),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_959),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1260),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1261),
.Y(n_1473)
);

CKINVDCx16_ASAP7_75t_R g1474 ( 
.A(n_936),
.Y(n_1474)
);

CKINVDCx16_ASAP7_75t_R g1475 ( 
.A(n_936),
.Y(n_1475)
);

INVxp67_ASAP7_75t_SL g1476 ( 
.A(n_959),
.Y(n_1476)
);

CKINVDCx14_ASAP7_75t_R g1477 ( 
.A(n_959),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_896),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1261),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1284),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1284),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1343),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1343),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_962),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_936),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_962),
.Y(n_1486)
);

NOR2xp67_ASAP7_75t_L g1487 ( 
.A(n_1016),
.B(n_1),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1352),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1429),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1421),
.Y(n_1490)
);

BUFx8_ASAP7_75t_L g1491 ( 
.A(n_1419),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1359),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1350),
.A2(n_1293),
.B(n_1129),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1363),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1365),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1421),
.Y(n_1496)
);

BUFx8_ASAP7_75t_SL g1497 ( 
.A(n_1405),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_1429),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1429),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1361),
.B(n_823),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1429),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1440),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1428),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1406),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1428),
.Y(n_1505)
);

CKINVDCx11_ASAP7_75t_R g1506 ( 
.A(n_1420),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1430),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1430),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1437),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1477),
.B(n_962),
.Y(n_1510)
);

BUFx12f_ASAP7_75t_L g1511 ( 
.A(n_1388),
.Y(n_1511)
);

BUFx8_ASAP7_75t_L g1512 ( 
.A(n_1423),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1433),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1370),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1433),
.Y(n_1515)
);

CKINVDCx11_ASAP7_75t_R g1516 ( 
.A(n_1422),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1439),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1454),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1441),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_1378),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1347),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1441),
.Y(n_1522)
);

BUFx12f_ASAP7_75t_L g1523 ( 
.A(n_1390),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1414),
.B(n_838),
.Y(n_1524)
);

INVx6_ASAP7_75t_L g1525 ( 
.A(n_1409),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1385),
.B(n_1477),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1461),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1380),
.B(n_1381),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1370),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1461),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1471),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1394),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1434),
.B(n_1000),
.Y(n_1533)
);

AOI22x1_ASAP7_75t_SL g1534 ( 
.A1(n_1435),
.A2(n_930),
.B1(n_932),
.B2(n_925),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1476),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1391),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1471),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1484),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1395),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1486),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1350),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1353),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1354),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1442),
.B(n_1000),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1355),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1356),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1354),
.Y(n_1547)
);

INVx5_ASAP7_75t_L g1548 ( 
.A(n_1474),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1458),
.B(n_851),
.Y(n_1549)
);

INVx4_ASAP7_75t_L g1550 ( 
.A(n_1467),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1469),
.B(n_962),
.Y(n_1551)
);

BUFx8_ASAP7_75t_L g1552 ( 
.A(n_1424),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1427),
.B(n_968),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1364),
.A2(n_850),
.B1(n_855),
.B2(n_825),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1376),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1362),
.B(n_968),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1396),
.B(n_851),
.Y(n_1557)
);

BUFx12f_ASAP7_75t_L g1558 ( 
.A(n_1403),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1376),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1431),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1379),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1357),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1358),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_SL g1564 ( 
.A(n_1377),
.B(n_925),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1360),
.Y(n_1565)
);

AOI22x1_ASAP7_75t_SL g1566 ( 
.A1(n_1457),
.A2(n_932),
.B1(n_944),
.B2(n_930),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1400),
.B(n_860),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1366),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1432),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1436),
.B(n_968),
.Y(n_1570)
);

BUFx8_ASAP7_75t_L g1571 ( 
.A(n_1443),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1417),
.B(n_1000),
.Y(n_1572)
);

BUFx8_ASAP7_75t_L g1573 ( 
.A(n_1444),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1445),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1446),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1367),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1349),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1368),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1369),
.Y(n_1579)
);

INVx6_ASAP7_75t_L g1580 ( 
.A(n_1475),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1371),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1397),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1372),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_L g1584 ( 
.A(n_1373),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1447),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1448),
.Y(n_1586)
);

OA21x2_ASAP7_75t_L g1587 ( 
.A1(n_1374),
.A2(n_926),
.B(n_917),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1450),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1375),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1383),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1417),
.A2(n_850),
.B1(n_855),
.B2(n_825),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1451),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1384),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1452),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1453),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1386),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1402),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1449),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1387),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1389),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1392),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1393),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1455),
.B(n_1456),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1398),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1401),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1407),
.Y(n_1606)
);

BUFx8_ASAP7_75t_SL g1607 ( 
.A(n_1478),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1462),
.B(n_968),
.Y(n_1608)
);

INVx5_ASAP7_75t_L g1609 ( 
.A(n_1426),
.Y(n_1609)
);

AOI22x1_ASAP7_75t_SL g1610 ( 
.A1(n_1463),
.A2(n_1336),
.B1(n_983),
.B2(n_992),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1426),
.B(n_1124),
.Y(n_1611)
);

AND2x2_ASAP7_75t_SL g1612 ( 
.A(n_1351),
.B(n_1382),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1408),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1521),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1569),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1489),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1489),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1503),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1574),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1583),
.B(n_1601),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1575),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1609),
.B(n_1399),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1585),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1489),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1609),
.B(n_1570),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1588),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_1561),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1592),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1609),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1594),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1498),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1595),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1503),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1583),
.B(n_1410),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1542),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1542),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1503),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1545),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1547),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1545),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1546),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1498),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1546),
.Y(n_1643)
);

BUFx6f_ASAP7_75t_L g1644 ( 
.A(n_1498),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1611),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1612),
.B(n_1459),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1562),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1562),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1565),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1502),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1565),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1541),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1593),
.Y(n_1653)
);

NAND3xp33_ASAP7_75t_L g1654 ( 
.A(n_1587),
.B(n_1438),
.C(n_1382),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1499),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1499),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1593),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1551),
.B(n_1468),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1513),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1563),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1499),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1513),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1563),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1497),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1563),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1555),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1557),
.A2(n_1485),
.B1(n_1399),
.B2(n_1425),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1577),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1513),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1515),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1578),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1578),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1578),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1601),
.B(n_1411),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1584),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1567),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1584),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1515),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1597),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1582),
.A2(n_983),
.B1(n_992),
.B2(n_944),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1510),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1584),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1501),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_SL g1684 ( 
.A1(n_1554),
.A2(n_1017),
.B1(n_1018),
.B2(n_994),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1589),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1589),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1589),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1590),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1526),
.B(n_1418),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1568),
.B(n_1412),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1590),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1590),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1596),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1515),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1556),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1596),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1519),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1576),
.B(n_1413),
.Y(n_1698)
);

XNOR2xp5_ASAP7_75t_L g1699 ( 
.A(n_1534),
.B(n_1418),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1572),
.B(n_1425),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1519),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1504),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1509),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1541),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1501),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1596),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1500),
.B(n_1415),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1602),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1519),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1602),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1522),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1533),
.B(n_1460),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1602),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1544),
.B(n_1524),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1501),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1522),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1605),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1522),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_1541),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1506),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1605),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1500),
.B(n_1416),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1605),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1527),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1613),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1527),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1598),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1613),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1548),
.B(n_1487),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1517),
.B(n_1348),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1549),
.B(n_1460),
.Y(n_1731)
);

OAI21x1_ASAP7_75t_L g1732 ( 
.A1(n_1493),
.A2(n_1465),
.B(n_1464),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1556),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1613),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1527),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1560),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1530),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1518),
.B(n_1348),
.Y(n_1738)
);

OAI21x1_ASAP7_75t_L g1739 ( 
.A1(n_1579),
.A2(n_1470),
.B(n_1466),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1530),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1581),
.Y(n_1741)
);

BUFx6f_ASAP7_75t_L g1742 ( 
.A(n_1543),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1516),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1570),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1548),
.B(n_1052),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1599),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1600),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1530),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1604),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1543),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1639),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1627),
.B(n_1548),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1639),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1739),
.Y(n_1754)
);

AND2x6_ASAP7_75t_L g1755 ( 
.A(n_1714),
.B(n_1528),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1731),
.B(n_1550),
.Y(n_1756)
);

INVx4_ASAP7_75t_L g1757 ( 
.A(n_1719),
.Y(n_1757)
);

AO22x2_ASAP7_75t_L g1758 ( 
.A1(n_1676),
.A2(n_1610),
.B1(n_1566),
.B2(n_1534),
.Y(n_1758)
);

INVx4_ASAP7_75t_L g1759 ( 
.A(n_1719),
.Y(n_1759)
);

BUFx10_ASAP7_75t_L g1760 ( 
.A(n_1664),
.Y(n_1760)
);

OR2x6_ASAP7_75t_L g1761 ( 
.A(n_1614),
.B(n_1650),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1627),
.B(n_1550),
.Y(n_1762)
);

OR2x6_ASAP7_75t_L g1763 ( 
.A(n_1668),
.B(n_1525),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1664),
.Y(n_1764)
);

INVx5_ASAP7_75t_L g1765 ( 
.A(n_1616),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1744),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1654),
.A2(n_1587),
.B1(n_1606),
.B2(n_1535),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1744),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1645),
.A2(n_1520),
.B1(n_1494),
.B2(n_1495),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1615),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1720),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1619),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1666),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1679),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1666),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1712),
.B(n_1492),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1689),
.B(n_1492),
.Y(n_1777)
);

INVx5_ASAP7_75t_L g1778 ( 
.A(n_1616),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1700),
.B(n_1495),
.Y(n_1779)
);

INVx1_ASAP7_75t_SL g1780 ( 
.A(n_1727),
.Y(n_1780)
);

BUFx3_ASAP7_75t_L g1781 ( 
.A(n_1736),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1621),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1741),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1623),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1626),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1746),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1681),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1676),
.B(n_1532),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1681),
.B(n_1543),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1645),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1720),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1628),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1658),
.B(n_1625),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1658),
.B(n_1559),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1646),
.B(n_1525),
.Y(n_1795)
);

CKINVDCx20_ASAP7_75t_R g1796 ( 
.A(n_1743),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1747),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1622),
.B(n_1738),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1749),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1654),
.A2(n_1438),
.B1(n_1559),
.B2(n_1608),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1635),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1730),
.B(n_1586),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_1743),
.Y(n_1803)
);

INVx3_ASAP7_75t_L g1804 ( 
.A(n_1719),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1742),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1636),
.A2(n_1559),
.B1(n_1608),
.B2(n_1053),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1625),
.B(n_1564),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1630),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1632),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1646),
.B(n_1580),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1702),
.B(n_1514),
.Y(n_1811)
);

INVx2_ASAP7_75t_SL g1812 ( 
.A(n_1629),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1638),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1640),
.Y(n_1814)
);

AND3x1_ASAP7_75t_L g1815 ( 
.A(n_1667),
.B(n_1473),
.C(n_1472),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1641),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1643),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1647),
.B(n_1537),
.Y(n_1818)
);

BUFx10_ASAP7_75t_L g1819 ( 
.A(n_1730),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1629),
.B(n_1580),
.Y(n_1820)
);

BUFx3_ASAP7_75t_L g1821 ( 
.A(n_1702),
.Y(n_1821)
);

AOI21x1_ASAP7_75t_L g1822 ( 
.A1(n_1620),
.A2(n_1496),
.B(n_1490),
.Y(n_1822)
);

BUFx3_ASAP7_75t_L g1823 ( 
.A(n_1703),
.Y(n_1823)
);

INVxp33_ASAP7_75t_L g1824 ( 
.A(n_1680),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1648),
.A2(n_1053),
.B1(n_1117),
.B2(n_1052),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1649),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1695),
.B(n_1591),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1651),
.B(n_1537),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1703),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1653),
.Y(n_1830)
);

OR2x6_ASAP7_75t_L g1831 ( 
.A(n_1684),
.B(n_1511),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1657),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_1745),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1620),
.B(n_1537),
.Y(n_1834)
);

INVxp33_ASAP7_75t_L g1835 ( 
.A(n_1699),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1695),
.Y(n_1836)
);

AND2x6_ASAP7_75t_L g1837 ( 
.A(n_1704),
.B(n_1750),
.Y(n_1837)
);

AND3x2_ASAP7_75t_L g1838 ( 
.A(n_1733),
.B(n_1539),
.C(n_1536),
.Y(n_1838)
);

BUFx3_ASAP7_75t_L g1839 ( 
.A(n_1733),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1707),
.A2(n_1053),
.B1(n_1117),
.B2(n_1052),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1732),
.Y(n_1841)
);

OAI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1707),
.A2(n_818),
.B1(n_852),
.B2(n_816),
.Y(n_1842)
);

INVx4_ASAP7_75t_L g1843 ( 
.A(n_1742),
.Y(n_1843)
);

BUFx10_ASAP7_75t_L g1844 ( 
.A(n_1660),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1690),
.Y(n_1845)
);

NAND3xp33_ASAP7_75t_L g1846 ( 
.A(n_1722),
.B(n_1603),
.C(n_1480),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1722),
.B(n_1404),
.Y(n_1847)
);

OAI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1634),
.A2(n_1674),
.B1(n_1698),
.B2(n_1690),
.Y(n_1848)
);

NAND2xp33_ASAP7_75t_L g1849 ( 
.A(n_1704),
.B(n_1750),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1663),
.B(n_1505),
.Y(n_1850)
);

BUFx3_ASAP7_75t_L g1851 ( 
.A(n_1618),
.Y(n_1851)
);

NAND2xp33_ASAP7_75t_L g1852 ( 
.A(n_1633),
.B(n_1052),
.Y(n_1852)
);

BUFx4f_ASAP7_75t_L g1853 ( 
.A(n_1665),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1671),
.B(n_1507),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1745),
.B(n_1523),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1698),
.Y(n_1856)
);

AO22x2_ASAP7_75t_L g1857 ( 
.A1(n_1729),
.A2(n_1610),
.B1(n_1566),
.B2(n_933),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1634),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1729),
.B(n_1404),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1674),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_SL g1861 ( 
.A(n_1672),
.B(n_1488),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1637),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1673),
.B(n_1479),
.Y(n_1863)
);

OR2x6_ASAP7_75t_L g1864 ( 
.A(n_1659),
.B(n_1558),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_SL g1865 ( 
.A(n_1742),
.B(n_1514),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_SL g1866 ( 
.A1(n_1675),
.A2(n_1017),
.B1(n_1018),
.B2(n_994),
.Y(n_1866)
);

INVx4_ASAP7_75t_SL g1867 ( 
.A(n_1616),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1677),
.B(n_1508),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1662),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1682),
.B(n_1538),
.Y(n_1870)
);

INVx4_ASAP7_75t_L g1871 ( 
.A(n_1624),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1669),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1685),
.B(n_1529),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1686),
.A2(n_1553),
.B1(n_1529),
.B2(n_1540),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1687),
.B(n_1481),
.Y(n_1875)
);

OR2x6_ASAP7_75t_L g1876 ( 
.A(n_1670),
.B(n_860),
.Y(n_1876)
);

AND2x2_ASAP7_75t_SL g1877 ( 
.A(n_1678),
.B(n_846),
.Y(n_1877)
);

OAI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1688),
.A2(n_853),
.B1(n_871),
.B2(n_854),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1691),
.B(n_1607),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1694),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1697),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1701),
.Y(n_1882)
);

INVx4_ASAP7_75t_L g1883 ( 
.A(n_1624),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1692),
.B(n_1053),
.Y(n_1884)
);

NAND2xp33_ASAP7_75t_L g1885 ( 
.A(n_1709),
.B(n_1737),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1693),
.B(n_1696),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1706),
.B(n_1538),
.Y(n_1887)
);

BUFx4f_ASAP7_75t_L g1888 ( 
.A(n_1708),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1710),
.B(n_875),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1711),
.Y(n_1890)
);

BUFx3_ASAP7_75t_L g1891 ( 
.A(n_1718),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1726),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1713),
.B(n_1117),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1740),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1748),
.Y(n_1895)
);

INVx4_ASAP7_75t_L g1896 ( 
.A(n_1624),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1717),
.B(n_909),
.Y(n_1897)
);

OR2x6_ASAP7_75t_L g1898 ( 
.A(n_1721),
.B(n_933),
.Y(n_1898)
);

NOR2x1p5_ASAP7_75t_L g1899 ( 
.A(n_1723),
.B(n_856),
.Y(n_1899)
);

INVx2_ASAP7_75t_SL g1900 ( 
.A(n_1617),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1725),
.B(n_1540),
.Y(n_1901)
);

INVx3_ASAP7_75t_L g1902 ( 
.A(n_1716),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1728),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1734),
.A2(n_1191),
.B1(n_1231),
.B2(n_1117),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1716),
.B(n_1482),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1617),
.Y(n_1906)
);

INVx5_ASAP7_75t_L g1907 ( 
.A(n_1631),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1661),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1652),
.B(n_1531),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1724),
.Y(n_1910)
);

AND2x6_ASAP7_75t_L g1911 ( 
.A(n_1724),
.B(n_846),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1788),
.B(n_1652),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1756),
.B(n_1631),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1845),
.B(n_1856),
.Y(n_1914)
);

INVx8_ASAP7_75t_L g1915 ( 
.A(n_1763),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1816),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1858),
.B(n_1735),
.Y(n_1917)
);

AOI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1755),
.A2(n_1735),
.B1(n_1661),
.B2(n_1642),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1817),
.Y(n_1919)
);

AOI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1860),
.A2(n_1231),
.B1(n_1236),
.B2(n_1191),
.Y(n_1920)
);

NAND2xp33_ASAP7_75t_L g1921 ( 
.A(n_1755),
.B(n_1631),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1751),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1777),
.B(n_1642),
.Y(n_1923)
);

INVx2_ASAP7_75t_SL g1924 ( 
.A(n_1774),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1794),
.B(n_1642),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1780),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1819),
.B(n_1787),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1802),
.B(n_1644),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1798),
.B(n_1644),
.Y(n_1929)
);

NOR2x2_ASAP7_75t_L g1930 ( 
.A(n_1761),
.B(n_1831),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1753),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1773),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1789),
.B(n_1644),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1819),
.B(n_1779),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1755),
.B(n_1848),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1755),
.B(n_1655),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1847),
.B(n_1655),
.Y(n_1937)
);

O2A1O1Ixp5_ASAP7_75t_L g1938 ( 
.A1(n_1822),
.A2(n_914),
.B(n_941),
.C(n_882),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1821),
.B(n_1655),
.Y(n_1939)
);

AOI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1827),
.A2(n_1034),
.B1(n_1078),
.B2(n_1042),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1801),
.B(n_1656),
.Y(n_1941)
);

AOI22xp33_ASAP7_75t_L g1942 ( 
.A1(n_1800),
.A2(n_1231),
.B1(n_1236),
.B2(n_1191),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1813),
.B(n_1656),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1775),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1814),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1766),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_SL g1947 ( 
.A(n_1823),
.B(n_1656),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1826),
.B(n_1683),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1834),
.A2(n_1705),
.B(n_1683),
.Y(n_1949)
);

AO221x1_ASAP7_75t_L g1950 ( 
.A1(n_1758),
.A2(n_1236),
.B1(n_1290),
.B2(n_1231),
.C(n_1191),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_SL g1951 ( 
.A(n_1829),
.B(n_1683),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1830),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1768),
.Y(n_1953)
);

INVx4_ASAP7_75t_L g1954 ( 
.A(n_1867),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1811),
.B(n_1705),
.Y(n_1955)
);

NOR2xp33_ASAP7_75t_L g1956 ( 
.A(n_1790),
.B(n_1034),
.Y(n_1956)
);

BUFx5_ASAP7_75t_L g1957 ( 
.A(n_1841),
.Y(n_1957)
);

AND2x6_ASAP7_75t_SL g1958 ( 
.A(n_1831),
.B(n_1344),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1770),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1832),
.B(n_1705),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1772),
.B(n_1715),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_SL g1962 ( 
.A(n_1764),
.B(n_1042),
.Y(n_1962)
);

NAND2xp33_ASAP7_75t_L g1963 ( 
.A(n_1911),
.B(n_1715),
.Y(n_1963)
);

NOR3xp33_ASAP7_75t_L g1964 ( 
.A(n_1795),
.B(n_1483),
.C(n_961),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1782),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1859),
.B(n_1124),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1793),
.B(n_1078),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1839),
.B(n_1101),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1767),
.A2(n_1849),
.B(n_1909),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1784),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1910),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1785),
.B(n_1715),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1792),
.B(n_1531),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1910),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1808),
.B(n_1809),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1877),
.B(n_984),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1905),
.B(n_984),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1811),
.B(n_1571),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1783),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1836),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1889),
.B(n_1897),
.Y(n_1981)
);

AND2x2_ASAP7_75t_SL g1982 ( 
.A(n_1861),
.B(n_882),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1833),
.B(n_1068),
.Y(n_1983)
);

INVx2_ASAP7_75t_SL g1984 ( 
.A(n_1761),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1894),
.B(n_1068),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_SL g1986 ( 
.A(n_1769),
.B(n_1491),
.Y(n_1986)
);

AOI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1842),
.A2(n_1290),
.B1(n_1321),
.B2(n_1236),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1812),
.B(n_1491),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1786),
.Y(n_1989)
);

INVxp67_ASAP7_75t_L g1990 ( 
.A(n_1815),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1797),
.B(n_1258),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1875),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1810),
.B(n_1101),
.Y(n_1993)
);

NAND2xp33_ASAP7_75t_L g1994 ( 
.A(n_1911),
.B(n_1290),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1799),
.B(n_1902),
.Y(n_1995)
);

NAND2xp33_ASAP7_75t_L g1996 ( 
.A(n_1911),
.B(n_1837),
.Y(n_1996)
);

A2O1A1Ixp33_ASAP7_75t_L g1997 ( 
.A1(n_1853),
.A2(n_1283),
.B(n_1346),
.C(n_1258),
.Y(n_1997)
);

NAND2x1_ASAP7_75t_L g1998 ( 
.A(n_1837),
.B(n_1290),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1875),
.Y(n_1999)
);

NOR3xp33_ASAP7_75t_L g2000 ( 
.A(n_1807),
.B(n_1062),
.C(n_912),
.Y(n_2000)
);

AOI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1758),
.A2(n_1109),
.B1(n_1147),
.B2(n_1131),
.Y(n_2001)
);

AOI22x1_ASAP7_75t_L g2002 ( 
.A1(n_1892),
.A2(n_1283),
.B1(n_1346),
.B2(n_858),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1902),
.B(n_1321),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1863),
.Y(n_2004)
);

NAND2x1_ASAP7_75t_L g2005 ( 
.A(n_1837),
.B(n_1321),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1850),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1892),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1804),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1886),
.B(n_1321),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1854),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1868),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1853),
.B(n_1888),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1804),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1805),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1824),
.B(n_1109),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1888),
.B(n_1512),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1818),
.B(n_832),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1776),
.B(n_1820),
.Y(n_2018)
);

AOI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_1857),
.A2(n_1911),
.B1(n_1846),
.B2(n_1866),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1805),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1903),
.Y(n_2021)
);

BUFx2_ASAP7_75t_L g2022 ( 
.A(n_1763),
.Y(n_2022)
);

NAND2xp33_ASAP7_75t_L g2023 ( 
.A(n_1837),
.B(n_837),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1828),
.B(n_840),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1870),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1851),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1762),
.B(n_1855),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1781),
.B(n_1571),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1765),
.B(n_1573),
.Y(n_2029)
);

NAND2xp33_ASAP7_75t_SL g2030 ( 
.A(n_1899),
.B(n_1131),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1887),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_R g2032 ( 
.A(n_1803),
.B(n_1512),
.Y(n_2032)
);

O2A1O1Ixp33_ASAP7_75t_L g2033 ( 
.A1(n_1884),
.A2(n_1163),
.B(n_1216),
.C(n_1102),
.Y(n_2033)
);

OR2x2_ASAP7_75t_L g2034 ( 
.A(n_1791),
.B(n_1229),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1900),
.B(n_841),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1898),
.B(n_1124),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1765),
.B(n_1573),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1862),
.B(n_845),
.Y(n_2038)
);

NOR2x1_ASAP7_75t_L g2039 ( 
.A(n_1879),
.B(n_1147),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1857),
.A2(n_1232),
.B1(n_1235),
.B2(n_1199),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1869),
.B(n_849),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1901),
.Y(n_2042)
);

O2A1O1Ixp5_ASAP7_75t_L g2043 ( 
.A1(n_1873),
.A2(n_941),
.B(n_1014),
.C(n_914),
.Y(n_2043)
);

AOI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1872),
.A2(n_1232),
.B1(n_1235),
.B2(n_1199),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1765),
.B(n_1552),
.Y(n_2045)
);

AOI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_1840),
.A2(n_1266),
.B1(n_1277),
.B2(n_1265),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1880),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1778),
.B(n_1552),
.Y(n_2048)
);

BUFx6f_ASAP7_75t_L g2049 ( 
.A(n_1778),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1881),
.B(n_889),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1882),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1891),
.Y(n_2052)
);

BUFx3_ASAP7_75t_L g2053 ( 
.A(n_1796),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1752),
.B(n_1265),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1890),
.B(n_890),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1895),
.B(n_891),
.Y(n_2056)
);

INVx5_ASAP7_75t_L g2057 ( 
.A(n_1864),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1906),
.B(n_892),
.Y(n_2058)
);

INVx2_ASAP7_75t_SL g2059 ( 
.A(n_1876),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1908),
.Y(n_2060)
);

NOR2xp67_ASAP7_75t_L g2061 ( 
.A(n_1874),
.B(n_1865),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1778),
.B(n_1266),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1754),
.Y(n_2063)
);

OAI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_1898),
.A2(n_1336),
.B1(n_1294),
.B2(n_1314),
.Y(n_2064)
);

AND2x4_ASAP7_75t_SL g2065 ( 
.A(n_1760),
.B(n_1168),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1907),
.B(n_1277),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_SL g2067 ( 
.A(n_1907),
.B(n_1294),
.Y(n_2067)
);

NAND2xp33_ASAP7_75t_L g2068 ( 
.A(n_1754),
.B(n_894),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_1771),
.B(n_1279),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1757),
.B(n_895),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1867),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1907),
.B(n_1757),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_1878),
.A2(n_1316),
.B1(n_1317),
.B2(n_1314),
.Y(n_2073)
);

NOR2xp33_ASAP7_75t_L g2074 ( 
.A(n_1844),
.B(n_1835),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1759),
.B(n_899),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1759),
.B(n_900),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1843),
.B(n_903),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1843),
.B(n_910),
.Y(n_2078)
);

INVx2_ASAP7_75t_SL g2079 ( 
.A(n_1876),
.Y(n_2079)
);

NAND3x1_ASAP7_75t_L g2080 ( 
.A(n_1760),
.B(n_843),
.C(n_820),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1871),
.B(n_1883),
.Y(n_2081)
);

INVxp67_ASAP7_75t_L g2082 ( 
.A(n_1864),
.Y(n_2082)
);

O2A1O1Ixp33_ASAP7_75t_L g2083 ( 
.A1(n_1893),
.A2(n_1339),
.B(n_1019),
.C(n_1032),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1844),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1754),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1916),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1919),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1971),
.Y(n_2088)
);

AO22x1_ASAP7_75t_L g2089 ( 
.A1(n_1993),
.A2(n_858),
.B1(n_861),
.B2(n_856),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1959),
.Y(n_2090)
);

AOI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_1981),
.A2(n_1885),
.B1(n_1871),
.B2(n_1883),
.Y(n_2091)
);

BUFx3_ASAP7_75t_L g2092 ( 
.A(n_1915),
.Y(n_2092)
);

AND2x6_ASAP7_75t_L g2093 ( 
.A(n_1935),
.B(n_1014),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1914),
.B(n_1912),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1974),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2007),
.Y(n_2096)
);

INVx2_ASAP7_75t_SL g2097 ( 
.A(n_1926),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2006),
.B(n_2010),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2011),
.B(n_1806),
.Y(n_2099)
);

NAND3xp33_ASAP7_75t_SL g2100 ( 
.A(n_1940),
.B(n_1317),
.C(n_1316),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1928),
.B(n_1896),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1934),
.B(n_1896),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1965),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2025),
.B(n_1825),
.Y(n_2104)
);

INVxp67_ASAP7_75t_SL g2105 ( 
.A(n_1937),
.Y(n_2105)
);

INVx2_ASAP7_75t_SL g2106 ( 
.A(n_1915),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_R g2107 ( 
.A(n_2030),
.B(n_1924),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_R g2108 ( 
.A(n_1915),
.B(n_1838),
.Y(n_2108)
);

AND2x6_ASAP7_75t_L g2109 ( 
.A(n_2063),
.B(n_1019),
.Y(n_2109)
);

O2A1O1Ixp33_ASAP7_75t_L g2110 ( 
.A1(n_1997),
.A2(n_1852),
.B(n_815),
.C(n_817),
.Y(n_2110)
);

OAI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_2027),
.A2(n_1904),
.B1(n_1320),
.B2(n_1332),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2031),
.B(n_2042),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1970),
.Y(n_2113)
);

BUFx3_ASAP7_75t_L g2114 ( 
.A(n_2022),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1975),
.B(n_911),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_2069),
.B(n_861),
.Y(n_2116)
);

AOI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_1969),
.A2(n_829),
.B(n_813),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1946),
.Y(n_2118)
);

INVx5_ASAP7_75t_L g2119 ( 
.A(n_1954),
.Y(n_2119)
);

AND2x4_ASAP7_75t_SL g2120 ( 
.A(n_1954),
.B(n_1168),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1922),
.Y(n_2121)
);

HB1xp67_ASAP7_75t_L g2122 ( 
.A(n_2053),
.Y(n_2122)
);

AOI21xp5_ASAP7_75t_L g2123 ( 
.A1(n_1994),
.A2(n_833),
.B(n_831),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1953),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1931),
.Y(n_2125)
);

INVx2_ASAP7_75t_SL g2126 ( 
.A(n_2034),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1980),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_1982),
.B(n_1318),
.Y(n_2128)
);

INVx2_ASAP7_75t_SL g2129 ( 
.A(n_2059),
.Y(n_2129)
);

INVxp67_ASAP7_75t_SL g2130 ( 
.A(n_1929),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_1999),
.B(n_834),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_L g2132 ( 
.A(n_2015),
.B(n_1318),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1966),
.B(n_913),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1932),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1944),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_1967),
.B(n_1320),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2047),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_2049),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2004),
.B(n_921),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_2049),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1977),
.B(n_922),
.Y(n_2141)
);

BUFx8_ASAP7_75t_L g2142 ( 
.A(n_1984),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_SL g2143 ( 
.A(n_2019),
.B(n_1332),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2018),
.A2(n_927),
.B1(n_928),
.B2(n_924),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2051),
.Y(n_2145)
);

HB1xp67_ASAP7_75t_L g2146 ( 
.A(n_1990),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1945),
.B(n_929),
.Y(n_2147)
);

A2O1A1Ixp33_ASAP7_75t_L g2148 ( 
.A1(n_2019),
.A2(n_839),
.B(n_842),
.C(n_835),
.Y(n_2148)
);

NOR2xp33_ASAP7_75t_L g2149 ( 
.A(n_1927),
.B(n_934),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1952),
.B(n_937),
.Y(n_2150)
);

O2A1O1Ixp33_ASAP7_75t_L g2151 ( 
.A1(n_1976),
.A2(n_1983),
.B(n_1964),
.C(n_2012),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2021),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1979),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1989),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_1956),
.B(n_1940),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_SL g2156 ( 
.A(n_2026),
.B(n_939),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_2060),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1917),
.Y(n_2158)
);

OAI21xp5_ASAP7_75t_L g2159 ( 
.A1(n_1938),
.A2(n_847),
.B(n_844),
.Y(n_2159)
);

OR2x2_ASAP7_75t_SL g2160 ( 
.A(n_2084),
.B(n_1032),
.Y(n_2160)
);

BUFx3_ASAP7_75t_L g2161 ( 
.A(n_2057),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1933),
.B(n_940),
.Y(n_2162)
);

AND3x2_ASAP7_75t_SL g2163 ( 
.A(n_2073),
.B(n_1047),
.C(n_1037),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_2052),
.B(n_945),
.Y(n_2164)
);

BUFx6f_ASAP7_75t_L g2165 ( 
.A(n_2049),
.Y(n_2165)
);

AND2x4_ASAP7_75t_L g2166 ( 
.A(n_1992),
.B(n_859),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2017),
.B(n_946),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_L g2168 ( 
.A(n_1968),
.B(n_947),
.Y(n_2168)
);

A2O1A1Ixp33_ASAP7_75t_L g2169 ( 
.A1(n_2061),
.A2(n_865),
.B(n_869),
.C(n_862),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1991),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_2008),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2013),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1973),
.Y(n_2173)
);

NAND3xp33_ASAP7_75t_SL g2174 ( 
.A(n_1962),
.B(n_864),
.C(n_863),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2014),
.Y(n_2175)
);

INVx5_ASAP7_75t_L g2176 ( 
.A(n_2057),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_2062),
.B(n_948),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1995),
.Y(n_2178)
);

AOI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_2000),
.A2(n_953),
.B1(n_958),
.B2(n_951),
.Y(n_2179)
);

AOI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2039),
.A2(n_963),
.B1(n_965),
.B2(n_960),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2024),
.B(n_967),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1925),
.B(n_970),
.Y(n_2182)
);

BUFx6f_ASAP7_75t_L g2183 ( 
.A(n_2071),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_2020),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1961),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1972),
.Y(n_2186)
);

AOI22xp33_ASAP7_75t_SL g2187 ( 
.A1(n_2054),
.A2(n_1345),
.B1(n_1251),
.B2(n_1172),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_1985),
.B(n_2044),
.Y(n_2188)
);

INVxp33_ASAP7_75t_L g2189 ( 
.A(n_2074),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1941),
.Y(n_2190)
);

NOR2x2_ASAP7_75t_L g2191 ( 
.A(n_2073),
.B(n_1037),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_2057),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1943),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2085),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1942),
.B(n_971),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1948),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2070),
.B(n_974),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1960),
.Y(n_2198)
);

NAND2x1p5_ASAP7_75t_L g2199 ( 
.A(n_2072),
.B(n_870),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2003),
.Y(n_2200)
);

INVx2_ASAP7_75t_SL g2201 ( 
.A(n_2079),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1955),
.Y(n_2202)
);

OAI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_2046),
.A2(n_976),
.B1(n_977),
.B2(n_975),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2043),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_SL g2205 ( 
.A(n_2075),
.B(n_2076),
.Y(n_2205)
);

INVxp67_ASAP7_75t_L g2206 ( 
.A(n_2036),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1957),
.Y(n_2207)
);

INVx4_ASAP7_75t_L g2208 ( 
.A(n_2065),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2038),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2041),
.Y(n_2210)
);

BUFx6f_ASAP7_75t_L g2211 ( 
.A(n_1936),
.Y(n_2211)
);

O2A1O1Ixp33_ASAP7_75t_L g2212 ( 
.A1(n_2058),
.A2(n_881),
.B(n_883),
.C(n_880),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2050),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_2032),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2077),
.B(n_978),
.Y(n_2215)
);

BUFx3_ASAP7_75t_L g2216 ( 
.A(n_2035),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_2066),
.B(n_2067),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2078),
.B(n_980),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1913),
.B(n_981),
.Y(n_2219)
);

INVxp67_ASAP7_75t_SL g2220 ( 
.A(n_2081),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2055),
.Y(n_2221)
);

OR2x2_ASAP7_75t_L g2222 ( 
.A(n_2056),
.B(n_863),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1957),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1957),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1957),
.Y(n_2225)
);

NOR2xp33_ASAP7_75t_L g2226 ( 
.A(n_2064),
.B(n_987),
.Y(n_2226)
);

O2A1O1Ixp5_ASAP7_75t_L g2227 ( 
.A1(n_1998),
.A2(n_1058),
.B(n_1064),
.C(n_1047),
.Y(n_2227)
);

OAI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2046),
.A2(n_990),
.B1(n_991),
.B2(n_988),
.Y(n_2228)
);

INVx1_ASAP7_75t_SL g2229 ( 
.A(n_1930),
.Y(n_2229)
);

BUFx3_ASAP7_75t_L g2230 ( 
.A(n_2040),
.Y(n_2230)
);

OR2x2_ASAP7_75t_L g2231 ( 
.A(n_1939),
.B(n_864),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1923),
.B(n_993),
.Y(n_2232)
);

AOI22xp33_ASAP7_75t_SL g2233 ( 
.A1(n_2002),
.A2(n_1238),
.B1(n_1172),
.B2(n_1184),
.Y(n_2233)
);

INVx4_ASAP7_75t_L g2234 ( 
.A(n_1958),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1987),
.B(n_996),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2009),
.Y(n_2236)
);

INVx3_ASAP7_75t_L g2237 ( 
.A(n_2080),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_1947),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1920),
.B(n_997),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_SL g2240 ( 
.A(n_2126),
.B(n_2040),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_2097),
.B(n_2001),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_2094),
.B(n_2001),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_2098),
.B(n_1988),
.Y(n_2243)
);

NAND2xp33_ASAP7_75t_SL g2244 ( 
.A(n_2107),
.B(n_1986),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_2155),
.B(n_2016),
.Y(n_2245)
);

NAND2xp33_ASAP7_75t_SL g2246 ( 
.A(n_2140),
.B(n_1978),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_SL g2247 ( 
.A(n_2189),
.B(n_2082),
.Y(n_2247)
);

NAND2xp33_ASAP7_75t_SL g2248 ( 
.A(n_2140),
.B(n_2029),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2112),
.B(n_2068),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_SL g2250 ( 
.A(n_2136),
.B(n_2028),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_2217),
.B(n_2188),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_2176),
.B(n_2037),
.Y(n_2252)
);

NAND2xp33_ASAP7_75t_SL g2253 ( 
.A(n_2140),
.B(n_2045),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_SL g2254 ( 
.A(n_2176),
.B(n_2048),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_SL g2255 ( 
.A(n_2176),
.B(n_2033),
.Y(n_2255)
);

AND2x4_ASAP7_75t_L g2256 ( 
.A(n_2106),
.B(n_1951),
.Y(n_2256)
);

NAND2xp33_ASAP7_75t_SL g2257 ( 
.A(n_2165),
.B(n_2005),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_SL g2258 ( 
.A(n_2208),
.B(n_2083),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_SL g2259 ( 
.A(n_2209),
.B(n_1957),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_2210),
.B(n_1918),
.Y(n_2260)
);

NAND2xp33_ASAP7_75t_SL g2261 ( 
.A(n_2165),
.B(n_866),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_2213),
.B(n_1949),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2105),
.B(n_1950),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_2221),
.B(n_866),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2130),
.B(n_2023),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_2128),
.B(n_867),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_2151),
.B(n_867),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2158),
.B(n_1921),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_2132),
.B(n_868),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2143),
.B(n_1168),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2216),
.B(n_868),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_2149),
.B(n_872),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_2187),
.B(n_2111),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_2168),
.B(n_872),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_2192),
.B(n_873),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_SL g2276 ( 
.A(n_2192),
.B(n_873),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_SL g2277 ( 
.A(n_2146),
.B(n_874),
.Y(n_2277)
);

AND2x4_ASAP7_75t_L g2278 ( 
.A(n_2092),
.B(n_884),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_2119),
.B(n_874),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_SL g2280 ( 
.A(n_2119),
.B(n_2177),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_2119),
.B(n_876),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_2206),
.B(n_876),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_SL g2283 ( 
.A(n_2102),
.B(n_877),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_2185),
.B(n_877),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_SL g2285 ( 
.A(n_2186),
.B(n_878),
.Y(n_2285)
);

AND2x4_ASAP7_75t_L g2286 ( 
.A(n_2118),
.B(n_897),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_2165),
.B(n_878),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_SL g2288 ( 
.A(n_2197),
.B(n_2215),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_2218),
.B(n_879),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_2133),
.B(n_879),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_2152),
.B(n_886),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2178),
.B(n_1963),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_SL g2293 ( 
.A(n_2238),
.B(n_886),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2238),
.B(n_887),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_2238),
.B(n_887),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_2170),
.B(n_888),
.Y(n_2296)
);

NAND2xp33_ASAP7_75t_SL g2297 ( 
.A(n_2108),
.B(n_888),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_SL g2298 ( 
.A(n_2124),
.B(n_1100),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_2230),
.B(n_1172),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_2100),
.B(n_999),
.Y(n_2300)
);

AND2x4_ASAP7_75t_L g2301 ( 
.A(n_2127),
.B(n_898),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_2122),
.B(n_1100),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2115),
.B(n_1252),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_2157),
.B(n_1252),
.Y(n_2304)
);

NAND2xp33_ASAP7_75t_SL g2305 ( 
.A(n_2183),
.B(n_1254),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2190),
.B(n_1996),
.Y(n_2306)
);

NAND2xp33_ASAP7_75t_SL g2307 ( 
.A(n_2183),
.B(n_1254),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_2173),
.B(n_1256),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2193),
.B(n_901),
.Y(n_2309)
);

AND2x4_ASAP7_75t_L g2310 ( 
.A(n_2138),
.B(n_904),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_2167),
.B(n_1256),
.Y(n_2311)
);

NAND2xp33_ASAP7_75t_SL g2312 ( 
.A(n_2183),
.B(n_1257),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_2181),
.B(n_1257),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_2086),
.B(n_1259),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2087),
.B(n_2090),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_SL g2316 ( 
.A(n_2103),
.B(n_1259),
.Y(n_2316)
);

NAND2xp33_ASAP7_75t_SL g2317 ( 
.A(n_2214),
.B(n_1264),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2198),
.B(n_2196),
.Y(n_2318)
);

NAND2xp33_ASAP7_75t_SL g2319 ( 
.A(n_2113),
.B(n_2137),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2237),
.B(n_1264),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_2222),
.B(n_1267),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_2121),
.B(n_1267),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_2125),
.B(n_1269),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_2116),
.B(n_2145),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_SL g2325 ( 
.A(n_2154),
.B(n_1269),
.Y(n_2325)
);

AND2x4_ASAP7_75t_L g2326 ( 
.A(n_2114),
.B(n_906),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_2211),
.B(n_1270),
.Y(n_2327)
);

NAND2xp33_ASAP7_75t_SL g2328 ( 
.A(n_2211),
.B(n_1270),
.Y(n_2328)
);

AND2x4_ASAP7_75t_L g2329 ( 
.A(n_2161),
.B(n_2129),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_SL g2330 ( 
.A(n_2211),
.B(n_2180),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_SL g2331 ( 
.A(n_2141),
.B(n_1271),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_SL g2332 ( 
.A(n_2096),
.B(n_1271),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_SL g2333 ( 
.A(n_2226),
.B(n_1273),
.Y(n_2333)
);

NAND2xp33_ASAP7_75t_SL g2334 ( 
.A(n_2099),
.B(n_2202),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_2153),
.B(n_1273),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_2134),
.B(n_1184),
.Y(n_2336)
);

NAND2xp33_ASAP7_75t_SL g2337 ( 
.A(n_2201),
.B(n_1058),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2220),
.B(n_907),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_2135),
.B(n_1184),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_2229),
.B(n_1238),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2182),
.B(n_908),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_2162),
.B(n_1238),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2131),
.B(n_1251),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_SL g2344 ( 
.A(n_2179),
.B(n_1251),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2088),
.B(n_1345),
.Y(n_2345)
);

NAND2xp33_ASAP7_75t_SL g2346 ( 
.A(n_2104),
.B(n_1064),
.Y(n_2346)
);

NAND2xp33_ASAP7_75t_SL g2347 ( 
.A(n_2156),
.B(n_1127),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_2095),
.B(n_1345),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_2139),
.B(n_1001),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_2101),
.B(n_1003),
.Y(n_2350)
);

NAND2xp33_ASAP7_75t_SL g2351 ( 
.A(n_2164),
.B(n_1127),
.Y(n_2351)
);

NAND2xp33_ASAP7_75t_SL g2352 ( 
.A(n_2219),
.B(n_1155),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_SL g2353 ( 
.A(n_2091),
.B(n_1007),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_SL g2354 ( 
.A(n_2231),
.B(n_1009),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_SL g2355 ( 
.A(n_2171),
.B(n_1010),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2236),
.B(n_915),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_2172),
.B(n_2175),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2184),
.B(n_1012),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2131),
.B(n_1013),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_2205),
.B(n_1021),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_SL g2361 ( 
.A(n_2144),
.B(n_1023),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_2147),
.B(n_1025),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_SL g2363 ( 
.A(n_2150),
.B(n_1026),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_2166),
.B(n_1029),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_SL g2365 ( 
.A(n_2166),
.B(n_1031),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_2232),
.B(n_1033),
.Y(n_2366)
);

NAND2xp33_ASAP7_75t_SL g2367 ( 
.A(n_2235),
.B(n_1155),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_2233),
.B(n_1036),
.Y(n_2368)
);

AND2x4_ASAP7_75t_L g2369 ( 
.A(n_2194),
.B(n_919),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_2212),
.B(n_1038),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_SL g2371 ( 
.A(n_2169),
.B(n_1039),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2199),
.B(n_1043),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2089),
.B(n_1045),
.Y(n_2373)
);

NAND2xp33_ASAP7_75t_SL g2374 ( 
.A(n_2195),
.B(n_2207),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2148),
.B(n_1046),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2093),
.B(n_920),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_SL g2377 ( 
.A(n_2142),
.B(n_1048),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_SL g2378 ( 
.A(n_2142),
.B(n_1051),
.Y(n_2378)
);

NAND2xp33_ASAP7_75t_SL g2379 ( 
.A(n_2223),
.B(n_1182),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_2203),
.B(n_2228),
.Y(n_2380)
);

AND2x4_ASAP7_75t_L g2381 ( 
.A(n_2224),
.B(n_931),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_2225),
.B(n_943),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2120),
.B(n_1056),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_2200),
.B(n_1057),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_SL g2385 ( 
.A(n_2239),
.B(n_1059),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2093),
.B(n_950),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_2117),
.B(n_1061),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_2110),
.B(n_1063),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2093),
.B(n_952),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_SL g2390 ( 
.A(n_2234),
.B(n_1066),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_SL g2391 ( 
.A(n_2159),
.B(n_1067),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_SL g2392 ( 
.A(n_2163),
.B(n_1069),
.Y(n_2392)
);

NAND2xp33_ASAP7_75t_SL g2393 ( 
.A(n_2204),
.B(n_1182),
.Y(n_2393)
);

OAI22xp5_ASAP7_75t_SL g2394 ( 
.A1(n_2300),
.A2(n_2160),
.B1(n_2191),
.B2(n_2249),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2251),
.B(n_2174),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2270),
.B(n_2109),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_L g2397 ( 
.A(n_2288),
.B(n_2109),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2318),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2242),
.B(n_2109),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2273),
.B(n_2123),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2359),
.B(n_2299),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2338),
.B(n_1070),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2369),
.B(n_956),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2369),
.B(n_2343),
.Y(n_2404)
);

INVx3_ASAP7_75t_L g2405 ( 
.A(n_2256),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2315),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_2247),
.Y(n_2407)
);

HB1xp67_ASAP7_75t_L g2408 ( 
.A(n_2329),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2245),
.B(n_1075),
.Y(n_2409)
);

CKINVDCx5p33_ASAP7_75t_R g2410 ( 
.A(n_2329),
.Y(n_2410)
);

OR2x2_ASAP7_75t_L g2411 ( 
.A(n_2324),
.B(n_957),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2341),
.B(n_1076),
.Y(n_2412)
);

OAI21x1_ASAP7_75t_L g2413 ( 
.A1(n_2262),
.A2(n_2227),
.B(n_1253),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2381),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_2317),
.Y(n_2415)
);

INVx4_ASAP7_75t_L g2416 ( 
.A(n_2256),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2309),
.B(n_1077),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_2244),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_2250),
.B(n_1330),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_SL g2420 ( 
.A(n_2243),
.B(n_1331),
.Y(n_2420)
);

CKINVDCx8_ASAP7_75t_R g2421 ( 
.A(n_2326),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2373),
.B(n_964),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_SL g2423 ( 
.A(n_2258),
.B(n_2292),
.Y(n_2423)
);

AND2x4_ASAP7_75t_L g2424 ( 
.A(n_2280),
.B(n_792),
.Y(n_2424)
);

AND2x4_ASAP7_75t_L g2425 ( 
.A(n_2327),
.B(n_795),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2381),
.Y(n_2426)
);

INVx8_ASAP7_75t_L g2427 ( 
.A(n_2278),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2310),
.B(n_966),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2382),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_SL g2430 ( 
.A(n_2265),
.B(n_1338),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2356),
.B(n_1080),
.Y(n_2431)
);

OAI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_2380),
.A2(n_1082),
.B1(n_1083),
.B2(n_1081),
.Y(n_2432)
);

OAI22xp5_ASAP7_75t_L g2433 ( 
.A1(n_2272),
.A2(n_1088),
.B1(n_1090),
.B2(n_1086),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2382),
.Y(n_2434)
);

CKINVDCx5p33_ASAP7_75t_R g2435 ( 
.A(n_2297),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2357),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2274),
.B(n_1091),
.Y(n_2437)
);

BUFx6f_ASAP7_75t_L g2438 ( 
.A(n_2278),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2286),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2266),
.B(n_1092),
.Y(n_2440)
);

HB1xp67_ASAP7_75t_L g2441 ( 
.A(n_2310),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2286),
.Y(n_2442)
);

AND2x4_ASAP7_75t_L g2443 ( 
.A(n_2330),
.B(n_796),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2269),
.B(n_1093),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2301),
.Y(n_2445)
);

CKINVDCx5p33_ASAP7_75t_R g2446 ( 
.A(n_2277),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2246),
.B(n_1333),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2301),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2240),
.B(n_1094),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2283),
.B(n_1095),
.Y(n_2450)
);

HB1xp67_ASAP7_75t_L g2451 ( 
.A(n_2326),
.Y(n_2451)
);

BUFx4f_ASAP7_75t_L g2452 ( 
.A(n_2248),
.Y(n_2452)
);

CKINVDCx5p33_ASAP7_75t_R g2453 ( 
.A(n_2390),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2321),
.B(n_969),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2319),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_2241),
.B(n_1337),
.Y(n_2456)
);

INVxp67_ASAP7_75t_SL g2457 ( 
.A(n_2306),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2384),
.B(n_1096),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2333),
.B(n_1098),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2376),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2386),
.Y(n_2461)
);

AND2x2_ASAP7_75t_L g2462 ( 
.A(n_2264),
.B(n_972),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2389),
.Y(n_2463)
);

AOI22xp5_ASAP7_75t_L g2464 ( 
.A1(n_2260),
.A2(n_2344),
.B1(n_2267),
.B2(n_2253),
.Y(n_2464)
);

INVx1_ASAP7_75t_SL g2465 ( 
.A(n_2328),
.Y(n_2465)
);

AOI22xp33_ASAP7_75t_L g2466 ( 
.A1(n_2361),
.A2(n_979),
.B1(n_982),
.B2(n_973),
.Y(n_2466)
);

HB1xp67_ASAP7_75t_L g2467 ( 
.A(n_2293),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2284),
.B(n_986),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2285),
.B(n_989),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2296),
.B(n_995),
.Y(n_2470)
);

NOR2xp67_ASAP7_75t_L g2471 ( 
.A(n_2268),
.B(n_800),
.Y(n_2471)
);

AOI22xp5_ASAP7_75t_L g2472 ( 
.A1(n_2308),
.A2(n_1103),
.B1(n_1104),
.B2(n_1099),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2263),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_SL g2474 ( 
.A(n_2271),
.B(n_1334),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2367),
.Y(n_2475)
);

AND3x1_ASAP7_75t_SL g2476 ( 
.A(n_2340),
.B(n_1004),
.C(n_998),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2354),
.B(n_1005),
.Y(n_2477)
);

BUFx6f_ASAP7_75t_L g2478 ( 
.A(n_2252),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2259),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_2377),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2334),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2303),
.B(n_1108),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2355),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2298),
.B(n_1008),
.Y(n_2484)
);

AOI22xp33_ASAP7_75t_L g2485 ( 
.A1(n_2368),
.A2(n_1015),
.B1(n_1022),
.B2(n_1011),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2311),
.B(n_1111),
.Y(n_2486)
);

OAI22xp5_ASAP7_75t_L g2487 ( 
.A1(n_2290),
.A2(n_1114),
.B1(n_1118),
.B2(n_1112),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2313),
.B(n_1120),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2314),
.B(n_1027),
.Y(n_2489)
);

NOR2xp33_ASAP7_75t_L g2490 ( 
.A(n_2289),
.B(n_2342),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2331),
.B(n_1121),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2350),
.B(n_1122),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2358),
.Y(n_2493)
);

INVx3_ASAP7_75t_L g2494 ( 
.A(n_2257),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2316),
.B(n_1028),
.Y(n_2495)
);

CKINVDCx16_ASAP7_75t_R g2496 ( 
.A(n_2261),
.Y(n_2496)
);

CKINVDCx20_ASAP7_75t_R g2497 ( 
.A(n_2305),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2387),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2349),
.B(n_1123),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_SL g2500 ( 
.A(n_2360),
.B(n_1125),
.Y(n_2500)
);

AOI22xp33_ASAP7_75t_L g2501 ( 
.A1(n_2370),
.A2(n_1040),
.B1(n_1041),
.B2(n_1030),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2332),
.Y(n_2502)
);

BUFx6f_ASAP7_75t_L g2503 ( 
.A(n_2254),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2294),
.B(n_1132),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_2378),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2352),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2362),
.B(n_1134),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2325),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2295),
.B(n_1135),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2304),
.Y(n_2510)
);

CKINVDCx11_ASAP7_75t_R g2511 ( 
.A(n_2302),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2335),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2363),
.B(n_1136),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2364),
.B(n_2365),
.Y(n_2514)
);

BUFx12f_ASAP7_75t_L g2515 ( 
.A(n_2307),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2392),
.B(n_1044),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2291),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2322),
.B(n_1139),
.Y(n_2518)
);

HB1xp67_ASAP7_75t_L g2519 ( 
.A(n_2323),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2255),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2336),
.B(n_1140),
.Y(n_2521)
);

CKINVDCx16_ASAP7_75t_R g2522 ( 
.A(n_2312),
.Y(n_2522)
);

CKINVDCx20_ASAP7_75t_R g2523 ( 
.A(n_2383),
.Y(n_2523)
);

AOI22xp5_ASAP7_75t_L g2524 ( 
.A1(n_2339),
.A2(n_1142),
.B1(n_1144),
.B2(n_1141),
.Y(n_2524)
);

OAI22xp5_ASAP7_75t_SL g2525 ( 
.A1(n_2320),
.A2(n_1055),
.B1(n_1060),
.B2(n_1049),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2346),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2375),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_SL g2528 ( 
.A(n_2345),
.B(n_1145),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_2275),
.Y(n_2529)
);

AND2x2_ASAP7_75t_SL g2530 ( 
.A(n_2391),
.B(n_1239),
.Y(n_2530)
);

OAI22xp5_ASAP7_75t_L g2531 ( 
.A1(n_2348),
.A2(n_1148),
.B1(n_1149),
.B2(n_1146),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2353),
.Y(n_2532)
);

BUFx6f_ASAP7_75t_L g2533 ( 
.A(n_2276),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2379),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_L g2535 ( 
.A(n_2366),
.B(n_1150),
.Y(n_2535)
);

OR2x2_ASAP7_75t_L g2536 ( 
.A(n_2287),
.B(n_1065),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2282),
.B(n_1152),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_L g2538 ( 
.A(n_2478),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2473),
.Y(n_2539)
);

NAND2x1p5_ASAP7_75t_L g2540 ( 
.A(n_2494),
.B(n_2385),
.Y(n_2540)
);

INVx1_ASAP7_75t_SL g2541 ( 
.A(n_2405),
.Y(n_2541)
);

OR2x2_ASAP7_75t_L g2542 ( 
.A(n_2520),
.B(n_2279),
.Y(n_2542)
);

BUFx4f_ASAP7_75t_L g2543 ( 
.A(n_2515),
.Y(n_2543)
);

INVx3_ASAP7_75t_L g2544 ( 
.A(n_2416),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2406),
.Y(n_2545)
);

AOI21xp5_ASAP7_75t_L g2546 ( 
.A1(n_2423),
.A2(n_2393),
.B(n_2374),
.Y(n_2546)
);

INVx1_ASAP7_75t_SL g2547 ( 
.A(n_2405),
.Y(n_2547)
);

INVx4_ASAP7_75t_L g2548 ( 
.A(n_2410),
.Y(n_2548)
);

NAND2x1p5_ASAP7_75t_L g2549 ( 
.A(n_2494),
.B(n_2455),
.Y(n_2549)
);

AO21x2_ASAP7_75t_L g2550 ( 
.A1(n_2481),
.A2(n_2388),
.B(n_2371),
.Y(n_2550)
);

BUFx6f_ASAP7_75t_L g2551 ( 
.A(n_2478),
.Y(n_2551)
);

OA21x2_ASAP7_75t_L g2552 ( 
.A1(n_2413),
.A2(n_2372),
.B(n_1072),
.Y(n_2552)
);

BUFx24_ASAP7_75t_L g2553 ( 
.A(n_2443),
.Y(n_2553)
);

CKINVDCx11_ASAP7_75t_R g2554 ( 
.A(n_2421),
.Y(n_2554)
);

CKINVDCx11_ASAP7_75t_R g2555 ( 
.A(n_2497),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2479),
.Y(n_2556)
);

AO21x2_ASAP7_75t_L g2557 ( 
.A1(n_2464),
.A2(n_2281),
.B(n_1074),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2436),
.Y(n_2558)
);

AO21x2_ASAP7_75t_L g2559 ( 
.A1(n_2464),
.A2(n_1084),
.B(n_1071),
.Y(n_2559)
);

BUFx3_ASAP7_75t_L g2560 ( 
.A(n_2427),
.Y(n_2560)
);

BUFx2_ASAP7_75t_L g2561 ( 
.A(n_2416),
.Y(n_2561)
);

AO21x2_ASAP7_75t_L g2562 ( 
.A1(n_2400),
.A2(n_1087),
.B(n_1085),
.Y(n_2562)
);

NOR2xp67_ASAP7_75t_L g2563 ( 
.A(n_2460),
.B(n_802),
.Y(n_2563)
);

OAI21x1_ASAP7_75t_L g2564 ( 
.A1(n_2526),
.A2(n_1253),
.B(n_1239),
.Y(n_2564)
);

BUFx3_ASAP7_75t_L g2565 ( 
.A(n_2427),
.Y(n_2565)
);

BUFx6f_ASAP7_75t_L g2566 ( 
.A(n_2478),
.Y(n_2566)
);

AO21x2_ASAP7_75t_L g2567 ( 
.A1(n_2399),
.A2(n_1106),
.B(n_1097),
.Y(n_2567)
);

INVx2_ASAP7_75t_SL g2568 ( 
.A(n_2427),
.Y(n_2568)
);

OAI21x1_ASAP7_75t_L g2569 ( 
.A1(n_2475),
.A2(n_1305),
.B(n_1113),
.Y(n_2569)
);

AOI22x1_ASAP7_75t_L g2570 ( 
.A1(n_2418),
.A2(n_2506),
.B1(n_2465),
.B2(n_2443),
.Y(n_2570)
);

OAI21x1_ASAP7_75t_L g2571 ( 
.A1(n_2527),
.A2(n_1305),
.B(n_1116),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2398),
.Y(n_2572)
);

INVx3_ASAP7_75t_L g2573 ( 
.A(n_2452),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2457),
.Y(n_2574)
);

INVx5_ASAP7_75t_L g2575 ( 
.A(n_2503),
.Y(n_2575)
);

OAI21x1_ASAP7_75t_L g2576 ( 
.A1(n_2534),
.A2(n_1119),
.B(n_1110),
.Y(n_2576)
);

AO21x2_ASAP7_75t_L g2577 ( 
.A1(n_2456),
.A2(n_1128),
.B(n_1126),
.Y(n_2577)
);

OAI21x1_ASAP7_75t_L g2578 ( 
.A1(n_2498),
.A2(n_2532),
.B(n_2471),
.Y(n_2578)
);

OAI21x1_ASAP7_75t_L g2579 ( 
.A1(n_2471),
.A2(n_1133),
.B(n_1130),
.Y(n_2579)
);

BUFx6f_ASAP7_75t_L g2580 ( 
.A(n_2503),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2461),
.Y(n_2581)
);

NAND2x1p5_ASAP7_75t_L g2582 ( 
.A(n_2452),
.B(n_1137),
.Y(n_2582)
);

BUFx2_ASAP7_75t_SL g2583 ( 
.A(n_2404),
.Y(n_2583)
);

AO21x2_ASAP7_75t_L g2584 ( 
.A1(n_2397),
.A2(n_1151),
.B(n_1143),
.Y(n_2584)
);

AO21x2_ASAP7_75t_L g2585 ( 
.A1(n_2430),
.A2(n_1161),
.B(n_1160),
.Y(n_2585)
);

OAI21x1_ASAP7_75t_L g2586 ( 
.A1(n_2463),
.A2(n_1170),
.B(n_1164),
.Y(n_2586)
);

INVx1_ASAP7_75t_SL g2587 ( 
.A(n_2503),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2434),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2439),
.Y(n_2589)
);

INVx3_ASAP7_75t_L g2590 ( 
.A(n_2414),
.Y(n_2590)
);

AOI22x1_ASAP7_75t_L g2591 ( 
.A1(n_2465),
.A2(n_1154),
.B1(n_1156),
.B2(n_1153),
.Y(n_2591)
);

NAND2x1p5_ASAP7_75t_L g2592 ( 
.A(n_2424),
.B(n_1174),
.Y(n_2592)
);

OAI21x1_ASAP7_75t_L g2593 ( 
.A1(n_2426),
.A2(n_1192),
.B(n_1178),
.Y(n_2593)
);

OAI21x1_ASAP7_75t_L g2594 ( 
.A1(n_2429),
.A2(n_1227),
.B(n_1194),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2442),
.Y(n_2595)
);

INVx3_ASAP7_75t_L g2596 ( 
.A(n_2424),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2445),
.Y(n_2597)
);

CKINVDCx11_ASAP7_75t_R g2598 ( 
.A(n_2511),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2448),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2411),
.Y(n_2600)
);

OAI21x1_ASAP7_75t_L g2601 ( 
.A1(n_2420),
.A2(n_1240),
.B(n_1230),
.Y(n_2601)
);

INVx3_ASAP7_75t_L g2602 ( 
.A(n_2483),
.Y(n_2602)
);

OAI21x1_ASAP7_75t_L g2603 ( 
.A1(n_2395),
.A2(n_1245),
.B(n_1243),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2493),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2502),
.Y(n_2605)
);

INVx3_ASAP7_75t_L g2606 ( 
.A(n_2438),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2508),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2510),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_2415),
.Y(n_2609)
);

NAND2x1p5_ASAP7_75t_L g2610 ( 
.A(n_2438),
.B(n_1263),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2512),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2403),
.Y(n_2612)
);

AO21x2_ASAP7_75t_L g2613 ( 
.A1(n_2419),
.A2(n_1275),
.B(n_1268),
.Y(n_2613)
);

INVx3_ASAP7_75t_L g2614 ( 
.A(n_2438),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_L g2615 ( 
.A(n_2423),
.B(n_2394),
.Y(n_2615)
);

OAI21x1_ASAP7_75t_L g2616 ( 
.A1(n_2501),
.A2(n_1282),
.B(n_1280),
.Y(n_2616)
);

OAI21x1_ASAP7_75t_SL g2617 ( 
.A1(n_2409),
.A2(n_1292),
.B(n_1289),
.Y(n_2617)
);

BUFx3_ASAP7_75t_L g2618 ( 
.A(n_2408),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2517),
.Y(n_2619)
);

BUFx12f_ASAP7_75t_L g2620 ( 
.A(n_2529),
.Y(n_2620)
);

BUFx12f_ASAP7_75t_L g2621 ( 
.A(n_2435),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2519),
.Y(n_2622)
);

OAI21xp5_ASAP7_75t_L g2623 ( 
.A1(n_2530),
.A2(n_2351),
.B(n_2347),
.Y(n_2623)
);

AOI22xp33_ASAP7_75t_SL g2624 ( 
.A1(n_2394),
.A2(n_1158),
.B1(n_1159),
.B2(n_1157),
.Y(n_2624)
);

BUFx3_ASAP7_75t_L g2625 ( 
.A(n_2451),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2490),
.B(n_1298),
.Y(n_2626)
);

AOI21x1_ASAP7_75t_L g2627 ( 
.A1(n_2447),
.A2(n_1306),
.B(n_1303),
.Y(n_2627)
);

OAI21x1_ASAP7_75t_L g2628 ( 
.A1(n_2396),
.A2(n_1325),
.B(n_1313),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2441),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2425),
.B(n_1327),
.Y(n_2630)
);

INVx2_ASAP7_75t_SL g2631 ( 
.A(n_2533),
.Y(n_2631)
);

BUFx3_ASAP7_75t_L g2632 ( 
.A(n_2401),
.Y(n_2632)
);

OAI21x1_ASAP7_75t_L g2633 ( 
.A1(n_2500),
.A2(n_1340),
.B(n_1329),
.Y(n_2633)
);

NAND2x1p5_ASAP7_75t_L g2634 ( 
.A(n_2425),
.B(n_1341),
.Y(n_2634)
);

INVx8_ASAP7_75t_L g2635 ( 
.A(n_2533),
.Y(n_2635)
);

HB1xp67_ASAP7_75t_L g2636 ( 
.A(n_2467),
.Y(n_2636)
);

AO21x2_ASAP7_75t_L g2637 ( 
.A1(n_2449),
.A2(n_1342),
.B(n_2337),
.Y(n_2637)
);

OAI21x1_ASAP7_75t_SL g2638 ( 
.A1(n_2514),
.A2(n_2),
.B(n_4),
.Y(n_2638)
);

AOI22xp33_ASAP7_75t_L g2639 ( 
.A1(n_2525),
.A2(n_1165),
.B1(n_1166),
.B2(n_1162),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2516),
.Y(n_2640)
);

OAI21x1_ASAP7_75t_L g2641 ( 
.A1(n_2458),
.A2(n_806),
.B(n_804),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2428),
.Y(n_2642)
);

BUFx2_ASAP7_75t_L g2643 ( 
.A(n_2407),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2533),
.B(n_807),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2422),
.B(n_810),
.Y(n_2645)
);

INVx1_ASAP7_75t_SL g2646 ( 
.A(n_2477),
.Y(n_2646)
);

OAI21x1_ASAP7_75t_L g2647 ( 
.A1(n_2528),
.A2(n_2),
.B(n_4),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2556),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2574),
.Y(n_2649)
);

INVx8_ASAP7_75t_L g2650 ( 
.A(n_2635),
.Y(n_2650)
);

AOI22xp33_ASAP7_75t_SL g2651 ( 
.A1(n_2615),
.A2(n_2525),
.B1(n_2535),
.B2(n_2507),
.Y(n_2651)
);

INVx6_ASAP7_75t_L g2652 ( 
.A(n_2548),
.Y(n_2652)
);

BUFx8_ASAP7_75t_SL g2653 ( 
.A(n_2543),
.Y(n_2653)
);

INVx6_ASAP7_75t_L g2654 ( 
.A(n_2548),
.Y(n_2654)
);

AOI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2615),
.A2(n_2522),
.B1(n_2496),
.B2(n_2453),
.Y(n_2655)
);

AOI22xp33_ASAP7_75t_L g2656 ( 
.A1(n_2624),
.A2(n_2432),
.B1(n_2454),
.B2(n_2462),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2545),
.Y(n_2657)
);

AOI22xp33_ASAP7_75t_L g2658 ( 
.A1(n_2624),
.A2(n_2469),
.B1(n_2470),
.B2(n_2468),
.Y(n_2658)
);

BUFx2_ASAP7_75t_L g2659 ( 
.A(n_2625),
.Y(n_2659)
);

AOI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_2570),
.A2(n_2474),
.B1(n_2523),
.B2(n_2495),
.Y(n_2660)
);

CKINVDCx11_ASAP7_75t_R g2661 ( 
.A(n_2598),
.Y(n_2661)
);

NAND2x1p5_ASAP7_75t_L g2662 ( 
.A(n_2575),
.B(n_2544),
.Y(n_2662)
);

BUFx2_ASAP7_75t_SL g2663 ( 
.A(n_2573),
.Y(n_2663)
);

OAI22xp5_ASAP7_75t_L g2664 ( 
.A1(n_2634),
.A2(n_2446),
.B1(n_2485),
.B2(n_2466),
.Y(n_2664)
);

INVx3_ASAP7_75t_L g2665 ( 
.A(n_2538),
.Y(n_2665)
);

CKINVDCx8_ASAP7_75t_R g2666 ( 
.A(n_2609),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2556),
.Y(n_2667)
);

OAI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2634),
.A2(n_2480),
.B1(n_2505),
.B2(n_2524),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2572),
.Y(n_2669)
);

AOI22xp33_ASAP7_75t_L g2670 ( 
.A1(n_2559),
.A2(n_2484),
.B1(n_2489),
.B2(n_2459),
.Y(n_2670)
);

CKINVDCx11_ASAP7_75t_R g2671 ( 
.A(n_2598),
.Y(n_2671)
);

OAI22xp5_ASAP7_75t_L g2672 ( 
.A1(n_2639),
.A2(n_2592),
.B1(n_2646),
.B2(n_2573),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2539),
.Y(n_2673)
);

BUFx4f_ASAP7_75t_L g2674 ( 
.A(n_2621),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2572),
.Y(n_2675)
);

BUFx6f_ASAP7_75t_L g2676 ( 
.A(n_2538),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2558),
.Y(n_2677)
);

OR2x2_ASAP7_75t_L g2678 ( 
.A(n_2646),
.B(n_2636),
.Y(n_2678)
);

AOI22xp33_ASAP7_75t_L g2679 ( 
.A1(n_2559),
.A2(n_2499),
.B1(n_2513),
.B2(n_2492),
.Y(n_2679)
);

AOI22xp33_ASAP7_75t_SL g2680 ( 
.A1(n_2557),
.A2(n_2433),
.B1(n_2437),
.B2(n_2402),
.Y(n_2680)
);

AOI22xp33_ASAP7_75t_L g2681 ( 
.A1(n_2557),
.A2(n_2521),
.B1(n_2536),
.B2(n_2504),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2581),
.Y(n_2682)
);

OAI22xp5_ASAP7_75t_L g2683 ( 
.A1(n_2639),
.A2(n_2524),
.B1(n_2472),
.B2(n_2417),
.Y(n_2683)
);

OAI22xp5_ASAP7_75t_L g2684 ( 
.A1(n_2592),
.A2(n_2472),
.B1(n_2431),
.B2(n_2509),
.Y(n_2684)
);

BUFx8_ASAP7_75t_SL g2685 ( 
.A(n_2543),
.Y(n_2685)
);

CKINVDCx20_ASAP7_75t_R g2686 ( 
.A(n_2555),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2636),
.B(n_2412),
.Y(n_2687)
);

CKINVDCx20_ASAP7_75t_R g2688 ( 
.A(n_2555),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2588),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2605),
.Y(n_2690)
);

BUFx2_ASAP7_75t_R g2691 ( 
.A(n_2609),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2622),
.B(n_2444),
.Y(n_2692)
);

BUFx3_ASAP7_75t_L g2693 ( 
.A(n_2635),
.Y(n_2693)
);

AOI22xp33_ASAP7_75t_L g2694 ( 
.A1(n_2596),
.A2(n_2450),
.B1(n_2440),
.B2(n_2482),
.Y(n_2694)
);

NAND2x1p5_ASAP7_75t_L g2695 ( 
.A(n_2575),
.B(n_2486),
.Y(n_2695)
);

AOI22xp5_ASAP7_75t_SL g2696 ( 
.A1(n_2583),
.A2(n_2487),
.B1(n_1169),
.B2(n_1171),
.Y(n_2696)
);

INVxp67_ASAP7_75t_L g2697 ( 
.A(n_2632),
.Y(n_2697)
);

INVx1_ASAP7_75t_SL g2698 ( 
.A(n_2643),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2589),
.Y(n_2699)
);

CKINVDCx5p33_ASAP7_75t_R g2700 ( 
.A(n_2554),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2595),
.Y(n_2701)
);

BUFx2_ASAP7_75t_L g2702 ( 
.A(n_2625),
.Y(n_2702)
);

INVx6_ASAP7_75t_L g2703 ( 
.A(n_2635),
.Y(n_2703)
);

CKINVDCx11_ASAP7_75t_R g2704 ( 
.A(n_2554),
.Y(n_2704)
);

INVx3_ASAP7_75t_L g2705 ( 
.A(n_2538),
.Y(n_2705)
);

AND2x2_ASAP7_75t_L g2706 ( 
.A(n_2632),
.B(n_2537),
.Y(n_2706)
);

AOI22xp33_ASAP7_75t_L g2707 ( 
.A1(n_2596),
.A2(n_2491),
.B1(n_2488),
.B2(n_2518),
.Y(n_2707)
);

INVx4_ASAP7_75t_L g2708 ( 
.A(n_2575),
.Y(n_2708)
);

INVx3_ASAP7_75t_L g2709 ( 
.A(n_2551),
.Y(n_2709)
);

INVx1_ASAP7_75t_SL g2710 ( 
.A(n_2587),
.Y(n_2710)
);

AOI22xp33_ASAP7_75t_L g2711 ( 
.A1(n_2637),
.A2(n_2531),
.B1(n_1173),
.B2(n_1175),
.Y(n_2711)
);

OAI22xp33_ASAP7_75t_L g2712 ( 
.A1(n_2626),
.A2(n_1326),
.B1(n_1198),
.B2(n_1208),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2605),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2618),
.B(n_6),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2608),
.Y(n_2715)
);

AOI22xp33_ASAP7_75t_L g2716 ( 
.A1(n_2637),
.A2(n_1176),
.B1(n_1177),
.B2(n_1167),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2608),
.Y(n_2717)
);

AOI22xp33_ASAP7_75t_L g2718 ( 
.A1(n_2642),
.A2(n_1181),
.B1(n_1183),
.B2(n_1179),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2611),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2611),
.Y(n_2720)
);

AOI22xp5_ASAP7_75t_L g2721 ( 
.A1(n_2577),
.A2(n_2476),
.B1(n_1187),
.B2(n_1189),
.Y(n_2721)
);

AOI22xp33_ASAP7_75t_L g2722 ( 
.A1(n_2642),
.A2(n_1190),
.B1(n_1193),
.B2(n_1186),
.Y(n_2722)
);

INVx4_ASAP7_75t_L g2723 ( 
.A(n_2575),
.Y(n_2723)
);

INVx6_ASAP7_75t_L g2724 ( 
.A(n_2551),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2597),
.Y(n_2725)
);

AOI22xp33_ASAP7_75t_L g2726 ( 
.A1(n_2640),
.A2(n_1196),
.B1(n_1197),
.B2(n_1195),
.Y(n_2726)
);

AOI21xp5_ASAP7_75t_L g2727 ( 
.A1(n_2683),
.A2(n_2546),
.B(n_2562),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2678),
.B(n_2619),
.Y(n_2728)
);

OA21x2_ASAP7_75t_L g2729 ( 
.A1(n_2648),
.A2(n_2578),
.B(n_2603),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2682),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2657),
.Y(n_2731)
);

AOI21xp5_ASAP7_75t_L g2732 ( 
.A1(n_2684),
.A2(n_2546),
.B(n_2562),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2687),
.B(n_2604),
.Y(n_2733)
);

OAI21x1_ASAP7_75t_L g2734 ( 
.A1(n_2662),
.A2(n_2564),
.B(n_2571),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2648),
.Y(n_2735)
);

AND2x4_ASAP7_75t_L g2736 ( 
.A(n_2659),
.B(n_2618),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2649),
.B(n_2607),
.Y(n_2737)
);

OAI21x1_ASAP7_75t_L g2738 ( 
.A1(n_2695),
.A2(n_2549),
.B(n_2569),
.Y(n_2738)
);

OR2x6_ASAP7_75t_L g2739 ( 
.A(n_2663),
.B(n_2549),
.Y(n_2739)
);

BUFx3_ASAP7_75t_L g2740 ( 
.A(n_2686),
.Y(n_2740)
);

AO31x2_ASAP7_75t_L g2741 ( 
.A1(n_2708),
.A2(n_2597),
.A3(n_2561),
.B(n_2629),
.Y(n_2741)
);

OA21x2_ASAP7_75t_L g2742 ( 
.A1(n_2670),
.A2(n_2586),
.B(n_2628),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2673),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2677),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2689),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2702),
.B(n_2631),
.Y(n_2746)
);

AOI21xp5_ASAP7_75t_L g2747 ( 
.A1(n_2679),
.A2(n_2651),
.B(n_2680),
.Y(n_2747)
);

AO21x2_ASAP7_75t_L g2748 ( 
.A1(n_2692),
.A2(n_2638),
.B(n_2584),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2699),
.B(n_2602),
.Y(n_2749)
);

AOI21xp5_ASAP7_75t_L g2750 ( 
.A1(n_2681),
.A2(n_2623),
.B(n_2694),
.Y(n_2750)
);

AOI22xp33_ASAP7_75t_L g2751 ( 
.A1(n_2672),
.A2(n_2656),
.B1(n_2706),
.B2(n_2668),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2701),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2667),
.B(n_2602),
.Y(n_2753)
);

INVx4_ASAP7_75t_SL g2754 ( 
.A(n_2652),
.Y(n_2754)
);

OAI21x1_ASAP7_75t_L g2755 ( 
.A1(n_2690),
.A2(n_2576),
.B(n_2579),
.Y(n_2755)
);

AO31x2_ASAP7_75t_L g2756 ( 
.A1(n_2708),
.A2(n_2599),
.A3(n_2626),
.B(n_2630),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2675),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2713),
.Y(n_2758)
);

AND2x4_ASAP7_75t_L g2759 ( 
.A(n_2669),
.B(n_2541),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2715),
.Y(n_2760)
);

AOI21xp5_ASAP7_75t_L g2761 ( 
.A1(n_2707),
.A2(n_2623),
.B(n_2553),
.Y(n_2761)
);

AO21x2_ASAP7_75t_L g2762 ( 
.A1(n_2717),
.A2(n_2584),
.B(n_2567),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2719),
.Y(n_2763)
);

O2A1O1Ixp33_ASAP7_75t_L g2764 ( 
.A1(n_2712),
.A2(n_2630),
.B(n_2617),
.C(n_2582),
.Y(n_2764)
);

NOR2xp33_ASAP7_75t_L g2765 ( 
.A(n_2655),
.B(n_2612),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2720),
.Y(n_2766)
);

AOI21xp5_ASAP7_75t_L g2767 ( 
.A1(n_2716),
.A2(n_2553),
.B(n_2550),
.Y(n_2767)
);

OAI22xp5_ASAP7_75t_L g2768 ( 
.A1(n_2660),
.A2(n_2540),
.B1(n_2582),
.B2(n_2610),
.Y(n_2768)
);

INVx3_ASAP7_75t_L g2769 ( 
.A(n_2652),
.Y(n_2769)
);

AOI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2664),
.A2(n_2550),
.B(n_2567),
.Y(n_2770)
);

AOI21xp5_ASAP7_75t_L g2771 ( 
.A1(n_2711),
.A2(n_2540),
.B(n_2577),
.Y(n_2771)
);

OAI221xp5_ASAP7_75t_L g2772 ( 
.A1(n_2658),
.A2(n_2610),
.B1(n_2600),
.B2(n_2542),
.C(n_2591),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2697),
.B(n_2541),
.Y(n_2773)
);

OAI221xp5_ASAP7_75t_L g2774 ( 
.A1(n_2721),
.A2(n_2696),
.B1(n_2718),
.B2(n_2722),
.C(n_2726),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_2698),
.B(n_2547),
.Y(n_2775)
);

AOI21xp5_ASAP7_75t_L g2776 ( 
.A1(n_2723),
.A2(n_2585),
.B(n_2613),
.Y(n_2776)
);

OAI21x1_ASAP7_75t_L g2777 ( 
.A1(n_2665),
.A2(n_2552),
.B(n_2641),
.Y(n_2777)
);

AND2x2_ASAP7_75t_L g2778 ( 
.A(n_2710),
.B(n_2547),
.Y(n_2778)
);

OR2x2_ASAP7_75t_L g2779 ( 
.A(n_2725),
.B(n_2587),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2714),
.B(n_2590),
.Y(n_2780)
);

AOI21xp5_ASAP7_75t_L g2781 ( 
.A1(n_2723),
.A2(n_2585),
.B(n_2613),
.Y(n_2781)
);

INVxp67_ASAP7_75t_SL g2782 ( 
.A(n_2665),
.Y(n_2782)
);

OR2x2_ASAP7_75t_L g2783 ( 
.A(n_2705),
.B(n_2590),
.Y(n_2783)
);

AOI21xp5_ASAP7_75t_L g2784 ( 
.A1(n_2674),
.A2(n_2563),
.B(n_2552),
.Y(n_2784)
);

INVx3_ASAP7_75t_L g2785 ( 
.A(n_2654),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2705),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2709),
.B(n_2551),
.Y(n_2787)
);

OA21x2_ASAP7_75t_L g2788 ( 
.A1(n_2700),
.A2(n_2647),
.B(n_2594),
.Y(n_2788)
);

AOI21xp5_ASAP7_75t_L g2789 ( 
.A1(n_2674),
.A2(n_2544),
.B(n_2568),
.Y(n_2789)
);

AND2x4_ASAP7_75t_L g2790 ( 
.A(n_2709),
.B(n_2560),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_L g2791 ( 
.A(n_2654),
.B(n_2620),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2676),
.B(n_2566),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2676),
.Y(n_2793)
);

AOI21xp5_ASAP7_75t_L g2794 ( 
.A1(n_2650),
.A2(n_2601),
.B(n_2593),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2676),
.B(n_2566),
.Y(n_2795)
);

A2O1A1Ixp33_ASAP7_75t_L g2796 ( 
.A1(n_2688),
.A2(n_2645),
.B(n_2644),
.C(n_2633),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2724),
.B(n_2566),
.Y(n_2797)
);

AOI221xp5_ASAP7_75t_L g2798 ( 
.A1(n_2693),
.A2(n_1335),
.B1(n_1328),
.B2(n_1203),
.C(n_1204),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2724),
.B(n_2606),
.Y(n_2799)
);

INVx4_ASAP7_75t_SL g2800 ( 
.A(n_2756),
.Y(n_2800)
);

AOI22xp33_ASAP7_75t_L g2801 ( 
.A1(n_2747),
.A2(n_2644),
.B1(n_2671),
.B2(n_2661),
.Y(n_2801)
);

INVxp67_ASAP7_75t_L g2802 ( 
.A(n_2735),
.Y(n_2802)
);

O2A1O1Ixp33_ASAP7_75t_L g2803 ( 
.A1(n_2727),
.A2(n_2770),
.B(n_2774),
.C(n_2732),
.Y(n_2803)
);

AOI22xp33_ASAP7_75t_L g2804 ( 
.A1(n_2750),
.A2(n_2704),
.B1(n_2580),
.B2(n_2614),
.Y(n_2804)
);

AOI22xp33_ASAP7_75t_L g2805 ( 
.A1(n_2761),
.A2(n_2580),
.B1(n_2614),
.B2(n_2606),
.Y(n_2805)
);

AOI22xp33_ASAP7_75t_L g2806 ( 
.A1(n_2767),
.A2(n_2580),
.B1(n_2565),
.B2(n_2560),
.Y(n_2806)
);

BUFx2_ASAP7_75t_L g2807 ( 
.A(n_2736),
.Y(n_2807)
);

AOI22xp33_ASAP7_75t_L g2808 ( 
.A1(n_2772),
.A2(n_2565),
.B1(n_2703),
.B2(n_2685),
.Y(n_2808)
);

AOI22xp33_ASAP7_75t_L g2809 ( 
.A1(n_2768),
.A2(n_2703),
.B1(n_2653),
.B2(n_2650),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2743),
.Y(n_2810)
);

OAI221xp5_ASAP7_75t_L g2811 ( 
.A1(n_2751),
.A2(n_2666),
.B1(n_1205),
.B2(n_1206),
.C(n_1202),
.Y(n_2811)
);

AOI22xp33_ASAP7_75t_SL g2812 ( 
.A1(n_2748),
.A2(n_2616),
.B1(n_2691),
.B2(n_1207),
.Y(n_2812)
);

OAI21x1_ASAP7_75t_L g2813 ( 
.A1(n_2776),
.A2(n_2627),
.B(n_6),
.Y(n_2813)
);

AOI22xp33_ASAP7_75t_L g2814 ( 
.A1(n_2771),
.A2(n_1310),
.B1(n_1311),
.B2(n_1309),
.Y(n_2814)
);

OAI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2739),
.A2(n_1210),
.B1(n_1212),
.B2(n_1200),
.Y(n_2815)
);

NAND3xp33_ASAP7_75t_L g2816 ( 
.A(n_2781),
.B(n_1214),
.C(n_1213),
.Y(n_2816)
);

AND2x2_ASAP7_75t_L g2817 ( 
.A(n_2736),
.B(n_7),
.Y(n_2817)
);

AOI22xp33_ASAP7_75t_SL g2818 ( 
.A1(n_2765),
.A2(n_1218),
.B1(n_1219),
.B2(n_1217),
.Y(n_2818)
);

NAND4xp25_ASAP7_75t_L g2819 ( 
.A(n_2764),
.B(n_9),
.C(n_7),
.D(n_8),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2745),
.Y(n_2820)
);

CKINVDCx5p33_ASAP7_75t_R g2821 ( 
.A(n_2740),
.Y(n_2821)
);

A2O1A1Ixp33_ASAP7_75t_L g2822 ( 
.A1(n_2796),
.A2(n_2784),
.B(n_2789),
.C(n_2798),
.Y(n_2822)
);

AOI21xp5_ASAP7_75t_L g2823 ( 
.A1(n_2794),
.A2(n_2742),
.B(n_2762),
.Y(n_2823)
);

HB1xp67_ASAP7_75t_L g2824 ( 
.A(n_2741),
.Y(n_2824)
);

AOI22xp33_ASAP7_75t_L g2825 ( 
.A1(n_2788),
.A2(n_1301),
.B1(n_1302),
.B2(n_1300),
.Y(n_2825)
);

OAI22xp5_ASAP7_75t_L g2826 ( 
.A1(n_2739),
.A2(n_1221),
.B1(n_1222),
.B2(n_1220),
.Y(n_2826)
);

AOI22xp33_ASAP7_75t_L g2827 ( 
.A1(n_2788),
.A2(n_1319),
.B1(n_1322),
.B2(n_1315),
.Y(n_2827)
);

AOI22xp33_ASAP7_75t_L g2828 ( 
.A1(n_2742),
.A2(n_1324),
.B1(n_1323),
.B2(n_1224),
.Y(n_2828)
);

AND2x2_ASAP7_75t_L g2829 ( 
.A(n_2775),
.B(n_10),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2752),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2731),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2746),
.B(n_12),
.Y(n_2832)
);

INVx2_ASAP7_75t_SL g2833 ( 
.A(n_2769),
.Y(n_2833)
);

OAI22xp5_ASAP7_75t_L g2834 ( 
.A1(n_2769),
.A2(n_1225),
.B1(n_1228),
.B2(n_1223),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_2773),
.B(n_2778),
.Y(n_2835)
);

OAI21x1_ASAP7_75t_L g2836 ( 
.A1(n_2777),
.A2(n_12),
.B(n_13),
.Y(n_2836)
);

AOI22xp33_ASAP7_75t_L g2837 ( 
.A1(n_2785),
.A2(n_1286),
.B1(n_1287),
.B2(n_1285),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2757),
.Y(n_2838)
);

INVx4_ASAP7_75t_L g2839 ( 
.A(n_2754),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2733),
.B(n_1233),
.Y(n_2840)
);

OAI221xp5_ASAP7_75t_L g2841 ( 
.A1(n_2780),
.A2(n_1241),
.B1(n_1246),
.B2(n_1237),
.C(n_1234),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2730),
.Y(n_2842)
);

HB1xp67_ASAP7_75t_L g2843 ( 
.A(n_2802),
.Y(n_2843)
);

INVx1_ASAP7_75t_SL g2844 ( 
.A(n_2807),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2824),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2802),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2838),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2810),
.Y(n_2848)
);

HB1xp67_ASAP7_75t_L g2849 ( 
.A(n_2831),
.Y(n_2849)
);

OR2x2_ASAP7_75t_L g2850 ( 
.A(n_2842),
.B(n_2728),
.Y(n_2850)
);

AOI221x1_ASAP7_75t_L g2851 ( 
.A1(n_2819),
.A2(n_2786),
.B1(n_2795),
.B2(n_2792),
.C(n_2793),
.Y(n_2851)
);

AND2x2_ASAP7_75t_L g2852 ( 
.A(n_2835),
.B(n_2785),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2820),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2830),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2833),
.B(n_2782),
.Y(n_2855)
);

AND2x2_ASAP7_75t_L g2856 ( 
.A(n_2800),
.B(n_2753),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2800),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2800),
.B(n_2753),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2836),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2803),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2803),
.Y(n_2861)
);

HB1xp67_ASAP7_75t_L g2862 ( 
.A(n_2829),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2814),
.B(n_2756),
.Y(n_2863)
);

AND2x4_ASAP7_75t_L g2864 ( 
.A(n_2839),
.B(n_2754),
.Y(n_2864)
);

AND2x4_ASAP7_75t_L g2865 ( 
.A(n_2839),
.B(n_2741),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2817),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2813),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2832),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2806),
.B(n_2756),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2805),
.B(n_2744),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2840),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2816),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2804),
.B(n_2758),
.Y(n_2873)
);

OR2x2_ASAP7_75t_L g2874 ( 
.A(n_2823),
.B(n_2779),
.Y(n_2874)
);

BUFx3_ASAP7_75t_L g2875 ( 
.A(n_2821),
.Y(n_2875)
);

NOR2xp33_ASAP7_75t_L g2876 ( 
.A(n_2841),
.B(n_2791),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2826),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2834),
.Y(n_2878)
);

INVx5_ASAP7_75t_L g2879 ( 
.A(n_2825),
.Y(n_2879)
);

AOI22xp33_ASAP7_75t_SL g2880 ( 
.A1(n_2879),
.A2(n_2811),
.B1(n_2823),
.B2(n_2822),
.Y(n_2880)
);

OAI21x1_ASAP7_75t_L g2881 ( 
.A1(n_2857),
.A2(n_2766),
.B(n_2760),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2860),
.B(n_2827),
.Y(n_2882)
);

OA21x2_ASAP7_75t_L g2883 ( 
.A1(n_2861),
.A2(n_2845),
.B(n_2851),
.Y(n_2883)
);

AOI222xp33_ASAP7_75t_L g2884 ( 
.A1(n_2879),
.A2(n_2861),
.B1(n_2872),
.B2(n_2871),
.C1(n_2863),
.C2(n_2877),
.Y(n_2884)
);

HB1xp67_ASAP7_75t_L g2885 ( 
.A(n_2843),
.Y(n_2885)
);

AO31x2_ASAP7_75t_L g2886 ( 
.A1(n_2851),
.A2(n_2797),
.A3(n_2787),
.B(n_2763),
.Y(n_2886)
);

AOI31xp33_ASAP7_75t_L g2887 ( 
.A1(n_2864),
.A2(n_2801),
.A3(n_2808),
.B(n_2809),
.Y(n_2887)
);

INVx4_ASAP7_75t_L g2888 ( 
.A(n_2864),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2865),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2853),
.Y(n_2890)
);

OAI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2879),
.A2(n_2818),
.B(n_2828),
.Y(n_2891)
);

CKINVDCx5p33_ASAP7_75t_R g2892 ( 
.A(n_2875),
.Y(n_2892)
);

BUFx2_ASAP7_75t_L g2893 ( 
.A(n_2864),
.Y(n_2893)
);

INVxp67_ASAP7_75t_SL g2894 ( 
.A(n_2874),
.Y(n_2894)
);

OAI21xp33_ASAP7_75t_SL g2895 ( 
.A1(n_2869),
.A2(n_2738),
.B(n_2749),
.Y(n_2895)
);

AOI21xp33_ASAP7_75t_SL g2896 ( 
.A1(n_2872),
.A2(n_2818),
.B(n_2877),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2844),
.B(n_2799),
.Y(n_2897)
);

INVxp67_ASAP7_75t_L g2898 ( 
.A(n_2873),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2853),
.Y(n_2899)
);

INVx4_ASAP7_75t_SL g2900 ( 
.A(n_2875),
.Y(n_2900)
);

OR2x2_ASAP7_75t_L g2901 ( 
.A(n_2867),
.B(n_2759),
.Y(n_2901)
);

OAI21xp33_ASAP7_75t_L g2902 ( 
.A1(n_2878),
.A2(n_2812),
.B(n_2837),
.Y(n_2902)
);

NAND4xp25_ASAP7_75t_L g2903 ( 
.A(n_2871),
.B(n_2812),
.C(n_2737),
.D(n_2783),
.Y(n_2903)
);

AOI21xp5_ASAP7_75t_L g2904 ( 
.A1(n_2879),
.A2(n_2815),
.B(n_2790),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2847),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2865),
.Y(n_2906)
);

O2A1O1Ixp5_ASAP7_75t_L g2907 ( 
.A1(n_2865),
.A2(n_2759),
.B(n_2790),
.C(n_2741),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2852),
.B(n_2729),
.Y(n_2908)
);

INVxp67_ASAP7_75t_L g2909 ( 
.A(n_2878),
.Y(n_2909)
);

OAI22xp5_ASAP7_75t_L g2910 ( 
.A1(n_2879),
.A2(n_2868),
.B1(n_2862),
.B2(n_2859),
.Y(n_2910)
);

AOI21xp5_ASAP7_75t_L g2911 ( 
.A1(n_2876),
.A2(n_2729),
.B(n_2755),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2855),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2855),
.Y(n_2913)
);

NOR2xp33_ASAP7_75t_L g2914 ( 
.A(n_2866),
.B(n_1247),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2870),
.B(n_2734),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2870),
.B(n_1248),
.Y(n_2916)
);

AOI21xp5_ASAP7_75t_L g2917 ( 
.A1(n_2867),
.A2(n_1250),
.B(n_1249),
.Y(n_2917)
);

OAI22xp5_ASAP7_75t_L g2918 ( 
.A1(n_2868),
.A2(n_1278),
.B1(n_1281),
.B2(n_1274),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2850),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2893),
.B(n_2888),
.Y(n_2920)
);

AND2x2_ASAP7_75t_L g2921 ( 
.A(n_2888),
.B(n_2912),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2909),
.B(n_2846),
.Y(n_2922)
);

BUFx6f_ASAP7_75t_L g2923 ( 
.A(n_2883),
.Y(n_2923)
);

NAND5xp2_ASAP7_75t_L g2924 ( 
.A(n_2880),
.B(n_2858),
.C(n_2856),
.D(n_2852),
.E(n_2874),
.Y(n_2924)
);

AO21x2_ASAP7_75t_L g2925 ( 
.A1(n_2910),
.A2(n_2845),
.B(n_2856),
.Y(n_2925)
);

AND2x2_ASAP7_75t_L g2926 ( 
.A(n_2913),
.B(n_2858),
.Y(n_2926)
);

AOI222xp33_ASAP7_75t_L g2927 ( 
.A1(n_2891),
.A2(n_1299),
.B1(n_1295),
.B2(n_1304),
.C1(n_1296),
.C2(n_1288),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2890),
.Y(n_2928)
);

BUFx3_ASAP7_75t_L g2929 ( 
.A(n_2892),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2919),
.B(n_2849),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2881),
.Y(n_2931)
);

INVxp67_ASAP7_75t_SL g2932 ( 
.A(n_2885),
.Y(n_2932)
);

INVx5_ASAP7_75t_L g2933 ( 
.A(n_2889),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2899),
.Y(n_2934)
);

BUFx3_ASAP7_75t_L g2935 ( 
.A(n_2883),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2898),
.B(n_2848),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2886),
.Y(n_2937)
);

AND2x2_ASAP7_75t_L g2938 ( 
.A(n_2906),
.B(n_2848),
.Y(n_2938)
);

INVxp67_ASAP7_75t_SL g2939 ( 
.A(n_2904),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2905),
.Y(n_2940)
);

OR2x2_ASAP7_75t_L g2941 ( 
.A(n_2894),
.B(n_2854),
.Y(n_2941)
);

INVx2_ASAP7_75t_SL g2942 ( 
.A(n_2900),
.Y(n_2942)
);

AND2x2_ASAP7_75t_L g2943 ( 
.A(n_2897),
.B(n_2908),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_2886),
.B(n_2854),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2901),
.Y(n_2945)
);

INVxp67_ASAP7_75t_SL g2946 ( 
.A(n_2882),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2886),
.Y(n_2947)
);

BUFx3_ASAP7_75t_L g2948 ( 
.A(n_2916),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2900),
.B(n_2850),
.Y(n_2949)
);

AOI211xp5_ASAP7_75t_L g2950 ( 
.A1(n_2896),
.A2(n_2902),
.B(n_2917),
.C(n_2903),
.Y(n_2950)
);

AOI221xp5_ASAP7_75t_L g2951 ( 
.A1(n_2896),
.A2(n_1312),
.B1(n_1308),
.B2(n_15),
.C(n_13),
.Y(n_2951)
);

HB1xp67_ASAP7_75t_L g2952 ( 
.A(n_2915),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2907),
.Y(n_2953)
);

AOI22xp33_ASAP7_75t_L g2954 ( 
.A1(n_2884),
.A2(n_2902),
.B1(n_2911),
.B2(n_2914),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2895),
.B(n_14),
.Y(n_2955)
);

OR2x2_ASAP7_75t_L g2956 ( 
.A(n_2932),
.B(n_2887),
.Y(n_2956)
);

AND2x4_ASAP7_75t_L g2957 ( 
.A(n_2920),
.B(n_15),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2920),
.B(n_2895),
.Y(n_2958)
);

NOR2x1_ASAP7_75t_L g2959 ( 
.A(n_2935),
.B(n_2918),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2923),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2928),
.Y(n_2961)
);

AND2x2_ASAP7_75t_L g2962 ( 
.A(n_2921),
.B(n_16),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2950),
.B(n_16),
.Y(n_2963)
);

NOR2x1_ASAP7_75t_L g2964 ( 
.A(n_2935),
.B(n_17),
.Y(n_2964)
);

INVx2_ASAP7_75t_SL g2965 ( 
.A(n_2933),
.Y(n_2965)
);

OR2x2_ASAP7_75t_L g2966 ( 
.A(n_2945),
.B(n_17),
.Y(n_2966)
);

OAI22xp5_ASAP7_75t_L g2967 ( 
.A1(n_2954),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2923),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2923),
.Y(n_2969)
);

INVx2_ASAP7_75t_SL g2970 ( 
.A(n_2933),
.Y(n_2970)
);

INVx3_ASAP7_75t_L g2971 ( 
.A(n_2923),
.Y(n_2971)
);

AND2x2_ASAP7_75t_L g2972 ( 
.A(n_2949),
.B(n_19),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2950),
.B(n_21),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2928),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2934),
.Y(n_2975)
);

NOR2x1_ASAP7_75t_SL g2976 ( 
.A(n_2925),
.B(n_23),
.Y(n_2976)
);

OR2x2_ASAP7_75t_L g2977 ( 
.A(n_2945),
.B(n_781),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2923),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2949),
.B(n_22),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2921),
.B(n_22),
.Y(n_2980)
);

AND2x4_ASAP7_75t_L g2981 ( 
.A(n_2935),
.B(n_24),
.Y(n_2981)
);

HB1xp67_ASAP7_75t_L g2982 ( 
.A(n_2941),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2934),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2926),
.B(n_24),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2946),
.B(n_25),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2933),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2926),
.B(n_26),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2948),
.B(n_27),
.Y(n_2988)
);

HB1xp67_ASAP7_75t_L g2989 ( 
.A(n_2941),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2939),
.B(n_28),
.Y(n_2990)
);

INVx1_ASAP7_75t_SL g2991 ( 
.A(n_2929),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2940),
.Y(n_2992)
);

AND2x2_ASAP7_75t_L g2993 ( 
.A(n_2942),
.B(n_28),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2948),
.B(n_30),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2933),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2940),
.Y(n_2996)
);

OR2x2_ASAP7_75t_L g2997 ( 
.A(n_2922),
.B(n_788),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2936),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2930),
.Y(n_2999)
);

AND2x2_ASAP7_75t_L g3000 ( 
.A(n_2942),
.B(n_32),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2948),
.B(n_32),
.Y(n_3001)
);

AND2x4_ASAP7_75t_SL g3002 ( 
.A(n_2957),
.B(n_2930),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2957),
.B(n_2927),
.Y(n_3003)
);

NOR3xp33_ASAP7_75t_L g3004 ( 
.A(n_2959),
.B(n_2951),
.C(n_2924),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2982),
.Y(n_3005)
);

XNOR2xp5_ASAP7_75t_L g3006 ( 
.A(n_2991),
.B(n_2929),
.Y(n_3006)
);

INVx1_ASAP7_75t_SL g3007 ( 
.A(n_2972),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2965),
.Y(n_3008)
);

INVx4_ASAP7_75t_L g3009 ( 
.A(n_2981),
.Y(n_3009)
);

NAND4xp75_ASAP7_75t_SL g3010 ( 
.A(n_2958),
.B(n_2955),
.C(n_2944),
.D(n_2943),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2957),
.B(n_2955),
.Y(n_3011)
);

NAND4xp75_ASAP7_75t_L g3012 ( 
.A(n_2964),
.B(n_2953),
.C(n_2947),
.D(n_2937),
.Y(n_3012)
);

XNOR2xp5_ASAP7_75t_L g3013 ( 
.A(n_2967),
.B(n_2929),
.Y(n_3013)
);

BUFx8_ASAP7_75t_L g3014 ( 
.A(n_2993),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2982),
.Y(n_3015)
);

NOR3xp33_ASAP7_75t_SL g3016 ( 
.A(n_2963),
.B(n_2925),
.C(n_2933),
.Y(n_3016)
);

XNOR2xp5_ASAP7_75t_L g3017 ( 
.A(n_2956),
.B(n_2943),
.Y(n_3017)
);

NAND4xp75_ASAP7_75t_SL g3018 ( 
.A(n_2990),
.B(n_2944),
.C(n_2938),
.D(n_2925),
.Y(n_3018)
);

INVx2_ASAP7_75t_SL g3019 ( 
.A(n_2965),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2989),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2973),
.B(n_2953),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2972),
.B(n_2938),
.Y(n_3022)
);

INVx2_ASAP7_75t_SL g3023 ( 
.A(n_2970),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2979),
.B(n_2952),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2989),
.Y(n_3025)
);

NOR3xp33_ASAP7_75t_SL g3026 ( 
.A(n_2998),
.B(n_2933),
.C(n_2937),
.Y(n_3026)
);

INVx3_ASAP7_75t_L g3027 ( 
.A(n_2970),
.Y(n_3027)
);

INVxp67_ASAP7_75t_SL g3028 ( 
.A(n_2976),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2979),
.B(n_2931),
.Y(n_3029)
);

NAND4xp75_ASAP7_75t_L g3030 ( 
.A(n_2990),
.B(n_2937),
.C(n_2947),
.D(n_2931),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2993),
.B(n_2947),
.Y(n_3031)
);

XOR2x2_ASAP7_75t_L g3032 ( 
.A(n_2988),
.B(n_33),
.Y(n_3032)
);

NOR3xp33_ASAP7_75t_L g3033 ( 
.A(n_2971),
.B(n_34),
.C(n_38),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2999),
.B(n_40),
.Y(n_3034)
);

NOR3xp33_ASAP7_75t_L g3035 ( 
.A(n_2971),
.B(n_40),
.C(n_41),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2971),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2960),
.Y(n_3037)
);

XNOR2xp5_ASAP7_75t_L g3038 ( 
.A(n_2962),
.B(n_41),
.Y(n_3038)
);

INVx3_ASAP7_75t_L g3039 ( 
.A(n_2986),
.Y(n_3039)
);

NAND4xp75_ASAP7_75t_SL g3040 ( 
.A(n_2980),
.B(n_2987),
.C(n_2984),
.D(n_3000),
.Y(n_3040)
);

AND2x4_ASAP7_75t_SL g3041 ( 
.A(n_2981),
.B(n_42),
.Y(n_3041)
);

AND2x2_ASAP7_75t_SL g3042 ( 
.A(n_2997),
.B(n_42),
.Y(n_3042)
);

NAND4xp75_ASAP7_75t_L g3043 ( 
.A(n_2960),
.B(n_45),
.C(n_43),
.D(n_44),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2981),
.B(n_43),
.Y(n_3044)
);

NAND3xp33_ASAP7_75t_L g3045 ( 
.A(n_2968),
.B(n_2978),
.C(n_2969),
.Y(n_3045)
);

NOR3xp33_ASAP7_75t_L g3046 ( 
.A(n_2985),
.B(n_45),
.C(n_46),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2986),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2995),
.Y(n_3048)
);

NOR2xp33_ASAP7_75t_L g3049 ( 
.A(n_2994),
.B(n_782),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2995),
.Y(n_3050)
);

XOR2xp5_ASAP7_75t_L g3051 ( 
.A(n_2966),
.B(n_46),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2968),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_2969),
.B(n_47),
.Y(n_3053)
);

XNOR2xp5_ASAP7_75t_L g3054 ( 
.A(n_3001),
.B(n_48),
.Y(n_3054)
);

NAND3xp33_ASAP7_75t_L g3055 ( 
.A(n_2978),
.B(n_51),
.C(n_50),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_2977),
.B(n_49),
.Y(n_3056)
);

AOI22xp5_ASAP7_75t_L g3057 ( 
.A1(n_2992),
.A2(n_52),
.B1(n_49),
.B2(n_50),
.Y(n_3057)
);

NAND4xp75_ASAP7_75t_L g3058 ( 
.A(n_2996),
.B(n_55),
.C(n_53),
.D(n_54),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_2961),
.B(n_56),
.Y(n_3059)
);

XNOR2xp5_ASAP7_75t_L g3060 ( 
.A(n_2974),
.B(n_57),
.Y(n_3060)
);

XOR2xp5_ASAP7_75t_L g3061 ( 
.A(n_2975),
.B(n_58),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2983),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2957),
.B(n_58),
.Y(n_3063)
);

NAND4xp75_ASAP7_75t_L g3064 ( 
.A(n_2959),
.B(n_61),
.C(n_59),
.D(n_60),
.Y(n_3064)
);

XOR2xp5_ASAP7_75t_L g3065 ( 
.A(n_2956),
.B(n_59),
.Y(n_3065)
);

NAND4xp75_ASAP7_75t_L g3066 ( 
.A(n_2959),
.B(n_64),
.C(n_62),
.D(n_63),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_SL g3067 ( 
.A(n_2991),
.B(n_62),
.Y(n_3067)
);

NAND4xp75_ASAP7_75t_SL g3068 ( 
.A(n_2958),
.B(n_65),
.C(n_63),
.D(n_64),
.Y(n_3068)
);

NOR2xp67_ASAP7_75t_L g3069 ( 
.A(n_3009),
.B(n_785),
.Y(n_3069)
);

INVx3_ASAP7_75t_SL g3070 ( 
.A(n_3041),
.Y(n_3070)
);

INVxp67_ASAP7_75t_L g3071 ( 
.A(n_3014),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_3025),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_3022),
.B(n_786),
.Y(n_3073)
);

INVx2_ASAP7_75t_SL g3074 ( 
.A(n_3002),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_3025),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_3005),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_3028),
.B(n_65),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_3015),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_3020),
.Y(n_3079)
);

AND2x2_ASAP7_75t_L g3080 ( 
.A(n_3007),
.B(n_3006),
.Y(n_3080)
);

AND2x2_ASAP7_75t_L g3081 ( 
.A(n_3042),
.B(n_789),
.Y(n_3081)
);

NAND4xp75_ASAP7_75t_L g3082 ( 
.A(n_3016),
.B(n_68),
.C(n_66),
.D(n_67),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_3037),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_3014),
.Y(n_3084)
);

OR2x2_ASAP7_75t_L g3085 ( 
.A(n_3011),
.B(n_67),
.Y(n_3085)
);

OAI211xp5_ASAP7_75t_SL g3086 ( 
.A1(n_3004),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_3086)
);

NOR2xp33_ASAP7_75t_L g3087 ( 
.A(n_3065),
.B(n_772),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_3052),
.Y(n_3088)
);

OR2x2_ASAP7_75t_L g3089 ( 
.A(n_3024),
.B(n_3029),
.Y(n_3089)
);

AOI221xp5_ASAP7_75t_L g3090 ( 
.A1(n_3021),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.C(n_72),
.Y(n_3090)
);

NOR2xp33_ASAP7_75t_L g3091 ( 
.A(n_3009),
.B(n_777),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_3017),
.B(n_777),
.Y(n_3092)
);

INVx1_ASAP7_75t_SL g3093 ( 
.A(n_3040),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_3064),
.B(n_73),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_3066),
.B(n_74),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_3046),
.B(n_74),
.Y(n_3096)
);

AND2x4_ASAP7_75t_L g3097 ( 
.A(n_3027),
.B(n_78),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_3053),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_3034),
.B(n_780),
.Y(n_3099)
);

AND2x4_ASAP7_75t_L g3100 ( 
.A(n_3027),
.B(n_78),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_3019),
.B(n_76),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_3008),
.B(n_782),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_3039),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_3039),
.Y(n_3104)
);

OR2x2_ASAP7_75t_L g3105 ( 
.A(n_3003),
.B(n_76),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_3023),
.B(n_784),
.Y(n_3106)
);

AND2x2_ASAP7_75t_L g3107 ( 
.A(n_3013),
.B(n_787),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_SL g3108 ( 
.A(n_3055),
.B(n_79),
.Y(n_3108)
);

AND2x2_ASAP7_75t_L g3109 ( 
.A(n_3056),
.B(n_787),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_3026),
.B(n_789),
.Y(n_3110)
);

O2A1O1Ixp33_ASAP7_75t_SL g3111 ( 
.A1(n_3067),
.A2(n_3031),
.B(n_3063),
.C(n_3044),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_3045),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_3036),
.B(n_790),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_3047),
.Y(n_3114)
);

AOI31xp33_ASAP7_75t_L g3115 ( 
.A1(n_3038),
.A2(n_81),
.A3(n_79),
.B(n_80),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_3048),
.Y(n_3116)
);

AND2x4_ASAP7_75t_L g3117 ( 
.A(n_3050),
.B(n_82),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_3033),
.B(n_81),
.Y(n_3118)
);

AND2x2_ASAP7_75t_L g3119 ( 
.A(n_3059),
.B(n_3032),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_3030),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_3062),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_3049),
.B(n_766),
.Y(n_3122)
);

OR2x2_ASAP7_75t_L g3123 ( 
.A(n_3012),
.B(n_82),
.Y(n_3123)
);

AND2x2_ASAP7_75t_L g3124 ( 
.A(n_3051),
.B(n_768),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_3035),
.B(n_84),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_3054),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_3043),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_3060),
.Y(n_3128)
);

OR2x2_ASAP7_75t_L g3129 ( 
.A(n_3061),
.B(n_84),
.Y(n_3129)
);

INVx2_ASAP7_75t_L g3130 ( 
.A(n_3058),
.Y(n_3130)
);

OR2x2_ASAP7_75t_L g3131 ( 
.A(n_3057),
.B(n_3010),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_3018),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_3068),
.Y(n_3133)
);

INVx1_ASAP7_75t_SL g3134 ( 
.A(n_3002),
.Y(n_3134)
);

OR2x2_ASAP7_75t_L g3135 ( 
.A(n_3007),
.B(n_85),
.Y(n_3135)
);

OR2x2_ASAP7_75t_L g3136 ( 
.A(n_3007),
.B(n_85),
.Y(n_3136)
);

AND2x2_ASAP7_75t_L g3137 ( 
.A(n_3022),
.B(n_770),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_3028),
.B(n_86),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_3025),
.Y(n_3139)
);

INVx1_ASAP7_75t_SL g3140 ( 
.A(n_3002),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_3022),
.B(n_771),
.Y(n_3141)
);

OR2x2_ASAP7_75t_L g3142 ( 
.A(n_3007),
.B(n_87),
.Y(n_3142)
);

HB1xp67_ASAP7_75t_L g3143 ( 
.A(n_3014),
.Y(n_3143)
);

OR2x2_ASAP7_75t_L g3144 ( 
.A(n_3007),
.B(n_88),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_3025),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_3025),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_3025),
.Y(n_3147)
);

NOR2x1_ASAP7_75t_R g3148 ( 
.A(n_3028),
.B(n_88),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_3014),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_3025),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_3022),
.B(n_775),
.Y(n_3151)
);

OR2x2_ASAP7_75t_L g3152 ( 
.A(n_3007),
.B(n_89),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_3022),
.B(n_778),
.Y(n_3153)
);

NOR2xp33_ASAP7_75t_L g3154 ( 
.A(n_3065),
.B(n_779),
.Y(n_3154)
);

INVx1_ASAP7_75t_SL g3155 ( 
.A(n_3002),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_3014),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_3025),
.Y(n_3157)
);

NOR2x1_ASAP7_75t_L g3158 ( 
.A(n_3064),
.B(n_90),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_3028),
.B(n_91),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_3025),
.Y(n_3160)
);

AND2x4_ASAP7_75t_SL g3161 ( 
.A(n_3009),
.B(n_91),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_3143),
.B(n_92),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_3072),
.Y(n_3163)
);

AOI211xp5_ASAP7_75t_L g3164 ( 
.A1(n_3086),
.A2(n_95),
.B(n_92),
.C(n_93),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_3072),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_3070),
.B(n_93),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_3145),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_3145),
.Y(n_3168)
);

AOI22xp5_ASAP7_75t_L g3169 ( 
.A1(n_3112),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_3169)
);

AOI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_3111),
.A2(n_96),
.B(n_99),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_3084),
.B(n_100),
.Y(n_3171)
);

A2O1A1Ixp33_ASAP7_75t_L g3172 ( 
.A1(n_3158),
.A2(n_102),
.B(n_100),
.C(n_101),
.Y(n_3172)
);

INVx1_ASAP7_75t_SL g3173 ( 
.A(n_3134),
.Y(n_3173)
);

INVx3_ASAP7_75t_L g3174 ( 
.A(n_3097),
.Y(n_3174)
);

XOR2xp5_ASAP7_75t_L g3175 ( 
.A(n_3149),
.B(n_3156),
.Y(n_3175)
);

AO21x1_ASAP7_75t_L g3176 ( 
.A1(n_3123),
.A2(n_3112),
.B(n_3115),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_3140),
.B(n_102),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3157),
.Y(n_3178)
);

A2O1A1Ixp33_ASAP7_75t_L g3179 ( 
.A1(n_3120),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_3157),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_3155),
.B(n_103),
.Y(n_3181)
);

NAND3xp33_ASAP7_75t_L g3182 ( 
.A(n_3071),
.B(n_104),
.C(n_105),
.Y(n_3182)
);

AOI22xp33_ASAP7_75t_SL g3183 ( 
.A1(n_3093),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_3183)
);

OAI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_3082),
.A2(n_106),
.B(n_107),
.Y(n_3184)
);

NOR2x1_ASAP7_75t_L g3185 ( 
.A(n_3069),
.B(n_108),
.Y(n_3185)
);

OR2x2_ASAP7_75t_L g3186 ( 
.A(n_3130),
.B(n_110),
.Y(n_3186)
);

O2A1O1Ixp5_ASAP7_75t_L g3187 ( 
.A1(n_3104),
.A2(n_114),
.B(n_111),
.C(n_113),
.Y(n_3187)
);

INVx2_ASAP7_75t_L g3188 ( 
.A(n_3161),
.Y(n_3188)
);

XOR2x2_ASAP7_75t_L g3189 ( 
.A(n_3119),
.B(n_111),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_3160),
.Y(n_3190)
);

OAI21x1_ASAP7_75t_L g3191 ( 
.A1(n_3103),
.A2(n_113),
.B(n_116),
.Y(n_3191)
);

OAI22xp5_ASAP7_75t_L g3192 ( 
.A1(n_3131),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_3192)
);

OAI22xp5_ASAP7_75t_L g3193 ( 
.A1(n_3127),
.A2(n_121),
.B1(n_117),
.B2(n_120),
.Y(n_3193)
);

NOR3xp33_ASAP7_75t_L g3194 ( 
.A(n_3080),
.B(n_120),
.C(n_122),
.Y(n_3194)
);

OAI21xp33_ASAP7_75t_SL g3195 ( 
.A1(n_3074),
.A2(n_3103),
.B(n_3110),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_3160),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3075),
.Y(n_3197)
);

AOI21xp5_ASAP7_75t_L g3198 ( 
.A1(n_3108),
.A2(n_122),
.B(n_123),
.Y(n_3198)
);

AOI22xp5_ASAP7_75t_L g3199 ( 
.A1(n_3092),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_3199)
);

OAI22xp33_ASAP7_75t_L g3200 ( 
.A1(n_3096),
.A2(n_128),
.B1(n_125),
.B2(n_127),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_3148),
.B(n_128),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_3073),
.B(n_129),
.Y(n_3202)
);

INVxp67_ASAP7_75t_L g3203 ( 
.A(n_3081),
.Y(n_3203)
);

OAI21xp33_ASAP7_75t_L g3204 ( 
.A1(n_3132),
.A2(n_130),
.B(n_131),
.Y(n_3204)
);

AOI22x1_ASAP7_75t_L g3205 ( 
.A1(n_3098),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_3205)
);

XOR2x2_ASAP7_75t_L g3206 ( 
.A(n_3126),
.B(n_132),
.Y(n_3206)
);

OAI22x1_ASAP7_75t_L g3207 ( 
.A1(n_3133),
.A2(n_136),
.B1(n_133),
.B2(n_135),
.Y(n_3207)
);

OAI22xp33_ASAP7_75t_SL g3208 ( 
.A1(n_3076),
.A2(n_766),
.B1(n_768),
.B2(n_765),
.Y(n_3208)
);

AOI22xp5_ASAP7_75t_L g3209 ( 
.A1(n_3107),
.A2(n_138),
.B1(n_135),
.B2(n_137),
.Y(n_3209)
);

AOI22xp5_ASAP7_75t_L g3210 ( 
.A1(n_3128),
.A2(n_140),
.B1(n_137),
.B2(n_138),
.Y(n_3210)
);

OAI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_3077),
.A2(n_142),
.B(n_143),
.Y(n_3211)
);

INVxp67_ASAP7_75t_SL g3212 ( 
.A(n_3138),
.Y(n_3212)
);

AND2x2_ASAP7_75t_L g3213 ( 
.A(n_3137),
.B(n_143),
.Y(n_3213)
);

OAI22xp33_ASAP7_75t_L g3214 ( 
.A1(n_3118),
.A2(n_147),
.B1(n_144),
.B2(n_146),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3139),
.Y(n_3215)
);

INVxp67_ASAP7_75t_L g3216 ( 
.A(n_3091),
.Y(n_3216)
);

OAI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_3159),
.A2(n_146),
.B(n_149),
.Y(n_3217)
);

OAI22xp5_ASAP7_75t_L g3218 ( 
.A1(n_3089),
.A2(n_152),
.B1(n_149),
.B2(n_151),
.Y(n_3218)
);

XOR2x2_ASAP7_75t_L g3219 ( 
.A(n_3090),
.B(n_152),
.Y(n_3219)
);

OAI31xp33_ASAP7_75t_SL g3220 ( 
.A1(n_3078),
.A2(n_156),
.A3(n_154),
.B(n_155),
.Y(n_3220)
);

OAI22xp5_ASAP7_75t_L g3221 ( 
.A1(n_3094),
.A2(n_157),
.B1(n_154),
.B2(n_155),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_3097),
.Y(n_3222)
);

OAI21xp5_ASAP7_75t_L g3223 ( 
.A1(n_3125),
.A2(n_158),
.B(n_159),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_3141),
.B(n_159),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_3151),
.B(n_160),
.Y(n_3225)
);

BUFx2_ASAP7_75t_L g3226 ( 
.A(n_3100),
.Y(n_3226)
);

AOI22xp5_ASAP7_75t_L g3227 ( 
.A1(n_3079),
.A2(n_3100),
.B1(n_3106),
.B2(n_3153),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_3117),
.Y(n_3228)
);

AOI22xp5_ASAP7_75t_L g3229 ( 
.A1(n_3102),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_3229)
);

OAI22xp5_ASAP7_75t_L g3230 ( 
.A1(n_3095),
.A2(n_164),
.B1(n_161),
.B2(n_163),
.Y(n_3230)
);

OAI21xp33_ASAP7_75t_L g3231 ( 
.A1(n_3114),
.A2(n_163),
.B(n_165),
.Y(n_3231)
);

INVxp67_ASAP7_75t_SL g3232 ( 
.A(n_3087),
.Y(n_3232)
);

AOI21xp5_ASAP7_75t_L g3233 ( 
.A1(n_3105),
.A2(n_165),
.B(n_166),
.Y(n_3233)
);

AOI22xp5_ASAP7_75t_L g3234 ( 
.A1(n_3116),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_3234)
);

AOI22xp33_ASAP7_75t_SL g3235 ( 
.A1(n_3146),
.A2(n_172),
.B1(n_168),
.B2(n_171),
.Y(n_3235)
);

NAND3xp33_ASAP7_75t_L g3236 ( 
.A(n_3121),
.B(n_171),
.C(n_172),
.Y(n_3236)
);

AOI22xp33_ASAP7_75t_L g3237 ( 
.A1(n_3147),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_3237)
);

INVxp67_ASAP7_75t_SL g3238 ( 
.A(n_3154),
.Y(n_3238)
);

AOI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_3101),
.A2(n_173),
.B(n_174),
.Y(n_3239)
);

NAND3xp33_ASAP7_75t_L g3240 ( 
.A(n_3150),
.B(n_175),
.C(n_176),
.Y(n_3240)
);

OAI22xp33_ASAP7_75t_L g3241 ( 
.A1(n_3135),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_3241)
);

INVxp33_ASAP7_75t_L g3242 ( 
.A(n_3122),
.Y(n_3242)
);

XNOR2x1_ASAP7_75t_L g3243 ( 
.A(n_3129),
.B(n_177),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3113),
.B(n_3109),
.Y(n_3244)
);

OAI221xp5_ASAP7_75t_L g3245 ( 
.A1(n_3085),
.A2(n_182),
.B1(n_179),
.B2(n_181),
.C(n_183),
.Y(n_3245)
);

OAI211xp5_ASAP7_75t_L g3246 ( 
.A1(n_3083),
.A2(n_184),
.B(n_181),
.C(n_183),
.Y(n_3246)
);

NOR3x1_ASAP7_75t_L g3247 ( 
.A(n_3136),
.B(n_186),
.C(n_187),
.Y(n_3247)
);

AND2x2_ASAP7_75t_L g3248 ( 
.A(n_3099),
.B(n_186),
.Y(n_3248)
);

INVx2_ASAP7_75t_SL g3249 ( 
.A(n_3117),
.Y(n_3249)
);

AOI22xp5_ASAP7_75t_L g3250 ( 
.A1(n_3088),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3142),
.Y(n_3251)
);

OAI22xp33_ASAP7_75t_L g3252 ( 
.A1(n_3152),
.A2(n_192),
.B1(n_188),
.B2(n_190),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3144),
.Y(n_3253)
);

INVx4_ASAP7_75t_L g3254 ( 
.A(n_3124),
.Y(n_3254)
);

OAI221xp5_ASAP7_75t_L g3255 ( 
.A1(n_3071),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.C(n_196),
.Y(n_3255)
);

INVx1_ASAP7_75t_SL g3256 ( 
.A(n_3070),
.Y(n_3256)
);

AND2x2_ASAP7_75t_L g3257 ( 
.A(n_3143),
.B(n_193),
.Y(n_3257)
);

XOR2x2_ASAP7_75t_L g3258 ( 
.A(n_3082),
.B(n_196),
.Y(n_3258)
);

INVxp67_ASAP7_75t_L g3259 ( 
.A(n_3148),
.Y(n_3259)
);

INVxp67_ASAP7_75t_L g3260 ( 
.A(n_3148),
.Y(n_3260)
);

OR4x1_ASAP7_75t_L g3261 ( 
.A(n_3074),
.B(n_199),
.C(n_197),
.D(n_198),
.Y(n_3261)
);

AOI21xp33_ASAP7_75t_L g3262 ( 
.A1(n_3071),
.A2(n_772),
.B(n_770),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3072),
.Y(n_3263)
);

AOI21xp33_ASAP7_75t_SL g3264 ( 
.A1(n_3070),
.A2(n_197),
.B(n_198),
.Y(n_3264)
);

OAI211xp5_ASAP7_75t_L g3265 ( 
.A1(n_3112),
.A2(n_201),
.B(n_199),
.C(n_200),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3072),
.Y(n_3266)
);

AOI22xp5_ASAP7_75t_L g3267 ( 
.A1(n_3112),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_3267)
);

INVx1_ASAP7_75t_SL g3268 ( 
.A(n_3070),
.Y(n_3268)
);

AOI22xp5_ASAP7_75t_L g3269 ( 
.A1(n_3112),
.A2(n_206),
.B1(n_202),
.B2(n_205),
.Y(n_3269)
);

OAI21xp33_ASAP7_75t_L g3270 ( 
.A1(n_3071),
.A2(n_207),
.B(n_208),
.Y(n_3270)
);

AOI211xp5_ASAP7_75t_L g3271 ( 
.A1(n_3086),
.A2(n_212),
.B(n_209),
.C(n_211),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3072),
.Y(n_3272)
);

INVxp67_ASAP7_75t_L g3273 ( 
.A(n_3148),
.Y(n_3273)
);

HB1xp67_ASAP7_75t_L g3274 ( 
.A(n_3069),
.Y(n_3274)
);

INVx1_ASAP7_75t_SL g3275 ( 
.A(n_3070),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3072),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3072),
.Y(n_3277)
);

OAI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_3082),
.A2(n_211),
.B(n_212),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3072),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3072),
.Y(n_3280)
);

NOR2xp33_ASAP7_75t_L g3281 ( 
.A(n_3070),
.B(n_214),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_3143),
.B(n_215),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_3084),
.Y(n_3283)
);

XNOR2xp5_ASAP7_75t_L g3284 ( 
.A(n_3143),
.B(n_774),
.Y(n_3284)
);

AOI22xp33_ASAP7_75t_L g3285 ( 
.A1(n_3112),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3072),
.Y(n_3286)
);

AOI22xp5_ASAP7_75t_L g3287 ( 
.A1(n_3112),
.A2(n_220),
.B1(n_217),
.B2(n_218),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3072),
.Y(n_3288)
);

AOI22xp5_ASAP7_75t_L g3289 ( 
.A1(n_3112),
.A2(n_222),
.B1(n_218),
.B2(n_221),
.Y(n_3289)
);

AOI22xp5_ASAP7_75t_L g3290 ( 
.A1(n_3112),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_3072),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3072),
.Y(n_3292)
);

AOI22xp5_ASAP7_75t_L g3293 ( 
.A1(n_3112),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_3111),
.A2(n_228),
.B(n_229),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3072),
.Y(n_3295)
);

INVxp67_ASAP7_75t_L g3296 ( 
.A(n_3148),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3143),
.B(n_228),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3072),
.Y(n_3298)
);

NOR3xp33_ASAP7_75t_L g3299 ( 
.A(n_3071),
.B(n_230),
.C(n_231),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3072),
.Y(n_3300)
);

XNOR2x1_ASAP7_75t_L g3301 ( 
.A(n_3082),
.B(n_230),
.Y(n_3301)
);

OAI22xp5_ASAP7_75t_L g3302 ( 
.A1(n_3082),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_3302)
);

NAND3xp33_ASAP7_75t_L g3303 ( 
.A(n_3112),
.B(n_233),
.C(n_234),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3072),
.Y(n_3304)
);

OR2x2_ASAP7_75t_L g3305 ( 
.A(n_3130),
.B(n_234),
.Y(n_3305)
);

OR2x2_ASAP7_75t_L g3306 ( 
.A(n_3130),
.B(n_235),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3084),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_3072),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3072),
.Y(n_3309)
);

OAI22xp33_ASAP7_75t_R g3310 ( 
.A1(n_3093),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_3310)
);

XNOR2xp5_ASAP7_75t_L g3311 ( 
.A(n_3143),
.B(n_783),
.Y(n_3311)
);

BUFx3_ASAP7_75t_L g3312 ( 
.A(n_3070),
.Y(n_3312)
);

OAI22xp33_ASAP7_75t_L g3313 ( 
.A1(n_3112),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_3313)
);

AOI211xp5_ASAP7_75t_SL g3314 ( 
.A1(n_3071),
.A2(n_242),
.B(n_239),
.C(n_241),
.Y(n_3314)
);

OA22x2_ASAP7_75t_L g3315 ( 
.A1(n_3112),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_3315)
);

AOI22xp5_ASAP7_75t_L g3316 ( 
.A1(n_3112),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_3316)
);

AOI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_3112),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.Y(n_3317)
);

OAI22xp5_ASAP7_75t_L g3318 ( 
.A1(n_3256),
.A2(n_250),
.B1(n_247),
.B2(n_248),
.Y(n_3318)
);

OR2x2_ASAP7_75t_L g3319 ( 
.A(n_3274),
.B(n_250),
.Y(n_3319)
);

OR2x2_ASAP7_75t_L g3320 ( 
.A(n_3173),
.B(n_251),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3268),
.B(n_251),
.Y(n_3321)
);

OR2x2_ASAP7_75t_L g3322 ( 
.A(n_3249),
.B(n_252),
.Y(n_3322)
);

OR2x2_ASAP7_75t_L g3323 ( 
.A(n_3226),
.B(n_254),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3275),
.B(n_255),
.Y(n_3324)
);

AND2x2_ASAP7_75t_L g3325 ( 
.A(n_3312),
.B(n_257),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3185),
.Y(n_3326)
);

AOI31xp33_ASAP7_75t_L g3327 ( 
.A1(n_3259),
.A2(n_790),
.A3(n_259),
.B(n_257),
.Y(n_3327)
);

INVxp67_ASAP7_75t_L g3328 ( 
.A(n_3175),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_3174),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_3260),
.B(n_258),
.Y(n_3330)
);

OAI22xp33_ASAP7_75t_L g3331 ( 
.A1(n_3314),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_3331)
);

OAI32xp33_ASAP7_75t_L g3332 ( 
.A1(n_3195),
.A2(n_263),
.A3(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_3332)
);

NAND4xp75_ASAP7_75t_L g3333 ( 
.A(n_3176),
.B(n_267),
.C(n_265),
.D(n_266),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3257),
.Y(n_3334)
);

AOI211xp5_ASAP7_75t_SL g3335 ( 
.A1(n_3273),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_3335)
);

INVx2_ASAP7_75t_SL g3336 ( 
.A(n_3174),
.Y(n_3336)
);

INVxp67_ASAP7_75t_L g3337 ( 
.A(n_3281),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3284),
.Y(n_3338)
);

AND2x2_ASAP7_75t_L g3339 ( 
.A(n_3296),
.B(n_269),
.Y(n_3339)
);

INVx2_ASAP7_75t_SL g3340 ( 
.A(n_3222),
.Y(n_3340)
);

AND2x4_ASAP7_75t_L g3341 ( 
.A(n_3188),
.B(n_269),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3311),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_3254),
.B(n_272),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3166),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3283),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3307),
.B(n_272),
.Y(n_3346)
);

INVx2_ASAP7_75t_L g3347 ( 
.A(n_3254),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3228),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3177),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3181),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3162),
.Y(n_3351)
);

OAI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_3170),
.A2(n_273),
.B(n_274),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3171),
.Y(n_3353)
);

A2O1A1Ixp33_ASAP7_75t_SL g3354 ( 
.A1(n_3216),
.A2(n_277),
.B(n_274),
.C(n_275),
.Y(n_3354)
);

INVxp67_ASAP7_75t_SL g3355 ( 
.A(n_3247),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_3203),
.B(n_275),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3294),
.A2(n_278),
.B(n_279),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3282),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3264),
.B(n_279),
.Y(n_3359)
);

OAI221xp5_ASAP7_75t_L g3360 ( 
.A1(n_3220),
.A2(n_283),
.B1(n_280),
.B2(n_281),
.C(n_284),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_3248),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3183),
.B(n_3172),
.Y(n_3362)
);

OR2x2_ASAP7_75t_L g3363 ( 
.A(n_3244),
.B(n_281),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3242),
.B(n_3232),
.Y(n_3364)
);

OAI221xp5_ASAP7_75t_SL g3365 ( 
.A1(n_3227),
.A2(n_289),
.B1(n_284),
.B2(n_287),
.C(n_291),
.Y(n_3365)
);

HB1xp67_ASAP7_75t_L g3366 ( 
.A(n_3243),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3297),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3213),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3238),
.B(n_287),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3163),
.Y(n_3370)
);

HB1xp67_ASAP7_75t_L g3371 ( 
.A(n_3207),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3189),
.B(n_289),
.Y(n_3372)
);

OAI22xp33_ASAP7_75t_L g3373 ( 
.A1(n_3184),
.A2(n_294),
.B1(n_291),
.B2(n_293),
.Y(n_3373)
);

AOI221xp5_ASAP7_75t_L g3374 ( 
.A1(n_3192),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.C(n_298),
.Y(n_3374)
);

HB1xp67_ASAP7_75t_L g3375 ( 
.A(n_3315),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3165),
.Y(n_3376)
);

AND2x4_ASAP7_75t_L g3377 ( 
.A(n_3251),
.B(n_297),
.Y(n_3377)
);

AOI221xp5_ASAP7_75t_L g3378 ( 
.A1(n_3302),
.A2(n_301),
.B1(n_298),
.B2(n_300),
.C(n_302),
.Y(n_3378)
);

OAI322xp33_ASAP7_75t_L g3379 ( 
.A1(n_3197),
.A2(n_306),
.A3(n_305),
.B1(n_303),
.B2(n_300),
.C1(n_301),
.C2(n_304),
.Y(n_3379)
);

NOR2xp33_ASAP7_75t_L g3380 ( 
.A(n_3204),
.B(n_303),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3278),
.B(n_304),
.Y(n_3381)
);

AOI21xp33_ASAP7_75t_SL g3382 ( 
.A1(n_3301),
.A2(n_3194),
.B(n_3253),
.Y(n_3382)
);

NAND3xp33_ASAP7_75t_L g3383 ( 
.A(n_3303),
.B(n_305),
.C(n_307),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3167),
.Y(n_3384)
);

AOI211x1_ASAP7_75t_L g3385 ( 
.A1(n_3265),
.A2(n_310),
.B(n_307),
.C(n_309),
.Y(n_3385)
);

AOI22xp5_ASAP7_75t_L g3386 ( 
.A1(n_3310),
.A2(n_312),
.B1(n_309),
.B2(n_311),
.Y(n_3386)
);

A2O1A1Ixp33_ASAP7_75t_L g3387 ( 
.A1(n_3187),
.A2(n_314),
.B(n_311),
.C(n_313),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3168),
.Y(n_3388)
);

AOI21xp33_ASAP7_75t_L g3389 ( 
.A1(n_3212),
.A2(n_3215),
.B(n_3186),
.Y(n_3389)
);

OAI21xp33_ASAP7_75t_L g3390 ( 
.A1(n_3206),
.A2(n_3180),
.B(n_3178),
.Y(n_3390)
);

AOI22xp33_ASAP7_75t_L g3391 ( 
.A1(n_3219),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3190),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3299),
.B(n_315),
.Y(n_3393)
);

AND2x2_ASAP7_75t_L g3394 ( 
.A(n_3211),
.B(n_316),
.Y(n_3394)
);

NOR2x1_ASAP7_75t_L g3395 ( 
.A(n_3182),
.B(n_781),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3196),
.Y(n_3396)
);

AND2x4_ASAP7_75t_L g3397 ( 
.A(n_3263),
.B(n_316),
.Y(n_3397)
);

AOI22xp5_ASAP7_75t_L g3398 ( 
.A1(n_3221),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3266),
.Y(n_3399)
);

AND2x2_ASAP7_75t_L g3400 ( 
.A(n_3217),
.B(n_318),
.Y(n_3400)
);

AOI221x1_ASAP7_75t_L g3401 ( 
.A1(n_3179),
.A2(n_3208),
.B1(n_3233),
.B2(n_3239),
.C(n_3230),
.Y(n_3401)
);

INVx2_ASAP7_75t_SL g3402 ( 
.A(n_3191),
.Y(n_3402)
);

AOI22xp5_ASAP7_75t_L g3403 ( 
.A1(n_3258),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3272),
.Y(n_3404)
);

AO22x2_ASAP7_75t_L g3405 ( 
.A1(n_3276),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.Y(n_3405)
);

OAI222xp33_ASAP7_75t_L g3406 ( 
.A1(n_3205),
.A2(n_325),
.B1(n_327),
.B2(n_323),
.C1(n_324),
.C2(n_326),
.Y(n_3406)
);

OAI21xp33_ASAP7_75t_L g3407 ( 
.A1(n_3277),
.A2(n_324),
.B(n_325),
.Y(n_3407)
);

OAI21xp33_ASAP7_75t_L g3408 ( 
.A1(n_3279),
.A2(n_326),
.B(n_328),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3280),
.Y(n_3409)
);

OAI31xp33_ASAP7_75t_L g3410 ( 
.A1(n_3246),
.A2(n_3200),
.A3(n_3214),
.B(n_3313),
.Y(n_3410)
);

AOI22xp5_ASAP7_75t_L g3411 ( 
.A1(n_3164),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_3411)
);

OAI21xp33_ASAP7_75t_L g3412 ( 
.A1(n_3286),
.A2(n_329),
.B(n_330),
.Y(n_3412)
);

AOI21xp33_ASAP7_75t_L g3413 ( 
.A1(n_3305),
.A2(n_331),
.B(n_332),
.Y(n_3413)
);

OAI22xp5_ASAP7_75t_L g3414 ( 
.A1(n_3285),
.A2(n_335),
.B1(n_331),
.B2(n_334),
.Y(n_3414)
);

OAI32xp33_ASAP7_75t_L g3415 ( 
.A1(n_3288),
.A2(n_338),
.A3(n_336),
.B1(n_337),
.B2(n_339),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3291),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3292),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_SL g3418 ( 
.A(n_3271),
.B(n_336),
.Y(n_3418)
);

AOI22xp33_ASAP7_75t_SL g3419 ( 
.A1(n_3295),
.A2(n_779),
.B1(n_340),
.B2(n_338),
.Y(n_3419)
);

AOI221xp5_ASAP7_75t_L g3420 ( 
.A1(n_3298),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.C(n_342),
.Y(n_3420)
);

AOI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_3270),
.A2(n_345),
.B1(n_342),
.B2(n_344),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3300),
.Y(n_3422)
);

NAND3xp33_ASAP7_75t_L g3423 ( 
.A(n_3235),
.B(n_345),
.C(n_346),
.Y(n_3423)
);

AOI21xp5_ASAP7_75t_L g3424 ( 
.A1(n_3198),
.A2(n_346),
.B(n_347),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_3223),
.B(n_347),
.Y(n_3425)
);

AOI322xp5_ASAP7_75t_L g3426 ( 
.A1(n_3304),
.A2(n_354),
.A3(n_353),
.B1(n_351),
.B2(n_349),
.C1(n_350),
.C2(n_352),
.Y(n_3426)
);

AOI21xp33_ASAP7_75t_L g3427 ( 
.A1(n_3306),
.A2(n_3309),
.B(n_3308),
.Y(n_3427)
);

OR2x2_ASAP7_75t_L g3428 ( 
.A(n_3201),
.B(n_349),
.Y(n_3428)
);

AOI221xp5_ASAP7_75t_L g3429 ( 
.A1(n_3261),
.A2(n_358),
.B1(n_354),
.B2(n_356),
.C(n_359),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3202),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3224),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3225),
.Y(n_3432)
);

INVx2_ASAP7_75t_SL g3433 ( 
.A(n_3236),
.Y(n_3433)
);

OAI22xp5_ASAP7_75t_L g3434 ( 
.A1(n_3169),
.A2(n_360),
.B1(n_356),
.B2(n_358),
.Y(n_3434)
);

AOI22xp5_ASAP7_75t_L g3435 ( 
.A1(n_3231),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_3435)
);

NAND2xp33_ASAP7_75t_SL g3436 ( 
.A(n_3218),
.B(n_361),
.Y(n_3436)
);

OR2x2_ASAP7_75t_L g3437 ( 
.A(n_3240),
.B(n_363),
.Y(n_3437)
);

AOI222xp33_ASAP7_75t_L g3438 ( 
.A1(n_3193),
.A2(n_366),
.B1(n_368),
.B2(n_364),
.C1(n_365),
.C2(n_367),
.Y(n_3438)
);

OAI22xp5_ASAP7_75t_L g3439 ( 
.A1(n_3267),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_3439)
);

NOR2xp33_ASAP7_75t_L g3440 ( 
.A(n_3262),
.B(n_369),
.Y(n_3440)
);

INVx1_ASAP7_75t_SL g3441 ( 
.A(n_3209),
.Y(n_3441)
);

OAI21xp33_ASAP7_75t_L g3442 ( 
.A1(n_3269),
.A2(n_369),
.B(n_370),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3326),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3323),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3336),
.Y(n_3445)
);

OAI21xp5_ASAP7_75t_L g3446 ( 
.A1(n_3328),
.A2(n_3289),
.B(n_3287),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_3355),
.B(n_3241),
.Y(n_3447)
);

OAI211xp5_ASAP7_75t_SL g3448 ( 
.A1(n_3390),
.A2(n_3293),
.B(n_3316),
.C(n_3290),
.Y(n_3448)
);

AND2x2_ASAP7_75t_L g3449 ( 
.A(n_3321),
.B(n_3210),
.Y(n_3449)
);

NAND2xp33_ASAP7_75t_SL g3450 ( 
.A(n_3402),
.B(n_3237),
.Y(n_3450)
);

OAI32xp33_ASAP7_75t_L g3451 ( 
.A1(n_3375),
.A2(n_3255),
.A3(n_3245),
.B1(n_3317),
.B2(n_3252),
.Y(n_3451)
);

NOR3xp33_ASAP7_75t_L g3452 ( 
.A(n_3382),
.B(n_3199),
.C(n_3229),
.Y(n_3452)
);

AOI22xp5_ASAP7_75t_L g3453 ( 
.A1(n_3340),
.A2(n_3234),
.B1(n_3250),
.B2(n_378),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_3357),
.A2(n_374),
.B(n_377),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3324),
.Y(n_3455)
);

NAND2x1p5_ASAP7_75t_L g3456 ( 
.A(n_3325),
.B(n_374),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3329),
.B(n_377),
.Y(n_3457)
);

AOI21xp33_ASAP7_75t_SL g3458 ( 
.A1(n_3331),
.A2(n_379),
.B(n_380),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3319),
.Y(n_3459)
);

AOI22xp5_ASAP7_75t_L g3460 ( 
.A1(n_3371),
.A2(n_382),
.B1(n_379),
.B2(n_381),
.Y(n_3460)
);

OR2x2_ASAP7_75t_L g3461 ( 
.A(n_3320),
.B(n_381),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3322),
.Y(n_3462)
);

AOI31xp33_ASAP7_75t_L g3463 ( 
.A1(n_3395),
.A2(n_384),
.A3(n_382),
.B(n_383),
.Y(n_3463)
);

OAI31xp33_ASAP7_75t_SL g3464 ( 
.A1(n_3441),
.A2(n_386),
.A3(n_384),
.B(n_385),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_3341),
.B(n_388),
.Y(n_3465)
);

OAI22xp33_ASAP7_75t_SL g3466 ( 
.A1(n_3362),
.A2(n_391),
.B1(n_389),
.B2(n_390),
.Y(n_3466)
);

OAI22xp5_ASAP7_75t_L g3467 ( 
.A1(n_3386),
.A2(n_392),
.B1(n_389),
.B2(n_391),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3339),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_3364),
.B(n_393),
.Y(n_3469)
);

NAND4xp25_ASAP7_75t_L g3470 ( 
.A(n_3401),
.B(n_776),
.C(n_395),
.D(n_393),
.Y(n_3470)
);

OAI22xp5_ASAP7_75t_L g3471 ( 
.A1(n_3391),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3341),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3334),
.Y(n_3473)
);

O2A1O1Ixp33_ASAP7_75t_L g3474 ( 
.A1(n_3354),
.A2(n_398),
.B(n_394),
.C(n_397),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3347),
.Y(n_3475)
);

O2A1O1Ixp33_ASAP7_75t_L g3476 ( 
.A1(n_3332),
.A2(n_3406),
.B(n_3387),
.C(n_3327),
.Y(n_3476)
);

INVxp67_ASAP7_75t_SL g3477 ( 
.A(n_3366),
.Y(n_3477)
);

INVx1_ASAP7_75t_SL g3478 ( 
.A(n_3436),
.Y(n_3478)
);

NOR2xp33_ASAP7_75t_L g3479 ( 
.A(n_3360),
.B(n_397),
.Y(n_3479)
);

OAI222xp33_ASAP7_75t_L g3480 ( 
.A1(n_3433),
.A2(n_400),
.B1(n_402),
.B2(n_398),
.C1(n_399),
.C2(n_401),
.Y(n_3480)
);

AOI221xp5_ASAP7_75t_L g3481 ( 
.A1(n_3427),
.A2(n_3389),
.B1(n_3410),
.B2(n_3385),
.C(n_3373),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3335),
.B(n_399),
.Y(n_3482)
);

AND2x2_ASAP7_75t_L g3483 ( 
.A(n_3348),
.B(n_401),
.Y(n_3483)
);

AO21x1_ASAP7_75t_L g3484 ( 
.A1(n_3352),
.A2(n_403),
.B(n_405),
.Y(n_3484)
);

AOI321xp33_ASAP7_75t_L g3485 ( 
.A1(n_3345),
.A2(n_407),
.A3(n_409),
.B1(n_403),
.B2(n_406),
.C(n_408),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3346),
.Y(n_3486)
);

AOI322xp5_ASAP7_75t_L g3487 ( 
.A1(n_3418),
.A2(n_406),
.A3(n_407),
.B1(n_409),
.B2(n_410),
.C1(n_411),
.C2(n_412),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3343),
.Y(n_3488)
);

AOI22xp5_ASAP7_75t_L g3489 ( 
.A1(n_3333),
.A2(n_413),
.B1(n_410),
.B2(n_412),
.Y(n_3489)
);

INVxp33_ASAP7_75t_L g3490 ( 
.A(n_3380),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3377),
.Y(n_3491)
);

OAI21xp33_ASAP7_75t_L g3492 ( 
.A1(n_3338),
.A2(n_414),
.B(n_415),
.Y(n_3492)
);

O2A1O1Ixp33_ASAP7_75t_L g3493 ( 
.A1(n_3365),
.A2(n_417),
.B(n_415),
.C(n_416),
.Y(n_3493)
);

INVxp67_ASAP7_75t_L g3494 ( 
.A(n_3372),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3405),
.Y(n_3495)
);

AOI22xp33_ASAP7_75t_L g3496 ( 
.A1(n_3342),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_3496)
);

AOI22xp5_ASAP7_75t_L g3497 ( 
.A1(n_3353),
.A2(n_423),
.B1(n_420),
.B2(n_422),
.Y(n_3497)
);

NAND2x1_ASAP7_75t_L g3498 ( 
.A(n_3377),
.B(n_422),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3405),
.Y(n_3499)
);

NOR2xp33_ASAP7_75t_L g3500 ( 
.A(n_3368),
.B(n_423),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3356),
.Y(n_3501)
);

AOI22xp5_ASAP7_75t_L g3502 ( 
.A1(n_3361),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3429),
.B(n_424),
.Y(n_3503)
);

AND2x2_ASAP7_75t_L g3504 ( 
.A(n_3394),
.B(n_426),
.Y(n_3504)
);

A2O1A1Ixp33_ASAP7_75t_L g3505 ( 
.A1(n_3423),
.A2(n_429),
.B(n_427),
.C(n_428),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3330),
.Y(n_3506)
);

OAI33xp33_ASAP7_75t_L g3507 ( 
.A1(n_3370),
.A2(n_429),
.A3(n_431),
.B1(n_427),
.B2(n_428),
.B3(n_430),
.Y(n_3507)
);

INVx2_ASAP7_75t_L g3508 ( 
.A(n_3397),
.Y(n_3508)
);

NAND3xp33_ASAP7_75t_L g3509 ( 
.A(n_3337),
.B(n_432),
.C(n_433),
.Y(n_3509)
);

AND2x2_ASAP7_75t_SL g3510 ( 
.A(n_3363),
.B(n_433),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3397),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3369),
.Y(n_3512)
);

O2A1O1Ixp5_ASAP7_75t_L g3513 ( 
.A1(n_3376),
.A2(n_437),
.B(n_434),
.C(n_435),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3403),
.B(n_3425),
.Y(n_3514)
);

NOR3xp33_ASAP7_75t_L g3515 ( 
.A(n_3344),
.B(n_437),
.C(n_438),
.Y(n_3515)
);

AOI221xp5_ASAP7_75t_L g3516 ( 
.A1(n_3379),
.A2(n_440),
.B1(n_438),
.B2(n_439),
.C(n_441),
.Y(n_3516)
);

OAI22xp5_ASAP7_75t_L g3517 ( 
.A1(n_3411),
.A2(n_3421),
.B1(n_3435),
.B2(n_3381),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_SL g3518 ( 
.A(n_3424),
.B(n_439),
.Y(n_3518)
);

OAI22xp5_ASAP7_75t_SL g3519 ( 
.A1(n_3419),
.A2(n_3393),
.B1(n_3383),
.B2(n_3349),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_SL g3520 ( 
.A(n_3438),
.B(n_3378),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3400),
.B(n_440),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3428),
.Y(n_3522)
);

AND2x2_ASAP7_75t_L g3523 ( 
.A(n_3350),
.B(n_441),
.Y(n_3523)
);

INVx1_ASAP7_75t_SL g3524 ( 
.A(n_3437),
.Y(n_3524)
);

NOR2xp33_ASAP7_75t_L g3525 ( 
.A(n_3407),
.B(n_442),
.Y(n_3525)
);

NOR3xp33_ASAP7_75t_L g3526 ( 
.A(n_3351),
.B(n_443),
.C(n_444),
.Y(n_3526)
);

OAI221xp5_ASAP7_75t_L g3527 ( 
.A1(n_3442),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.C(n_447),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3440),
.B(n_446),
.Y(n_3528)
);

AOI21xp33_ASAP7_75t_SL g3529 ( 
.A1(n_3413),
.A2(n_776),
.B(n_448),
.Y(n_3529)
);

INVx1_ASAP7_75t_SL g3530 ( 
.A(n_3359),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3408),
.B(n_449),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3384),
.Y(n_3532)
);

OR2x2_ASAP7_75t_L g3533 ( 
.A(n_3358),
.B(n_449),
.Y(n_3533)
);

NOR2x1_ASAP7_75t_L g3534 ( 
.A(n_3318),
.B(n_450),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3388),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_SL g3536 ( 
.A(n_3374),
.B(n_450),
.Y(n_3536)
);

OAI22xp5_ASAP7_75t_L g3537 ( 
.A1(n_3398),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3430),
.Y(n_3538)
);

OAI221xp5_ASAP7_75t_L g3539 ( 
.A1(n_3367),
.A2(n_454),
.B1(n_451),
.B2(n_453),
.C(n_455),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_3412),
.B(n_3431),
.Y(n_3540)
);

AND3x2_ASAP7_75t_L g3541 ( 
.A(n_3392),
.B(n_455),
.C(n_456),
.Y(n_3541)
);

AOI322xp5_ASAP7_75t_L g3542 ( 
.A1(n_3396),
.A2(n_774),
.A3(n_460),
.B1(n_461),
.B2(n_462),
.C1(n_463),
.C2(n_465),
.Y(n_3542)
);

AOI321xp33_ASAP7_75t_L g3543 ( 
.A1(n_3432),
.A2(n_459),
.A3(n_462),
.B1(n_463),
.B2(n_465),
.C(n_468),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3399),
.Y(n_3544)
);

BUFx2_ASAP7_75t_SL g3545 ( 
.A(n_3404),
.Y(n_3545)
);

AOI211xp5_ASAP7_75t_L g3546 ( 
.A1(n_3414),
.A2(n_769),
.B(n_469),
.C(n_459),
.Y(n_3546)
);

AOI22xp5_ASAP7_75t_L g3547 ( 
.A1(n_3434),
.A2(n_473),
.B1(n_468),
.B2(n_470),
.Y(n_3547)
);

OAI21xp5_ASAP7_75t_L g3548 ( 
.A1(n_3439),
.A2(n_470),
.B(n_473),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3409),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_3416),
.Y(n_3550)
);

OR2x2_ASAP7_75t_L g3551 ( 
.A(n_3417),
.B(n_474),
.Y(n_3551)
);

AND2x2_ASAP7_75t_L g3552 ( 
.A(n_3422),
.B(n_474),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3420),
.B(n_475),
.Y(n_3553)
);

NOR2xp67_ASAP7_75t_L g3554 ( 
.A(n_3415),
.B(n_765),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3426),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3326),
.Y(n_3556)
);

OAI22xp33_ASAP7_75t_L g3557 ( 
.A1(n_3386),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.Y(n_3557)
);

AOI21xp33_ASAP7_75t_SL g3558 ( 
.A1(n_3326),
.A2(n_477),
.B(n_479),
.Y(n_3558)
);

INVx1_ASAP7_75t_SL g3559 ( 
.A(n_3326),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3326),
.Y(n_3560)
);

OR2x2_ASAP7_75t_L g3561 ( 
.A(n_3336),
.B(n_479),
.Y(n_3561)
);

OAI22xp33_ASAP7_75t_L g3562 ( 
.A1(n_3386),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.Y(n_3562)
);

OR2x2_ASAP7_75t_L g3563 ( 
.A(n_3336),
.B(n_482),
.Y(n_3563)
);

OAI221xp5_ASAP7_75t_L g3564 ( 
.A1(n_3328),
.A2(n_485),
.B1(n_483),
.B2(n_484),
.C(n_486),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_SL g3565 ( 
.A(n_3326),
.B(n_485),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3326),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3326),
.Y(n_3567)
);

AOI221xp5_ASAP7_75t_L g3568 ( 
.A1(n_3382),
.A2(n_489),
.B1(n_486),
.B2(n_488),
.C(n_490),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3336),
.Y(n_3569)
);

OR2x2_ASAP7_75t_L g3570 ( 
.A(n_3336),
.B(n_489),
.Y(n_3570)
);

AND2x2_ASAP7_75t_L g3571 ( 
.A(n_3328),
.B(n_490),
.Y(n_3571)
);

OAI31xp33_ASAP7_75t_SL g3572 ( 
.A1(n_3355),
.A2(n_493),
.A3(n_491),
.B(n_492),
.Y(n_3572)
);

AND2x2_ASAP7_75t_L g3573 ( 
.A(n_3328),
.B(n_491),
.Y(n_3573)
);

INVx1_ASAP7_75t_SL g3574 ( 
.A(n_3326),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3326),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3326),
.Y(n_3576)
);

AOI221xp5_ASAP7_75t_L g3577 ( 
.A1(n_3382),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.C(n_496),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3328),
.B(n_494),
.Y(n_3578)
);

AOI21xp33_ASAP7_75t_L g3579 ( 
.A1(n_3326),
.A2(n_497),
.B(n_498),
.Y(n_3579)
);

AOI221xp5_ASAP7_75t_L g3580 ( 
.A1(n_3382),
.A2(n_500),
.B1(n_497),
.B2(n_499),
.C(n_503),
.Y(n_3580)
);

AOI22xp33_ASAP7_75t_SL g3581 ( 
.A1(n_3371),
.A2(n_504),
.B1(n_500),
.B2(n_503),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3328),
.B(n_504),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3326),
.Y(n_3583)
);

OR2x2_ASAP7_75t_L g3584 ( 
.A(n_3336),
.B(n_506),
.Y(n_3584)
);

NAND3xp33_ASAP7_75t_L g3585 ( 
.A(n_3326),
.B(n_507),
.C(n_508),
.Y(n_3585)
);

OAI322xp33_ASAP7_75t_L g3586 ( 
.A1(n_3326),
.A2(n_507),
.A3(n_508),
.B1(n_509),
.B2(n_510),
.C1(n_511),
.C2(n_512),
.Y(n_3586)
);

HB1xp67_ASAP7_75t_L g3587 ( 
.A(n_3326),
.Y(n_3587)
);

A2O1A1Ixp33_ASAP7_75t_L g3588 ( 
.A1(n_3357),
.A2(n_511),
.B(n_509),
.C(n_510),
.Y(n_3588)
);

A2O1A1Ixp33_ASAP7_75t_L g3589 ( 
.A1(n_3357),
.A2(n_515),
.B(n_513),
.C(n_514),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3326),
.Y(n_3590)
);

A2O1A1Ixp33_ASAP7_75t_L g3591 ( 
.A1(n_3357),
.A2(n_517),
.B(n_513),
.C(n_515),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3328),
.B(n_518),
.Y(n_3592)
);

OAI221xp5_ASAP7_75t_SL g3593 ( 
.A1(n_3410),
.A2(n_520),
.B1(n_518),
.B2(n_519),
.C(n_522),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3326),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3326),
.Y(n_3595)
);

AND2x2_ASAP7_75t_L g3596 ( 
.A(n_3328),
.B(n_519),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3326),
.Y(n_3597)
);

OAI21xp5_ASAP7_75t_L g3598 ( 
.A1(n_3328),
.A2(n_520),
.B(n_522),
.Y(n_3598)
);

NAND3xp33_ASAP7_75t_L g3599 ( 
.A(n_3326),
.B(n_523),
.C(n_524),
.Y(n_3599)
);

OAI22xp33_ASAP7_75t_L g3600 ( 
.A1(n_3386),
.A2(n_525),
.B1(n_523),
.B2(n_524),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3326),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3572),
.B(n_525),
.Y(n_3602)
);

NOR2xp33_ASAP7_75t_L g3603 ( 
.A(n_3472),
.B(n_526),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3498),
.Y(n_3604)
);

INVx2_ASAP7_75t_SL g3605 ( 
.A(n_3491),
.Y(n_3605)
);

NOR3x1_ASAP7_75t_L g3606 ( 
.A(n_3470),
.B(n_526),
.C(n_527),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3541),
.B(n_527),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_3477),
.A2(n_530),
.B(n_531),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3495),
.B(n_530),
.Y(n_3609)
);

O2A1O1Ixp33_ASAP7_75t_SL g3610 ( 
.A1(n_3499),
.A2(n_533),
.B(n_531),
.C(n_532),
.Y(n_3610)
);

OR2x2_ASAP7_75t_L g3611 ( 
.A(n_3478),
.B(n_3508),
.Y(n_3611)
);

NOR2xp33_ASAP7_75t_L g3612 ( 
.A(n_3511),
.B(n_535),
.Y(n_3612)
);

INVx2_ASAP7_75t_SL g3613 ( 
.A(n_3561),
.Y(n_3613)
);

NAND2xp33_ASAP7_75t_L g3614 ( 
.A(n_3587),
.B(n_3534),
.Y(n_3614)
);

AOI21xp5_ASAP7_75t_L g3615 ( 
.A1(n_3474),
.A2(n_3518),
.B(n_3450),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_L g3616 ( 
.A(n_3464),
.B(n_535),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3456),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3581),
.B(n_536),
.Y(n_3618)
);

AOI211xp5_ASAP7_75t_L g3619 ( 
.A1(n_3451),
.A2(n_539),
.B(n_536),
.C(n_538),
.Y(n_3619)
);

AOI21xp5_ASAP7_75t_L g3620 ( 
.A1(n_3481),
.A2(n_539),
.B(n_540),
.Y(n_3620)
);

NOR3x1_ASAP7_75t_L g3621 ( 
.A(n_3446),
.B(n_540),
.C(n_541),
.Y(n_3621)
);

INVx1_ASAP7_75t_SL g3622 ( 
.A(n_3510),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3563),
.Y(n_3623)
);

NOR2xp33_ASAP7_75t_L g3624 ( 
.A(n_3559),
.B(n_3574),
.Y(n_3624)
);

AOI22xp5_ASAP7_75t_SL g3625 ( 
.A1(n_3545),
.A2(n_764),
.B1(n_543),
.B2(n_541),
.Y(n_3625)
);

OAI21xp33_ASAP7_75t_L g3626 ( 
.A1(n_3555),
.A2(n_542),
.B(n_544),
.Y(n_3626)
);

NOR3xp33_ASAP7_75t_L g3627 ( 
.A(n_3447),
.B(n_542),
.C(n_545),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3570),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_SL g3629 ( 
.A(n_3489),
.B(n_3554),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3445),
.B(n_546),
.Y(n_3630)
);

AOI221xp5_ASAP7_75t_SL g3631 ( 
.A1(n_3476),
.A2(n_546),
.B1(n_547),
.B2(n_548),
.C(n_549),
.Y(n_3631)
);

OA22x2_ASAP7_75t_L g3632 ( 
.A1(n_3453),
.A2(n_551),
.B1(n_548),
.B2(n_550),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3569),
.B(n_551),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3584),
.Y(n_3634)
);

HB1xp67_ASAP7_75t_L g3635 ( 
.A(n_3554),
.Y(n_3635)
);

AOI22xp5_ASAP7_75t_L g3636 ( 
.A1(n_3452),
.A2(n_3448),
.B1(n_3519),
.B2(n_3571),
.Y(n_3636)
);

NOR2x1_ASAP7_75t_SL g3637 ( 
.A(n_3444),
.B(n_552),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3469),
.Y(n_3638)
);

NAND2xp33_ASAP7_75t_L g3639 ( 
.A(n_3515),
.B(n_552),
.Y(n_3639)
);

NOR3xp33_ASAP7_75t_SL g3640 ( 
.A(n_3593),
.B(n_553),
.C(n_554),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_3489),
.B(n_3455),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3558),
.B(n_555),
.Y(n_3642)
);

AOI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_3454),
.A2(n_555),
.B(n_556),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3465),
.Y(n_3644)
);

AOI221xp5_ASAP7_75t_L g3645 ( 
.A1(n_3517),
.A2(n_556),
.B1(n_557),
.B2(n_558),
.C(n_559),
.Y(n_3645)
);

NOR2xp33_ASAP7_75t_L g3646 ( 
.A(n_3463),
.B(n_557),
.Y(n_3646)
);

NOR2xp33_ASAP7_75t_L g3647 ( 
.A(n_3458),
.B(n_559),
.Y(n_3647)
);

AOI211xp5_ASAP7_75t_L g3648 ( 
.A1(n_3484),
.A2(n_562),
.B(n_560),
.C(n_561),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_3449),
.B(n_560),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_SL g3650 ( 
.A(n_3466),
.B(n_562),
.Y(n_3650)
);

NOR2xp33_ASAP7_75t_L g3651 ( 
.A(n_3482),
.B(n_563),
.Y(n_3651)
);

OAI221xp5_ASAP7_75t_L g3652 ( 
.A1(n_3516),
.A2(n_563),
.B1(n_564),
.B2(n_565),
.C(n_566),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3483),
.Y(n_3653)
);

O2A1O1Ixp33_ASAP7_75t_L g3654 ( 
.A1(n_3480),
.A2(n_566),
.B(n_564),
.C(n_565),
.Y(n_3654)
);

HB1xp67_ASAP7_75t_L g3655 ( 
.A(n_3459),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3461),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_SL g3657 ( 
.A(n_3485),
.B(n_567),
.Y(n_3657)
);

AOI22xp5_ASAP7_75t_L g3658 ( 
.A1(n_3573),
.A2(n_570),
.B1(n_567),
.B2(n_569),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3504),
.B(n_569),
.Y(n_3659)
);

NOR2xp33_ASAP7_75t_L g3660 ( 
.A(n_3492),
.B(n_570),
.Y(n_3660)
);

NOR2xp33_ASAP7_75t_L g3661 ( 
.A(n_3468),
.B(n_571),
.Y(n_3661)
);

INVx2_ASAP7_75t_L g3662 ( 
.A(n_3533),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_3551),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3596),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3487),
.B(n_572),
.Y(n_3665)
);

INVx2_ASAP7_75t_SL g3666 ( 
.A(n_3552),
.Y(n_3666)
);

OR2x2_ASAP7_75t_L g3667 ( 
.A(n_3578),
.B(n_572),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3460),
.B(n_573),
.Y(n_3668)
);

NOR3x1_ASAP7_75t_L g3669 ( 
.A(n_3548),
.B(n_573),
.C(n_574),
.Y(n_3669)
);

AOI21xp5_ASAP7_75t_L g3670 ( 
.A1(n_3565),
.A2(n_575),
.B(n_576),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3457),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3582),
.Y(n_3672)
);

NOR2x1_ASAP7_75t_L g3673 ( 
.A(n_3585),
.B(n_575),
.Y(n_3673)
);

NOR3x1_ASAP7_75t_L g3674 ( 
.A(n_3520),
.B(n_576),
.C(n_577),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3592),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3475),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3443),
.B(n_577),
.Y(n_3677)
);

OAI21xp33_ASAP7_75t_L g3678 ( 
.A1(n_3490),
.A2(n_578),
.B(n_579),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3523),
.Y(n_3679)
);

INVxp67_ASAP7_75t_L g3680 ( 
.A(n_3500),
.Y(n_3680)
);

NOR2xp67_ASAP7_75t_L g3681 ( 
.A(n_3599),
.B(n_3462),
.Y(n_3681)
);

AOI21xp33_ASAP7_75t_L g3682 ( 
.A1(n_3556),
.A2(n_764),
.B(n_581),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3560),
.B(n_582),
.Y(n_3683)
);

INVx1_ASAP7_75t_SL g3684 ( 
.A(n_3524),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3521),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3566),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3486),
.Y(n_3687)
);

NOR2xp33_ASAP7_75t_L g3688 ( 
.A(n_3501),
.B(n_582),
.Y(n_3688)
);

NOR2xp33_ASAP7_75t_L g3689 ( 
.A(n_3601),
.B(n_583),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3567),
.Y(n_3690)
);

OAI21xp5_ASAP7_75t_L g3691 ( 
.A1(n_3493),
.A2(n_584),
.B(n_585),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3575),
.B(n_584),
.Y(n_3692)
);

NAND3xp33_ASAP7_75t_L g3693 ( 
.A(n_3576),
.B(n_763),
.C(n_586),
.Y(n_3693)
);

NOR2xp33_ASAP7_75t_L g3694 ( 
.A(n_3583),
.B(n_586),
.Y(n_3694)
);

AOI211xp5_ASAP7_75t_L g3695 ( 
.A1(n_3557),
.A2(n_589),
.B(n_587),
.C(n_588),
.Y(n_3695)
);

AOI21xp5_ASAP7_75t_L g3696 ( 
.A1(n_3514),
.A2(n_587),
.B(n_589),
.Y(n_3696)
);

OAI21xp33_ASAP7_75t_L g3697 ( 
.A1(n_3540),
.A2(n_590),
.B(n_591),
.Y(n_3697)
);

AOI211xp5_ASAP7_75t_L g3698 ( 
.A1(n_3626),
.A2(n_3594),
.B(n_3595),
.C(n_3590),
.Y(n_3698)
);

NAND4xp75_ASAP7_75t_L g3699 ( 
.A(n_3674),
.B(n_3597),
.C(n_3473),
.D(n_3535),
.Y(n_3699)
);

AOI221xp5_ASAP7_75t_L g3700 ( 
.A1(n_3620),
.A2(n_3494),
.B1(n_3536),
.B2(n_3530),
.C(n_3529),
.Y(n_3700)
);

OAI222xp33_ASAP7_75t_L g3701 ( 
.A1(n_3622),
.A2(n_3544),
.B1(n_3549),
.B2(n_3532),
.C1(n_3550),
.C2(n_3488),
.Y(n_3701)
);

NOR2x1_ASAP7_75t_L g3702 ( 
.A(n_3604),
.B(n_3509),
.Y(n_3702)
);

OAI31xp33_ASAP7_75t_L g3703 ( 
.A1(n_3626),
.A2(n_3505),
.A3(n_3589),
.B(n_3588),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3637),
.Y(n_3704)
);

O2A1O1Ixp33_ASAP7_75t_L g3705 ( 
.A1(n_3657),
.A2(n_3513),
.B(n_3591),
.C(n_3503),
.Y(n_3705)
);

NOR3x1_ASAP7_75t_L g3706 ( 
.A(n_3652),
.B(n_3527),
.C(n_3598),
.Y(n_3706)
);

OAI21xp5_ASAP7_75t_SL g3707 ( 
.A1(n_3636),
.A2(n_3522),
.B(n_3506),
.Y(n_3707)
);

AOI221x1_ASAP7_75t_L g3708 ( 
.A1(n_3627),
.A2(n_3526),
.B1(n_3579),
.B2(n_3512),
.C(n_3538),
.Y(n_3708)
);

AOI221xp5_ASAP7_75t_L g3709 ( 
.A1(n_3615),
.A2(n_3580),
.B1(n_3577),
.B2(n_3568),
.C(n_3600),
.Y(n_3709)
);

AOI222xp33_ASAP7_75t_L g3710 ( 
.A1(n_3614),
.A2(n_3629),
.B1(n_3635),
.B2(n_3624),
.C1(n_3681),
.C2(n_3684),
.Y(n_3710)
);

NOR3xp33_ASAP7_75t_L g3711 ( 
.A(n_3617),
.B(n_3479),
.C(n_3553),
.Y(n_3711)
);

INVx2_ASAP7_75t_L g3712 ( 
.A(n_3611),
.Y(n_3712)
);

HB1xp67_ASAP7_75t_L g3713 ( 
.A(n_3655),
.Y(n_3713)
);

NAND4xp25_ASAP7_75t_SL g3714 ( 
.A(n_3631),
.B(n_3546),
.C(n_3547),
.D(n_3496),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3605),
.B(n_3638),
.Y(n_3715)
);

BUFx2_ASAP7_75t_L g3716 ( 
.A(n_3673),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3625),
.B(n_3562),
.Y(n_3717)
);

NOR3xp33_ASAP7_75t_SL g3718 ( 
.A(n_3641),
.B(n_3650),
.C(n_3691),
.Y(n_3718)
);

NAND2xp33_ASAP7_75t_SL g3719 ( 
.A(n_3640),
.B(n_3531),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3667),
.Y(n_3720)
);

AOI221xp5_ASAP7_75t_L g3721 ( 
.A1(n_3654),
.A2(n_3586),
.B1(n_3507),
.B2(n_3467),
.C(n_3471),
.Y(n_3721)
);

AOI221xp5_ASAP7_75t_L g3722 ( 
.A1(n_3619),
.A2(n_3537),
.B1(n_3525),
.B2(n_3564),
.C(n_3539),
.Y(n_3722)
);

OAI22xp33_ASAP7_75t_L g3723 ( 
.A1(n_3602),
.A2(n_3528),
.B1(n_3497),
.B2(n_3502),
.Y(n_3723)
);

NOR2xp33_ASAP7_75t_L g3724 ( 
.A(n_3697),
.B(n_3543),
.Y(n_3724)
);

AOI322xp5_ASAP7_75t_L g3725 ( 
.A1(n_3639),
.A2(n_3542),
.A3(n_591),
.B1(n_592),
.B2(n_594),
.C1(n_595),
.C2(n_596),
.Y(n_3725)
);

AOI211xp5_ASAP7_75t_L g3726 ( 
.A1(n_3676),
.A2(n_597),
.B(n_590),
.C(n_596),
.Y(n_3726)
);

A2O1A1Ixp33_ASAP7_75t_L g3727 ( 
.A1(n_3646),
.A2(n_762),
.B(n_600),
.C(n_598),
.Y(n_3727)
);

OAI21xp5_ASAP7_75t_L g3728 ( 
.A1(n_3616),
.A2(n_598),
.B(n_599),
.Y(n_3728)
);

NOR3xp33_ASAP7_75t_L g3729 ( 
.A(n_3649),
.B(n_599),
.C(n_600),
.Y(n_3729)
);

O2A1O1Ixp33_ASAP7_75t_L g3730 ( 
.A1(n_3610),
.A2(n_601),
.B(n_602),
.C(n_603),
.Y(n_3730)
);

OAI21xp5_ASAP7_75t_L g3731 ( 
.A1(n_3696),
.A2(n_602),
.B(n_603),
.Y(n_3731)
);

NAND3xp33_ASAP7_75t_L g3732 ( 
.A(n_3648),
.B(n_604),
.C(n_605),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3666),
.B(n_604),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3607),
.Y(n_3734)
);

OAI21xp5_ASAP7_75t_L g3735 ( 
.A1(n_3665),
.A2(n_605),
.B(n_606),
.Y(n_3735)
);

NAND5xp2_ASAP7_75t_L g3736 ( 
.A(n_3664),
.B(n_608),
.C(n_609),
.D(n_610),
.E(n_611),
.Y(n_3736)
);

NOR3xp33_ASAP7_75t_L g3737 ( 
.A(n_3680),
.B(n_3613),
.C(n_3628),
.Y(n_3737)
);

AOI21xp33_ASAP7_75t_SL g3738 ( 
.A1(n_3632),
.A2(n_610),
.B(n_611),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3679),
.Y(n_3739)
);

AOI22xp5_ASAP7_75t_L g3740 ( 
.A1(n_3647),
.A2(n_612),
.B1(n_613),
.B2(n_614),
.Y(n_3740)
);

NAND2x1_ASAP7_75t_L g3741 ( 
.A(n_3623),
.B(n_612),
.Y(n_3741)
);

OAI21xp5_ASAP7_75t_SL g3742 ( 
.A1(n_3634),
.A2(n_613),
.B(n_615),
.Y(n_3742)
);

AOI221xp5_ASAP7_75t_L g3743 ( 
.A1(n_3609),
.A2(n_616),
.B1(n_617),
.B2(n_618),
.C(n_619),
.Y(n_3743)
);

OAI21xp5_ASAP7_75t_SL g3744 ( 
.A1(n_3687),
.A2(n_617),
.B(n_618),
.Y(n_3744)
);

AOI22xp5_ASAP7_75t_L g3745 ( 
.A1(n_3651),
.A2(n_619),
.B1(n_620),
.B2(n_621),
.Y(n_3745)
);

INVx2_ASAP7_75t_SL g3746 ( 
.A(n_3656),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3612),
.B(n_620),
.Y(n_3747)
);

AOI221xp5_ASAP7_75t_L g3748 ( 
.A1(n_3686),
.A2(n_621),
.B1(n_622),
.B2(n_623),
.C(n_624),
.Y(n_3748)
);

NAND4xp25_ASAP7_75t_L g3749 ( 
.A(n_3606),
.B(n_624),
.C(n_625),
.D(n_626),
.Y(n_3749)
);

OR2x2_ASAP7_75t_L g3750 ( 
.A(n_3630),
.B(n_625),
.Y(n_3750)
);

XNOR2xp5_ASAP7_75t_L g3751 ( 
.A(n_3695),
.B(n_626),
.Y(n_3751)
);

NOR2xp33_ASAP7_75t_L g3752 ( 
.A(n_3697),
.B(n_627),
.Y(n_3752)
);

AOI211xp5_ASAP7_75t_SL g3753 ( 
.A1(n_3690),
.A2(n_627),
.B(n_628),
.C(n_629),
.Y(n_3753)
);

AOI21xp33_ASAP7_75t_L g3754 ( 
.A1(n_3653),
.A2(n_628),
.B(n_630),
.Y(n_3754)
);

AOI22xp33_ASAP7_75t_SL g3755 ( 
.A1(n_3663),
.A2(n_630),
.B1(n_631),
.B2(n_632),
.Y(n_3755)
);

AOI22xp33_ASAP7_75t_L g3756 ( 
.A1(n_3672),
.A2(n_631),
.B1(n_632),
.B2(n_633),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3662),
.Y(n_3757)
);

AOI21xp5_ASAP7_75t_L g3758 ( 
.A1(n_3643),
.A2(n_633),
.B(n_634),
.Y(n_3758)
);

NAND3xp33_ASAP7_75t_L g3759 ( 
.A(n_3608),
.B(n_3694),
.C(n_3689),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3704),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3713),
.Y(n_3761)
);

AOI22xp5_ASAP7_75t_L g3762 ( 
.A1(n_3724),
.A2(n_3660),
.B1(n_3675),
.B2(n_3685),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3741),
.Y(n_3763)
);

INVxp67_ASAP7_75t_SL g3764 ( 
.A(n_3730),
.Y(n_3764)
);

NOR2xp33_ASAP7_75t_L g3765 ( 
.A(n_3749),
.B(n_3678),
.Y(n_3765)
);

AOI31xp33_ASAP7_75t_L g3766 ( 
.A1(n_3698),
.A2(n_3633),
.A3(n_3618),
.B(n_3644),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3715),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3712),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3746),
.Y(n_3769)
);

AO22x2_ASAP7_75t_L g3770 ( 
.A1(n_3699),
.A2(n_3677),
.B1(n_3692),
.B2(n_3683),
.Y(n_3770)
);

OAI22xp5_ASAP7_75t_L g3771 ( 
.A1(n_3732),
.A2(n_3740),
.B1(n_3717),
.B2(n_3757),
.Y(n_3771)
);

INVxp67_ASAP7_75t_SL g3772 ( 
.A(n_3702),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3751),
.Y(n_3773)
);

AOI221xp5_ASAP7_75t_L g3774 ( 
.A1(n_3701),
.A2(n_3671),
.B1(n_3682),
.B2(n_3645),
.C(n_3670),
.Y(n_3774)
);

AND4x1_ASAP7_75t_L g3775 ( 
.A(n_3710),
.B(n_3718),
.C(n_3621),
.D(n_3753),
.Y(n_3775)
);

INVx2_ASAP7_75t_SL g3776 ( 
.A(n_3716),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3733),
.Y(n_3777)
);

AOI22xp5_ASAP7_75t_L g3778 ( 
.A1(n_3719),
.A2(n_3603),
.B1(n_3688),
.B2(n_3661),
.Y(n_3778)
);

OAI22xp5_ASAP7_75t_L g3779 ( 
.A1(n_3739),
.A2(n_3693),
.B1(n_3642),
.B2(n_3659),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3747),
.Y(n_3780)
);

AOI22xp5_ASAP7_75t_L g3781 ( 
.A1(n_3737),
.A2(n_3668),
.B1(n_3658),
.B2(n_3669),
.Y(n_3781)
);

BUFx2_ASAP7_75t_L g3782 ( 
.A(n_3731),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3752),
.Y(n_3783)
);

OAI22x1_ASAP7_75t_L g3784 ( 
.A1(n_3714),
.A2(n_634),
.B1(n_635),
.B2(n_636),
.Y(n_3784)
);

INVxp67_ASAP7_75t_L g3785 ( 
.A(n_3736),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3750),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3734),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3745),
.Y(n_3788)
);

AOI22xp5_ASAP7_75t_L g3789 ( 
.A1(n_3711),
.A2(n_637),
.B1(n_638),
.B2(n_639),
.Y(n_3789)
);

AOI221xp5_ASAP7_75t_L g3790 ( 
.A1(n_3738),
.A2(n_637),
.B1(n_638),
.B2(n_639),
.C(n_640),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3727),
.Y(n_3791)
);

AOI22xp5_ASAP7_75t_L g3792 ( 
.A1(n_3721),
.A2(n_640),
.B1(n_641),
.B2(n_642),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3720),
.Y(n_3793)
);

AOI22xp5_ASAP7_75t_L g3794 ( 
.A1(n_3709),
.A2(n_642),
.B1(n_643),
.B2(n_644),
.Y(n_3794)
);

AOI221xp5_ASAP7_75t_L g3795 ( 
.A1(n_3723),
.A2(n_644),
.B1(n_645),
.B2(n_646),
.C(n_647),
.Y(n_3795)
);

OAI22x1_ASAP7_75t_L g3796 ( 
.A1(n_3759),
.A2(n_645),
.B1(n_646),
.B2(n_648),
.Y(n_3796)
);

AND2x2_ASAP7_75t_L g3797 ( 
.A(n_3760),
.B(n_3728),
.Y(n_3797)
);

NAND5xp2_ASAP7_75t_L g3798 ( 
.A(n_3774),
.B(n_3707),
.C(n_3700),
.D(n_3705),
.E(n_3781),
.Y(n_3798)
);

AOI211xp5_ASAP7_75t_L g3799 ( 
.A1(n_3771),
.A2(n_3735),
.B(n_3722),
.C(n_3744),
.Y(n_3799)
);

AOI221xp5_ASAP7_75t_SL g3800 ( 
.A1(n_3766),
.A2(n_3758),
.B1(n_3743),
.B2(n_3748),
.C(n_3726),
.Y(n_3800)
);

AOI21xp33_ASAP7_75t_SL g3801 ( 
.A1(n_3763),
.A2(n_3729),
.B(n_3754),
.Y(n_3801)
);

AOI31xp33_ASAP7_75t_L g3802 ( 
.A1(n_3772),
.A2(n_3755),
.A3(n_3756),
.B(n_3725),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3764),
.B(n_3725),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3767),
.Y(n_3804)
);

HB1xp67_ASAP7_75t_L g3805 ( 
.A(n_3784),
.Y(n_3805)
);

NOR2xp33_ASAP7_75t_L g3806 ( 
.A(n_3785),
.B(n_3742),
.Y(n_3806)
);

AOI221xp5_ASAP7_75t_L g3807 ( 
.A1(n_3761),
.A2(n_3703),
.B1(n_3706),
.B2(n_3708),
.C(n_652),
.Y(n_3807)
);

OAI211xp5_ASAP7_75t_L g3808 ( 
.A1(n_3792),
.A2(n_3778),
.B(n_3762),
.C(n_3790),
.Y(n_3808)
);

NOR3xp33_ASAP7_75t_L g3809 ( 
.A(n_3779),
.B(n_649),
.C(n_650),
.Y(n_3809)
);

AOI221xp5_ASAP7_75t_L g3810 ( 
.A1(n_3776),
.A2(n_651),
.B1(n_653),
.B2(n_654),
.C(n_655),
.Y(n_3810)
);

NOR2xp67_ASAP7_75t_SL g3811 ( 
.A(n_3768),
.B(n_3769),
.Y(n_3811)
);

OAI22xp33_ASAP7_75t_L g3812 ( 
.A1(n_3794),
.A2(n_651),
.B1(n_653),
.B2(n_654),
.Y(n_3812)
);

XNOR2xp5_ASAP7_75t_L g3813 ( 
.A(n_3775),
.B(n_762),
.Y(n_3813)
);

AOI22xp5_ASAP7_75t_L g3814 ( 
.A1(n_3765),
.A2(n_655),
.B1(n_656),
.B2(n_657),
.Y(n_3814)
);

AOI221xp5_ASAP7_75t_L g3815 ( 
.A1(n_3770),
.A2(n_658),
.B1(n_659),
.B2(n_660),
.C(n_661),
.Y(n_3815)
);

AOI321xp33_ASAP7_75t_L g3816 ( 
.A1(n_3799),
.A2(n_3791),
.A3(n_3793),
.B1(n_3787),
.B2(n_3773),
.C(n_3788),
.Y(n_3816)
);

OAI222xp33_ASAP7_75t_L g3817 ( 
.A1(n_3811),
.A2(n_3782),
.B1(n_3783),
.B2(n_3786),
.C1(n_3777),
.C2(n_3780),
.Y(n_3817)
);

OAI211xp5_ASAP7_75t_SL g3818 ( 
.A1(n_3807),
.A2(n_3795),
.B(n_3789),
.C(n_3770),
.Y(n_3818)
);

OAI31xp33_ASAP7_75t_L g3819 ( 
.A1(n_3808),
.A2(n_3796),
.A3(n_659),
.B(n_660),
.Y(n_3819)
);

OAI221xp5_ASAP7_75t_L g3820 ( 
.A1(n_3815),
.A2(n_658),
.B1(n_662),
.B2(n_663),
.C(n_664),
.Y(n_3820)
);

AOI221xp5_ASAP7_75t_L g3821 ( 
.A1(n_3802),
.A2(n_662),
.B1(n_663),
.B2(n_665),
.C(n_666),
.Y(n_3821)
);

OAI211xp5_ASAP7_75t_SL g3822 ( 
.A1(n_3803),
.A2(n_668),
.B(n_669),
.C(n_670),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_SL g3823 ( 
.A(n_3812),
.B(n_670),
.Y(n_3823)
);

AOI221xp5_ASAP7_75t_L g3824 ( 
.A1(n_3801),
.A2(n_3798),
.B1(n_3806),
.B2(n_3804),
.C(n_3805),
.Y(n_3824)
);

OAI211xp5_ASAP7_75t_SL g3825 ( 
.A1(n_3809),
.A2(n_761),
.B(n_673),
.C(n_674),
.Y(n_3825)
);

O2A1O1Ixp33_ASAP7_75t_L g3826 ( 
.A1(n_3797),
.A2(n_671),
.B(n_673),
.C(n_675),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3813),
.Y(n_3827)
);

OAI211xp5_ASAP7_75t_L g3828 ( 
.A1(n_3800),
.A2(n_3810),
.B(n_3814),
.C(n_677),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3827),
.Y(n_3829)
);

AND2x2_ASAP7_75t_L g3830 ( 
.A(n_3824),
.B(n_675),
.Y(n_3830)
);

AOI221x1_ASAP7_75t_SL g3831 ( 
.A1(n_3816),
.A2(n_676),
.B1(n_677),
.B2(n_678),
.C(n_679),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3821),
.B(n_676),
.Y(n_3832)
);

AOI222xp33_ASAP7_75t_L g3833 ( 
.A1(n_3817),
.A2(n_678),
.B1(n_679),
.B2(n_680),
.C1(n_683),
.C2(n_684),
.Y(n_3833)
);

NAND3xp33_ASAP7_75t_L g3834 ( 
.A(n_3819),
.B(n_3822),
.C(n_3820),
.Y(n_3834)
);

INVx2_ASAP7_75t_SL g3835 ( 
.A(n_3823),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3826),
.Y(n_3836)
);

OAI22xp5_ASAP7_75t_L g3837 ( 
.A1(n_3828),
.A2(n_683),
.B1(n_684),
.B2(n_685),
.Y(n_3837)
);

A2O1A1Ixp33_ASAP7_75t_L g3838 ( 
.A1(n_3825),
.A2(n_685),
.B(n_686),
.C(n_688),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3833),
.B(n_3818),
.Y(n_3839)
);

AND2x4_ASAP7_75t_L g3840 ( 
.A(n_3829),
.B(n_3835),
.Y(n_3840)
);

NOR4xp75_ASAP7_75t_L g3841 ( 
.A(n_3837),
.B(n_689),
.C(n_690),
.D(n_693),
.Y(n_3841)
);

NAND4xp75_ASAP7_75t_L g3842 ( 
.A(n_3830),
.B(n_690),
.C(n_694),
.D(n_695),
.Y(n_3842)
);

BUFx4f_ASAP7_75t_SL g3843 ( 
.A(n_3840),
.Y(n_3843)
);

NOR3xp33_ASAP7_75t_L g3844 ( 
.A(n_3839),
.B(n_3836),
.C(n_3832),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3842),
.Y(n_3845)
);

OR2x2_ASAP7_75t_L g3846 ( 
.A(n_3845),
.B(n_3838),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3846),
.Y(n_3847)
);

AOI22xp5_ASAP7_75t_L g3848 ( 
.A1(n_3847),
.A2(n_3843),
.B1(n_3834),
.B2(n_3844),
.Y(n_3848)
);

AOI22xp5_ASAP7_75t_L g3849 ( 
.A1(n_3848),
.A2(n_3831),
.B1(n_3841),
.B2(n_698),
.Y(n_3849)
);

AOI31xp33_ASAP7_75t_L g3850 ( 
.A1(n_3849),
.A2(n_695),
.A3(n_697),
.B(n_698),
.Y(n_3850)
);

AOI22xp5_ASAP7_75t_L g3851 ( 
.A1(n_3850),
.A2(n_699),
.B1(n_700),
.B2(n_701),
.Y(n_3851)
);

AOI22xp33_ASAP7_75t_L g3852 ( 
.A1(n_3851),
.A2(n_699),
.B1(n_700),
.B2(n_702),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3852),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3853),
.Y(n_3854)
);

OR2x2_ASAP7_75t_L g3855 ( 
.A(n_3854),
.B(n_702),
.Y(n_3855)
);

AOI221xp5_ASAP7_75t_L g3856 ( 
.A1(n_3855),
.A2(n_703),
.B1(n_704),
.B2(n_705),
.C(n_707),
.Y(n_3856)
);

AOI211xp5_ASAP7_75t_L g3857 ( 
.A1(n_3856),
.A2(n_704),
.B(n_708),
.C(n_709),
.Y(n_3857)
);


endmodule