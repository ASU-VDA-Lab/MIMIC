module fake_jpeg_7721_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_39),
.Y(n_56)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_40),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_24),
.A2(n_1),
.B(n_2),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_1),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_24),
.B1(n_21),
.B2(n_30),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_54),
.B1(n_55),
.B2(n_23),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_24),
.B1(n_28),
.B2(n_19),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_37),
.B1(n_32),
.B2(n_39),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_56),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_19),
.B1(n_21),
.B2(n_26),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_29),
.B1(n_17),
.B2(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_65),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_37),
.B1(n_19),
.B2(n_32),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_75),
.B1(n_76),
.B2(n_52),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_44),
.B1(n_42),
.B2(n_47),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_32),
.B1(n_39),
.B2(n_34),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_74),
.B1(n_44),
.B2(n_52),
.Y(n_87)
);

CKINVDCx9p33_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_69),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_40),
.B(n_16),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_68),
.Y(n_83)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_18),
.B1(n_52),
.B2(n_46),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

CKINVDCx9p33_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_34),
.B1(n_39),
.B2(n_15),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_15),
.B1(n_29),
.B2(n_23),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_79),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_87),
.B1(n_90),
.B2(n_75),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_25),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_33),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_89),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_77),
.B(n_70),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_46),
.B1(n_33),
.B2(n_36),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_72),
.B1(n_67),
.B2(n_22),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_100),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_SL g98 ( 
.A(n_64),
.B(n_49),
.C(n_33),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_16),
.B(n_49),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_13),
.C(n_12),
.Y(n_100)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_3),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_71),
.B(n_40),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_111),
.B1(n_128),
.B2(n_130),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_68),
.C(n_78),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_119),
.C(n_88),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_102),
.B(n_63),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_12),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_120),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_36),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_73),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_122),
.B(n_94),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_40),
.B(n_71),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_84),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_75),
.B1(n_46),
.B2(n_22),
.Y(n_128)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_3),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_129),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_85),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_140),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_143),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_127),
.A2(n_108),
.B1(n_124),
.B2(n_115),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_137),
.A2(n_150),
.B1(n_36),
.B2(n_20),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_83),
.Y(n_141)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_86),
.B(n_101),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_145),
.B(n_146),
.Y(n_159)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_97),
.C(n_101),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_149),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_106),
.B(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_106),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_84),
.B1(n_72),
.B2(n_94),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_49),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_16),
.B(n_20),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_153),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_158),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_111),
.B(n_129),
.C(n_114),
.D(n_109),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_171),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_65),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_164),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_162),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_13),
.C(n_6),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_103),
.B1(n_91),
.B2(n_22),
.Y(n_163)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_150),
.B1(n_148),
.B2(n_136),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_133),
.B1(n_139),
.B2(n_137),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_140),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_136),
.C(n_169),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_172),
.B(n_151),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_185),
.Y(n_188)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_187),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_132),
.C(n_144),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_160),
.C(n_159),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_133),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_172),
.B(n_152),
.Y(n_185)
);

INVxp33_ASAP7_75t_SL g186 ( 
.A(n_168),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_SL g189 ( 
.A(n_186),
.B(n_142),
.C(n_159),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_192),
.B(n_190),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_194),
.C(n_195),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_174),
.A2(n_186),
.B(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_156),
.C(n_164),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_170),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_171),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_20),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_176),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_207),
.C(n_205),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_65),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_178),
.C(n_167),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_188),
.C(n_65),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_5),
.B(n_6),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_157),
.B(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_210),
.C(n_212),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_188),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_211),
.B(n_202),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_5),
.B(n_6),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_217),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_213),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_201),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_221),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_222),
.A3(n_201),
.B1(n_212),
.B2(n_203),
.C1(n_10),
.C2(n_5),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

OAI311xp33_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_224),
.A3(n_8),
.B1(n_9),
.C1(n_10),
.Y(n_227)
);

OAI221xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_11),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_11),
.Y(n_229)
);


endmodule