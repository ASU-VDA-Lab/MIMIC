module fake_jpeg_735_n_193 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_193);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_15),
.B(n_22),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_0),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx6f_ASAP7_75t_SL g82 ( 
.A(n_73),
.Y(n_82)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_88),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_75),
.A2(n_61),
.B1(n_48),
.B2(n_52),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_52),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_51),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_65),
.B1(n_66),
.B2(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_48),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_47),
.B(n_56),
.C(n_51),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_90),
.B(n_105),
.Y(n_126)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_46),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_98),
.Y(n_114)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_55),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_103),
.Y(n_122)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_67),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_26),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_83),
.B(n_87),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_108),
.A2(n_9),
.B(n_11),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_111),
.B(n_118),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_87),
.B1(n_59),
.B2(n_58),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_115),
.B1(n_117),
.B2(n_96),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_87),
.B1(n_59),
.B2(n_4),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_2),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_21),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_123),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_23),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_106),
.B1(n_104),
.B2(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_27),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_6),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_127),
.B(n_11),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_101),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_132),
.Y(n_166)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_91),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_135),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_137),
.B1(n_12),
.B2(n_13),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_140),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_122),
.B1(n_119),
.B2(n_120),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_12),
.B(n_14),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_29),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_28),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_144),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_122),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_149),
.Y(n_164)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_122),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_142),
.B1(n_143),
.B2(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_158),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_35),
.C(n_43),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_156),
.C(n_135),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_31),
.C(n_42),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_18),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_164),
.B(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_170),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_172),
.B1(n_150),
.B2(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_156),
.C(n_155),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_175),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

FAx1_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_153),
.CI(n_154),
.CON(n_178),
.SN(n_178)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_180),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_163),
.C(n_153),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_165),
.C(n_36),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_181),
.B(n_39),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_184),
.B(n_41),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_182),
.B(n_178),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_188),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_183),
.B(n_186),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_190),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_177),
.C(n_169),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_45),
.Y(n_193)
);


endmodule