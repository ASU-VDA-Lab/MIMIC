module fake_aes_3071_n_670 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_670);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_670;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx14_ASAP7_75t_R g77 ( .A(n_40), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_57), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_54), .Y(n_79) );
INVxp67_ASAP7_75t_L g80 ( .A(n_24), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_47), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_75), .Y(n_82) );
INVxp33_ASAP7_75t_SL g83 ( .A(n_36), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_67), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_76), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_22), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_8), .Y(n_87) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_70), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_9), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_69), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_15), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_66), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_15), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_64), .Y(n_95) );
NOR2xp33_ASAP7_75t_L g96 ( .A(n_73), .B(n_18), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_25), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_51), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_39), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_34), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_37), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_48), .Y(n_102) );
BUFx10_ASAP7_75t_L g103 ( .A(n_63), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_6), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_7), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_3), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_10), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_3), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_14), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_26), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_45), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_35), .B(n_28), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_21), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_65), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_50), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_41), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_52), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_9), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_14), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_7), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_19), .Y(n_122) );
BUFx2_ASAP7_75t_SL g123 ( .A(n_32), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_31), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_106), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_101), .Y(n_126) );
NOR2xp33_ASAP7_75t_R g127 ( .A(n_77), .B(n_29), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_101), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_78), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_106), .Y(n_130) );
NAND2x1_ASAP7_75t_L g131 ( .A(n_87), .B(n_0), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_82), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_112), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_78), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_112), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_84), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_115), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_86), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_122), .Y(n_140) );
INVx2_ASAP7_75t_SL g141 ( .A(n_103), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_122), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_105), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_120), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_88), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_103), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_81), .B(n_0), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_90), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_92), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_90), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_91), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_107), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_103), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_105), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_103), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_91), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_114), .B(n_1), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_114), .B(n_1), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_82), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_119), .B(n_2), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_93), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_104), .B(n_4), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_93), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_97), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_87), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_89), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_82), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_145), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_145), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_157), .A2(n_110), .B1(n_89), .B2(n_108), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_141), .B(n_121), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
INVx2_ASAP7_75t_SL g173 ( .A(n_141), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_149), .B(n_121), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_132), .Y(n_175) );
AO22x2_ASAP7_75t_L g176 ( .A1(n_131), .A2(n_124), .B1(n_117), .B2(n_97), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_157), .A2(n_94), .B1(n_108), .B2(n_109), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_145), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_146), .B(n_80), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_137), .Y(n_181) );
BUFx2_ASAP7_75t_L g182 ( .A(n_144), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_157), .B(n_119), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_159), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_145), .Y(n_186) );
OAI221xp5_ASAP7_75t_L g187 ( .A1(n_129), .A2(n_109), .B1(n_110), .B2(n_85), .C(n_100), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_159), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_160), .Y(n_189) );
OR2x2_ASAP7_75t_L g190 ( .A(n_142), .B(n_123), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_147), .B(n_123), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_153), .B(n_79), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_167), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_147), .B(n_124), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_155), .B(n_83), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_126), .B(n_95), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_138), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_160), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_167), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_160), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_129), .B(n_98), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_143), .Y(n_202) );
AND2x6_ASAP7_75t_L g203 ( .A(n_160), .B(n_118), .Y(n_203) );
INVx4_ASAP7_75t_L g204 ( .A(n_158), .Y(n_204) );
OR2x6_ASAP7_75t_L g205 ( .A(n_131), .B(n_118), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_143), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_143), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_134), .B(n_117), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_134), .Y(n_209) );
BUFx2_ASAP7_75t_L g210 ( .A(n_128), .Y(n_210) );
AO22x2_ASAP7_75t_L g211 ( .A1(n_136), .A2(n_111), .B1(n_102), .B2(n_99), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_136), .B(n_111), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_139), .B(n_102), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_154), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_139), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_148), .B(n_99), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_148), .B(n_116), .Y(n_217) );
OR2x2_ASAP7_75t_L g218 ( .A(n_133), .B(n_4), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_150), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_150), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_151), .B(n_116), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_151), .B(n_95), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_156), .B(n_88), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_135), .B(n_88), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_154), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_154), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_156), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_152), .Y(n_228) );
BUFx3_ASAP7_75t_L g229 ( .A(n_161), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_228), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_193), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_204), .B(n_161), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_219), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_204), .B(n_164), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_172), .Y(n_236) );
BUFx12f_ASAP7_75t_L g237 ( .A(n_182), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_204), .B(n_164), .Y(n_238) );
NOR2x1_ASAP7_75t_L g239 ( .A(n_205), .B(n_162), .Y(n_239) );
NAND2xp33_ASAP7_75t_SL g240 ( .A(n_204), .B(n_127), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_219), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_179), .B(n_130), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_194), .B(n_163), .Y(n_243) );
INVx3_ASAP7_75t_SL g244 ( .A(n_181), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_219), .B(n_158), .Y(n_245) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_220), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_220), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_220), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_182), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_194), .B(n_163), .Y(n_250) );
NOR2xp33_ASAP7_75t_R g251 ( .A(n_197), .B(n_140), .Y(n_251) );
INVx2_ASAP7_75t_SL g252 ( .A(n_229), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_229), .B(n_166), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_229), .B(n_165), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_172), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_175), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_203), .A2(n_96), .B1(n_88), .B2(n_113), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_209), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_198), .Y(n_259) );
BUFx4f_ASAP7_75t_SL g260 ( .A(n_210), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_175), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_209), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_203), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_191), .B(n_5), .Y(n_264) );
INVxp67_ASAP7_75t_SL g265 ( .A(n_189), .Y(n_265) );
NOR3xp33_ASAP7_75t_SL g266 ( .A(n_187), .B(n_125), .C(n_6), .Y(n_266) );
BUFx2_ASAP7_75t_L g267 ( .A(n_203), .Y(n_267) );
NOR3xp33_ASAP7_75t_SL g268 ( .A(n_196), .B(n_5), .C(n_8), .Y(n_268) );
AOI21x1_ASAP7_75t_L g269 ( .A1(n_223), .A2(n_88), .B(n_43), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_215), .Y(n_270) );
NOR3xp33_ASAP7_75t_L g271 ( .A(n_218), .B(n_10), .C(n_11), .Y(n_271) );
OR2x6_ASAP7_75t_L g272 ( .A(n_205), .B(n_176), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_191), .B(n_11), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_201), .B(n_88), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_185), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_198), .B(n_12), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_215), .Y(n_277) );
NOR3xp33_ASAP7_75t_SL g278 ( .A(n_192), .B(n_12), .C(n_13), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_227), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_185), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_205), .B(n_13), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_188), .Y(n_282) );
NOR2xp33_ASAP7_75t_R g283 ( .A(n_210), .B(n_46), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_188), .Y(n_284) );
INVxp67_ASAP7_75t_SL g285 ( .A(n_189), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_205), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_218), .B(n_16), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_227), .A2(n_16), .B(n_17), .C(n_18), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_174), .Y(n_289) );
OR2x6_ASAP7_75t_L g290 ( .A(n_205), .B(n_17), .Y(n_290) );
INVx4_ASAP7_75t_L g291 ( .A(n_203), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_203), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_199), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_199), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_208), .B(n_19), .Y(n_295) );
OR2x6_ASAP7_75t_L g296 ( .A(n_290), .B(n_198), .Y(n_296) );
INVxp67_ASAP7_75t_L g297 ( .A(n_249), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_234), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_253), .B(n_174), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_258), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_291), .B(n_173), .Y(n_301) );
NAND2xp33_ASAP7_75t_L g302 ( .A(n_286), .B(n_203), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_254), .B(n_190), .Y(n_303) );
BUFx4f_ASAP7_75t_L g304 ( .A(n_290), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_289), .B(n_190), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_243), .B(n_203), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_291), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_258), .A2(n_200), .B(n_180), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_237), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_262), .A2(n_200), .B(n_180), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_242), .B(n_195), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_281), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_281), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_250), .B(n_177), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_262), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_244), .B(n_177), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_270), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_270), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_264), .B(n_273), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_291), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_264), .B(n_208), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_264), .B(n_208), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_291), .B(n_173), .Y(n_323) );
AOI21x1_ASAP7_75t_L g324 ( .A1(n_269), .A2(n_211), .B(n_216), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_277), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_234), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_286), .A2(n_198), .B1(n_189), .B2(n_180), .Y(n_327) );
NAND2xp33_ASAP7_75t_L g328 ( .A(n_292), .B(n_211), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_260), .B(n_171), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_264), .A2(n_171), .B1(n_211), .B2(n_180), .Y(n_330) );
BUFx12f_ASAP7_75t_L g331 ( .A(n_237), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_277), .Y(n_332) );
O2A1O1Ixp5_ASAP7_75t_L g333 ( .A1(n_240), .A2(n_224), .B(n_183), .C(n_171), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_279), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_234), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_281), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_259), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_239), .B(n_171), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_273), .B(n_213), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_279), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_281), .B(n_212), .Y(n_341) );
INVx6_ASAP7_75t_L g342 ( .A(n_234), .Y(n_342) );
OAI21xp33_ASAP7_75t_SL g343 ( .A1(n_290), .A2(n_212), .B(n_213), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_231), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_234), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_236), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_318), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_320), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_300), .Y(n_349) );
AOI21xp33_ASAP7_75t_L g350 ( .A1(n_311), .A2(n_287), .B(n_239), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_304), .A2(n_290), .B1(n_272), .B2(n_276), .Y(n_351) );
BUFx12f_ASAP7_75t_L g352 ( .A(n_331), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_318), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_297), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_300), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_315), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_339), .B(n_287), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_304), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_339), .B(n_233), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_314), .A2(n_266), .B1(n_271), .B2(n_230), .C(n_251), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_304), .A2(n_272), .B1(n_290), .B2(n_259), .Y(n_361) );
AOI21xp33_ASAP7_75t_L g362 ( .A1(n_343), .A2(n_272), .B(n_295), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_320), .Y(n_363) );
INVx4_ASAP7_75t_L g364 ( .A(n_296), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_316), .B(n_244), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_330), .A2(n_272), .B1(n_276), .B2(n_211), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_341), .B(n_272), .Y(n_367) );
NAND2xp33_ASAP7_75t_SL g368 ( .A(n_312), .B(n_263), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_319), .A2(n_276), .B1(n_208), .B2(n_216), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_339), .B(n_235), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_325), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_325), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_305), .B(n_244), .Y(n_373) );
NAND3xp33_ASAP7_75t_SL g374 ( .A(n_309), .B(n_230), .C(n_283), .Y(n_374) );
OAI221xp5_ASAP7_75t_L g375 ( .A1(n_303), .A2(n_170), .B1(n_238), .B2(n_268), .C(n_278), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_316), .A2(n_259), .B1(n_263), .B2(n_267), .Y(n_376) );
BUFx6f_ASAP7_75t_SL g377 ( .A(n_296), .Y(n_377) );
AOI21xp33_ASAP7_75t_L g378 ( .A1(n_343), .A2(n_274), .B(n_257), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_366), .A2(n_296), .B1(n_312), .B2(n_336), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_360), .A2(n_299), .B1(n_329), .B2(n_305), .C(n_303), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_349), .B(n_341), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_347), .B(n_332), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_350), .A2(n_299), .B1(n_338), .B2(n_176), .C(n_183), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_349), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_369), .A2(n_328), .B(n_296), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_355), .Y(n_387) );
AOI211xp5_ASAP7_75t_L g388 ( .A1(n_351), .A2(n_328), .B(n_288), .C(n_302), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_355), .B(n_336), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_347), .B(n_332), .Y(n_390) );
OAI33xp33_ASAP7_75t_L g391 ( .A1(n_373), .A2(n_221), .A3(n_327), .B1(n_321), .B2(n_322), .B3(n_206), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_356), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_356), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_365), .A2(n_176), .B1(n_313), .B2(n_302), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_366), .A2(n_313), .B1(n_176), .B2(n_340), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_375), .A2(n_331), .B1(n_183), .B2(n_340), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_351), .A2(n_309), .B1(n_317), .B2(n_315), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_356), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_377), .A2(n_183), .B1(n_334), .B2(n_317), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g401 ( .A1(n_378), .A2(n_308), .B(n_310), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_353), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_357), .B(n_346), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_353), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_377), .A2(n_334), .B1(n_301), .B2(n_323), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_371), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_402), .B(n_406), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_404), .B(n_371), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_381), .B(n_372), .Y(n_409) );
OAI221xp5_ASAP7_75t_L g410 ( .A1(n_380), .A2(n_397), .B1(n_373), .B2(n_396), .C(n_395), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_402), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_381), .B(n_372), .Y(n_412) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_396), .A2(n_369), .B1(n_364), .B2(n_358), .Y(n_413) );
AOI31xp33_ASAP7_75t_L g414 ( .A1(n_386), .A2(n_361), .A3(n_362), .B(n_377), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_391), .A2(n_354), .B1(n_374), .B2(n_370), .C(n_359), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_379), .A2(n_377), .B1(n_367), .B2(n_362), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_398), .A2(n_367), .B1(n_364), .B2(n_358), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_406), .B(n_346), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_384), .A2(n_378), .B1(n_245), .B2(n_217), .C(n_222), .Y(n_419) );
OA21x2_ASAP7_75t_L g420 ( .A1(n_401), .A2(n_324), .B(n_269), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_403), .A2(n_364), .B1(n_358), .B2(n_352), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_385), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_404), .B(n_402), .Y(n_423) );
NAND3xp33_ASAP7_75t_L g424 ( .A(n_388), .B(n_333), .C(n_364), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_385), .Y(n_425) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_385), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_400), .A2(n_376), .B1(n_368), .B2(n_306), .C(n_202), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_406), .A2(n_217), .B1(n_222), .B2(n_216), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_383), .B(n_348), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_405), .A2(n_217), .B1(n_222), .B2(n_216), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_388), .A2(n_275), .B1(n_236), .B2(n_294), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_383), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_389), .A2(n_217), .B1(n_222), .B2(n_352), .Y(n_434) );
NOR4xp25_ASAP7_75t_SL g435 ( .A(n_387), .B(n_267), .C(n_352), .D(n_324), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g436 ( .A(n_401), .B(n_348), .C(n_363), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_387), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_392), .Y(n_438) );
AOI221x1_ASAP7_75t_L g439 ( .A1(n_392), .A2(n_348), .B1(n_345), .B2(n_344), .C(n_301), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_382), .A2(n_225), .B1(n_206), .B2(n_207), .C(n_226), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_382), .A2(n_202), .B1(n_226), .B2(n_207), .C(n_214), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_407), .B(n_393), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_437), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_410), .B(n_390), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_407), .B(n_393), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_407), .B(n_394), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_422), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_407), .B(n_399), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_433), .Y(n_449) );
AOI211xp5_ASAP7_75t_L g450 ( .A1(n_421), .A2(n_214), .B(n_390), .C(n_225), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_433), .Y(n_451) );
INVx4_ASAP7_75t_L g452 ( .A(n_430), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_418), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_409), .B(n_399), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_438), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_438), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_415), .B(n_225), .C(n_399), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_418), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_411), .Y(n_459) );
INVx4_ASAP7_75t_L g460 ( .A(n_430), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_422), .B(n_389), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_434), .A2(n_414), .B1(n_424), .B2(n_413), .C(n_409), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_430), .B(n_348), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_430), .Y(n_464) );
OAI321xp33_ASAP7_75t_L g465 ( .A1(n_424), .A2(n_225), .A3(n_261), .B1(n_255), .B2(n_256), .C(n_294), .Y(n_465) );
OAI21xp33_ASAP7_75t_L g466 ( .A1(n_414), .A2(n_225), .B(n_169), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_412), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_422), .B(n_363), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_416), .A2(n_301), .B1(n_323), .B2(n_337), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_423), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_417), .A2(n_363), .B1(n_344), .B2(n_323), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_425), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_412), .B(n_20), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_425), .B(n_280), .Y(n_474) );
AOI33xp33_ASAP7_75t_L g475 ( .A1(n_431), .A2(n_20), .A3(n_21), .B1(n_293), .B2(n_284), .B3(n_282), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_428), .B(n_261), .Y(n_476) );
AOI221xp5_ASAP7_75t_SL g477 ( .A1(n_408), .A2(n_225), .B1(n_255), .B2(n_293), .C(n_256), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_428), .B(n_284), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_428), .B(n_282), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_426), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_408), .B(n_275), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_419), .A2(n_337), .B1(n_265), .B2(n_285), .Y(n_482) );
BUFx2_ASAP7_75t_L g483 ( .A(n_432), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_420), .B(n_232), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_436), .B(n_231), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_432), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_429), .B(n_337), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_427), .B(n_232), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_436), .Y(n_489) );
INVx5_ASAP7_75t_L g490 ( .A(n_480), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_445), .B(n_420), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_449), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_445), .B(n_420), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_458), .B(n_420), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_452), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_451), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_459), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_467), .B(n_439), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_443), .B(n_441), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_444), .B(n_439), .Y(n_500) );
NOR2xp33_ASAP7_75t_R g501 ( .A(n_483), .B(n_298), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_446), .B(n_435), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_453), .B(n_298), .Y(n_503) );
NOR2xp33_ASAP7_75t_R g504 ( .A(n_473), .B(n_326), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_470), .B(n_435), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_454), .B(n_335), .Y(n_506) );
NAND2xp33_ASAP7_75t_R g507 ( .A(n_442), .B(n_23), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g508 ( .A1(n_444), .A2(n_440), .B1(n_342), .B2(n_335), .C(n_326), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_446), .B(n_27), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_455), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_472), .B(n_30), .Y(n_511) );
NOR2xp33_ASAP7_75t_R g512 ( .A(n_452), .B(n_345), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_456), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_442), .B(n_33), .Y(n_514) );
INVx4_ASAP7_75t_L g515 ( .A(n_442), .Y(n_515) );
NAND2xp33_ASAP7_75t_SL g516 ( .A(n_452), .B(n_460), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_461), .B(n_345), .Y(n_517) );
INVx5_ASAP7_75t_L g518 ( .A(n_480), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_448), .B(n_38), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_448), .B(n_42), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_461), .B(n_44), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_448), .B(n_49), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_468), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_464), .B(n_53), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_447), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_476), .B(n_342), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_460), .B(n_55), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_447), .B(n_56), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_484), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_460), .B(n_58), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_476), .B(n_342), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_489), .B(n_59), .Y(n_532) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_450), .B(n_186), .C(n_178), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_484), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_478), .B(n_342), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_468), .Y(n_536) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_466), .A2(n_184), .B(n_168), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_478), .B(n_60), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_462), .A2(n_241), .B1(n_247), .B2(n_307), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g540 ( .A(n_475), .B(n_184), .C(n_169), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_479), .B(n_61), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_474), .Y(n_542) );
OAI31xp67_ASAP7_75t_L g543 ( .A1(n_475), .A2(n_168), .A3(n_68), .B(n_71), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_497), .Y(n_544) );
NAND2x1_ASAP7_75t_L g545 ( .A(n_515), .B(n_463), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_507), .A2(n_486), .B1(n_463), .B2(n_457), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g547 ( .A(n_500), .B(n_477), .C(n_488), .Y(n_547) );
INVx2_ASAP7_75t_SL g548 ( .A(n_512), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_492), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_512), .Y(n_550) );
INVxp67_ASAP7_75t_SL g551 ( .A(n_507), .Y(n_551) );
OAI32xp33_ASAP7_75t_L g552 ( .A1(n_516), .A2(n_474), .A3(n_471), .B1(n_481), .B2(n_485), .Y(n_552) );
NAND3xp33_ASAP7_75t_SL g553 ( .A(n_504), .B(n_469), .C(n_482), .Y(n_553) );
NAND4xp25_ASAP7_75t_L g554 ( .A(n_500), .B(n_463), .C(n_487), .D(n_485), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_496), .B(n_479), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_490), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_539), .A2(n_465), .B1(n_186), .B2(n_178), .C(n_247), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_490), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_510), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_504), .A2(n_307), .B1(n_241), .B2(n_320), .Y(n_560) );
AOI21xp33_ASAP7_75t_SL g561 ( .A1(n_533), .A2(n_62), .B(n_72), .Y(n_561) );
AOI21xp33_ASAP7_75t_SL g562 ( .A1(n_543), .A2(n_292), .B(n_307), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_513), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_505), .B(n_178), .C(n_186), .Y(n_564) );
OAI322xp33_ASAP7_75t_L g565 ( .A1(n_499), .A2(n_178), .A3(n_186), .B1(n_246), .B2(n_248), .C1(n_252), .C2(n_320), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_515), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_515), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_523), .B(n_178), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_490), .A2(n_320), .B1(n_248), .B2(n_252), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_536), .B(n_178), .Y(n_570) );
OAI21xp33_ASAP7_75t_L g571 ( .A1(n_498), .A2(n_186), .B(n_501), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_542), .B(n_186), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_516), .A2(n_490), .B(n_518), .Y(n_573) );
INVx3_ASAP7_75t_L g574 ( .A(n_518), .Y(n_574) );
NAND2x1_ASAP7_75t_SL g575 ( .A(n_495), .B(n_527), .Y(n_575) );
NAND2xp33_ASAP7_75t_SL g576 ( .A(n_501), .B(n_495), .Y(n_576) );
INVxp67_ASAP7_75t_L g577 ( .A(n_514), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_518), .A2(n_521), .B1(n_530), .B2(n_495), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_514), .B(n_503), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_491), .B(n_493), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_511), .Y(n_581) );
XOR2x2_ASAP7_75t_L g582 ( .A(n_524), .B(n_520), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_518), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_525), .Y(n_584) );
INVx3_ASAP7_75t_L g585 ( .A(n_518), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_491), .B(n_493), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_524), .B(n_532), .C(n_502), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_529), .Y(n_588) );
NAND2x1p5_ASAP7_75t_L g589 ( .A(n_511), .B(n_522), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_538), .A2(n_541), .B(n_522), .Y(n_590) );
AOI222xp33_ASAP7_75t_L g591 ( .A1(n_494), .A2(n_502), .B1(n_509), .B2(n_520), .C1(n_519), .C2(n_534), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_580), .B(n_534), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_583), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_549), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_586), .B(n_509), .Y(n_595) );
BUFx2_ASAP7_75t_L g596 ( .A(n_576), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_544), .B(n_517), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_586), .B(n_532), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_574), .Y(n_599) );
O2A1O1Ixp5_ASAP7_75t_SL g600 ( .A1(n_561), .A2(n_535), .B(n_526), .C(n_531), .Y(n_600) );
INVx2_ASAP7_75t_SL g601 ( .A(n_574), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_550), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_559), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_563), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_588), .B(n_519), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_584), .Y(n_606) );
XNOR2xp5_ASAP7_75t_L g607 ( .A(n_582), .B(n_538), .Y(n_607) );
INVxp67_ASAP7_75t_SL g608 ( .A(n_585), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_555), .Y(n_609) );
NOR3xp33_ASAP7_75t_L g610 ( .A(n_547), .B(n_508), .C(n_540), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_555), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_591), .B(n_541), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_585), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_572), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_572), .Y(n_615) );
NOR4xp25_ASAP7_75t_SL g616 ( .A(n_551), .B(n_537), .C(n_506), .D(n_528), .Y(n_616) );
NOR2x1_ASAP7_75t_L g617 ( .A(n_573), .B(n_537), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_556), .Y(n_618) );
AOI21xp33_ASAP7_75t_L g619 ( .A1(n_552), .A2(n_591), .B(n_587), .Y(n_619) );
NOR3xp33_ASAP7_75t_SL g620 ( .A(n_553), .B(n_554), .C(n_571), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_566), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_558), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_581), .B(n_567), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_577), .B(n_566), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_603), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_603), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_604), .Y(n_627) );
AO22x1_ASAP7_75t_L g628 ( .A1(n_596), .A2(n_590), .B1(n_548), .B2(n_578), .Y(n_628) );
INVx2_ASAP7_75t_SL g629 ( .A(n_602), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_593), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_607), .A2(n_589), .B1(n_590), .B2(n_546), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_596), .A2(n_545), .B(n_578), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_619), .A2(n_564), .B(n_565), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_604), .Y(n_634) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_612), .A2(n_589), .B1(n_579), .B2(n_570), .Y(n_635) );
NOR2xp67_ASAP7_75t_SL g636 ( .A(n_599), .B(n_575), .Y(n_636) );
AOI32xp33_ASAP7_75t_L g637 ( .A1(n_612), .A2(n_560), .A3(n_557), .B1(n_569), .B2(n_568), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_623), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_610), .A2(n_557), .B1(n_569), .B2(n_562), .Y(n_639) );
AOI31xp33_ASAP7_75t_L g640 ( .A1(n_607), .A2(n_608), .A3(n_601), .B(n_617), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_609), .B(n_611), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_630), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_641), .Y(n_643) );
AOI211xp5_ASAP7_75t_L g644 ( .A1(n_631), .A2(n_624), .B(n_601), .C(n_599), .Y(n_644) );
NAND4xp25_ASAP7_75t_SL g645 ( .A(n_632), .B(n_595), .C(n_600), .D(n_598), .Y(n_645) );
AOI211xp5_ASAP7_75t_L g646 ( .A1(n_631), .A2(n_597), .B(n_621), .C(n_613), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_629), .Y(n_647) );
AOI31xp33_ASAP7_75t_L g648 ( .A1(n_633), .A2(n_620), .A3(n_595), .B(n_621), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_640), .A2(n_594), .B1(n_606), .B2(n_622), .C(n_618), .Y(n_649) );
NAND2xp33_ASAP7_75t_R g650 ( .A(n_633), .B(n_616), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_641), .Y(n_651) );
AND4x1_ASAP7_75t_L g652 ( .A(n_639), .B(n_622), .C(n_618), .D(n_592), .Y(n_652) );
AOI211xp5_ASAP7_75t_L g653 ( .A1(n_628), .A2(n_613), .B(n_614), .C(n_615), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_635), .A2(n_605), .B1(n_614), .B2(n_615), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_638), .A2(n_600), .B1(n_605), .B2(n_637), .C(n_626), .Y(n_655) );
NAND4xp75_ASAP7_75t_L g656 ( .A(n_625), .B(n_627), .C(n_634), .D(n_636), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_631), .A2(n_612), .B1(n_639), .B2(n_635), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_631), .A2(n_619), .B1(n_610), .B2(n_612), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_647), .Y(n_659) );
AND2x4_ASAP7_75t_L g660 ( .A(n_642), .B(n_657), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_656), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_658), .A2(n_645), .B1(n_655), .B2(n_649), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_659), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_661), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_662), .A2(n_648), .B1(n_644), .B2(n_646), .Y(n_665) );
OAI221xp5_ASAP7_75t_L g666 ( .A1(n_665), .A2(n_650), .B1(n_653), .B2(n_652), .C(n_654), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_663), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_667), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_664), .B1(n_660), .B2(n_666), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_669), .A2(n_660), .B1(n_650), .B2(n_651), .C(n_643), .Y(n_670) );
endmodule