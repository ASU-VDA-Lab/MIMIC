module fake_jpeg_2784_n_94 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_94);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_94;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_24),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_34),
.B1(n_28),
.B2(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_42),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_22),
.Y(n_42)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_27),
.B1(n_38),
.B2(n_35),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_1),
.C(n_2),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_28),
.B1(n_36),
.B2(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_40),
.B1(n_31),
.B2(n_4),
.Y(n_58)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_59),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_44),
.B(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_2),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_64),
.B1(n_53),
.B2(n_67),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_45),
.B(n_5),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_7),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_3),
.B(n_6),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_9),
.C(n_10),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_64)
);

AOI22x1_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_55),
.B1(n_52),
.B2(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_73),
.Y(n_81)
);

AO21x1_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_79),
.B(n_15),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_75),
.B(n_76),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_78),
.C(n_9),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_63),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_85),
.B1(n_79),
.B2(n_78),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_88),
.A2(n_87),
.B1(n_82),
.B2(n_84),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_89),
.A2(n_87),
.B1(n_80),
.B2(n_81),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_83),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_13),
.C(n_14),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_14),
.Y(n_94)
);


endmodule