module fake_jpeg_25614_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_73),
.Y(n_79)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_75),
.Y(n_81)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_48),
.B1(n_63),
.B2(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_78),
.B1(n_80),
.B2(n_49),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_67),
.B1(n_65),
.B2(n_58),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_87),
.B1(n_86),
.B2(n_59),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_62),
.B1(n_56),
.B2(n_51),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_67),
.B1(n_65),
.B2(n_44),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_50),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_45),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_87),
.Y(n_107)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_86),
.Y(n_110)
);

AOI211xp5_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_50),
.B(n_72),
.C(n_58),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_98),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_103),
.B(n_108),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_54),
.C(n_52),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_0),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_112),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_46),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_57),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_110),
.A2(n_102),
.B1(n_55),
.B2(n_53),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_117),
.B1(n_3),
.B2(n_4),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_118),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_104),
.A2(n_16),
.B1(n_40),
.B2(n_37),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_14),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_119),
.B(n_122),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_106),
.B1(n_4),
.B2(n_5),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_109),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_132),
.B1(n_134),
.B2(n_10),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_129),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_3),
.B(n_5),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_131),
.B(n_9),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_21),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_130),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_121),
.B(n_8),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_135),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_139),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_128),
.C(n_127),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_133),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_140),
.B1(n_141),
.B2(n_125),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_145),
.A2(n_142),
.B(n_138),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_136),
.C(n_123),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_132),
.B1(n_18),
.B2(n_20),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_28),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_149),
.B(n_22),
.C(n_23),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_26),
.Y(n_152)
);


endmodule