module fake_jpeg_24894_n_61 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_61);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_55;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_24;
wire n_26;
wire n_36;
wire n_31;
wire n_56;
wire n_25;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_7),
.B(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_15),
.B(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

OR2x2_ASAP7_75t_SL g38 ( 
.A(n_37),
.B(n_1),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_47)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_34),
.B1(n_23),
.B2(n_36),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_41),
.B1(n_45),
.B2(n_29),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_23),
.A2(n_29),
.B1(n_28),
.B2(n_37),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_40),
.B1(n_42),
.B2(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_46),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_49),
.B(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_27),
.B(n_48),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_18),
.C(n_24),
.Y(n_58)
);

AOI322xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.A3(n_24),
.B1(n_25),
.B2(n_30),
.C1(n_35),
.C2(n_44),
.Y(n_59)
);

FAx1_ASAP7_75t_SL g60 ( 
.A(n_59),
.B(n_26),
.CI(n_48),
.CON(n_60),
.SN(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_58),
.Y(n_61)
);


endmodule