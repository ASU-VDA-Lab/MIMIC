module fake_jpeg_27722_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_47),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_10),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

HAxp5_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_0),
.CON(n_70),
.SN(n_70)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_53),
.B1(n_66),
.B2(n_56),
.Y(n_78)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_75),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_78),
.Y(n_94)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_51),
.B1(n_65),
.B2(n_52),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_88),
.B1(n_55),
.B2(n_49),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_71),
.B1(n_57),
.B2(n_50),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_68),
.B1(n_64),
.B2(n_60),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_57),
.B1(n_69),
.B2(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_1),
.Y(n_107)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_54),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_103),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_69),
.B(n_50),
.C(n_64),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_99),
.B(n_18),
.C(n_40),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_62),
.B(n_26),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

BUFx2_ASAP7_75t_SL g114 ( 
.A(n_101),
.Y(n_114)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

CKINVDCx6p67_ASAP7_75t_R g113 ( 
.A(n_102),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_116)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_108),
.Y(n_112)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_110),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_68),
.C(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_17),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_105),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_21),
.B1(n_43),
.B2(n_42),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_97),
.B(n_106),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_127),
.Y(n_142)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_128),
.B(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_98),
.B(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_93),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_140)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_102),
.A3(n_113),
.B1(n_28),
.B2(n_32),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_141),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_100),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_146),
.C(n_11),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_10),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_143),
.B1(n_12),
.B2(n_13),
.Y(n_153)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_16),
.B(n_39),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_144),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_128),
.B(n_9),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_152),
.B(n_153),
.Y(n_159)
);

XNOR2x2_ASAP7_75t_SL g148 ( 
.A(n_142),
.B(n_11),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_151),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_145),
.A2(n_36),
.B1(n_14),
.B2(n_15),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_158),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.C(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_137),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_154),
.C(n_159),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_163),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_157),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_136),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_155),
.B(n_141),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_155),
.C(n_146),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_148),
.B(n_22),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_38),
.B(n_30),
.C(n_35),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_44),
.Y(n_172)
);


endmodule