module fake_ariane_794_n_1498 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1498);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1498;

wire n_913;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_334;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_552;
wire n_348;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_699;
wire n_590;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_887;
wire n_729;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1440;
wire n_1370;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_363;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_838;
wire n_383;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_208;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_140),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_66),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_88),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_157),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_177),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_51),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_107),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_51),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_33),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_47),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_24),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_45),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_191),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_27),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_63),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_2),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_101),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_110),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_85),
.Y(n_227)
);

INVx4_ASAP7_75t_R g228 ( 
.A(n_200),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_45),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_20),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_151),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_69),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_172),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_39),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_76),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_52),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_31),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_113),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_28),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_115),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_193),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_1),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_137),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_131),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_73),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_112),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_31),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_135),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_198),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_52),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_27),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_83),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_48),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_7),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_167),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_43),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_78),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_75),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_146),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_3),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_196),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_4),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_111),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_43),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_32),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_0),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_120),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_182),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_149),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_118),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_190),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_11),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_18),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_68),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_116),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_123),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_117),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_24),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_37),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_53),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_15),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_21),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_188),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_13),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_12),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_80),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_22),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_178),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_39),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_175),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_10),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_2),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_4),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_154),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_136),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_32),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_59),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_187),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_95),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_162),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_55),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_30),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_59),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_203),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_189),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_186),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_127),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_179),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_93),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_150),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_62),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_20),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_14),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_57),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_129),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_164),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_97),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_84),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_62),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_161),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_37),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_148),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_74),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_184),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_119),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_159),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_147),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_54),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_183),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_143),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_96),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_91),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_34),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_7),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_102),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_55),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_64),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_176),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_90),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_126),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_11),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_160),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_257),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_296),
.B(n_0),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_240),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_209),
.B(n_1),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_240),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_219),
.B(n_3),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_294),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_210),
.B(n_220),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_257),
.Y(n_356)
);

NOR2x1_ASAP7_75t_L g357 ( 
.A(n_221),
.B(n_77),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_289),
.Y(n_358)
);

BUFx8_ASAP7_75t_SL g359 ( 
.A(n_205),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_5),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_342),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_222),
.B(n_5),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_257),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_233),
.B(n_6),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_212),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_236),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_238),
.B(n_6),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_244),
.B(n_8),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_209),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_324),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_8),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_211),
.B(n_9),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_211),
.B(n_9),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_230),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_230),
.Y(n_376)
);

AND2x6_ASAP7_75t_L g377 ( 
.A(n_227),
.B(n_79),
.Y(n_377)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_240),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_212),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_240),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_286),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_213),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_240),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_213),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_286),
.B(n_10),
.Y(n_385)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_225),
.Y(n_386)
);

BUFx12f_ASAP7_75t_L g387 ( 
.A(n_320),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_246),
.B(n_12),
.Y(n_388)
);

INVx6_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_320),
.Y(n_390)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_249),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_343),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_227),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_251),
.B(n_13),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_323),
.B(n_14),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_225),
.B(n_15),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_332),
.B(n_16),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_343),
.Y(n_399)
);

BUFx12f_ASAP7_75t_L g400 ( 
.A(n_231),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_253),
.B(n_16),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_215),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_215),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_214),
.Y(n_404)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_263),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_268),
.B(n_17),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_272),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_204),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_224),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_275),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_280),
.B(n_17),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_257),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_241),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_288),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_204),
.Y(n_416)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_257),
.Y(n_417)
);

INVx5_ASAP7_75t_L g418 ( 
.A(n_257),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_329),
.B(n_18),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_334),
.B(n_19),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_217),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_257),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_247),
.B(n_19),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_242),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_257),
.B(n_21),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_273),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_217),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_252),
.B(n_22),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_285),
.B(n_23),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_274),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_273),
.B(n_23),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_255),
.B(n_25),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_243),
.Y(n_433)
);

BUFx8_ASAP7_75t_L g434 ( 
.A(n_228),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_391),
.B(n_218),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_396),
.A2(n_239),
.B1(n_297),
.B2(n_237),
.Y(n_436)
);

OR2x6_ASAP7_75t_L g437 ( 
.A(n_387),
.B(n_256),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_430),
.A2(n_341),
.B1(n_338),
.B2(n_218),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_391),
.B(n_279),
.Y(n_439)
);

OAI22xp33_ASAP7_75t_R g440 ( 
.A1(n_360),
.A2(n_346),
.B1(n_308),
.B2(n_258),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_396),
.A2(n_347),
.B1(n_310),
.B2(n_322),
.Y(n_441)
);

OAI22xp33_ASAP7_75t_R g442 ( 
.A1(n_429),
.A2(n_339),
.B1(n_265),
.B2(n_277),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_358),
.B(n_278),
.Y(n_444)
);

OAI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_353),
.A2(n_298),
.B1(n_279),
.B2(n_338),
.Y(n_445)
);

OAI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_355),
.A2(n_292),
.B1(n_229),
.B2(n_232),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_372),
.A2(n_307),
.B1(n_306),
.B2(n_235),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_390),
.A2(n_370),
.B1(n_402),
.B2(n_382),
.Y(n_448)
);

OAI22xp33_ASAP7_75t_SL g449 ( 
.A1(n_397),
.A2(n_284),
.B1(n_301),
.B2(n_259),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_391),
.B(n_321),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_351),
.A2(n_261),
.B1(n_267),
.B2(n_269),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_390),
.A2(n_318),
.B1(n_270),
.B2(n_271),
.Y(n_452)
);

OAI22xp33_ASAP7_75t_SL g453 ( 
.A1(n_397),
.A2(n_398),
.B1(n_362),
.B2(n_368),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_406),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_361),
.B(n_283),
.Y(n_455)
);

OAI22xp33_ASAP7_75t_SL g456 ( 
.A1(n_397),
.A2(n_302),
.B1(n_319),
.B2(n_287),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_424),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_406),
.Y(n_458)
);

BUFx10_ASAP7_75t_L g459 ( 
.A(n_389),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_366),
.B(n_206),
.Y(n_460)
);

OAI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_397),
.A2(n_326),
.B1(n_317),
.B2(n_316),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_351),
.A2(n_374),
.B1(n_385),
.B2(n_354),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_391),
.B(n_290),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_393),
.B(n_399),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_371),
.B(n_234),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_394),
.Y(n_467)
);

AO22x2_ASAP7_75t_L g468 ( 
.A1(n_371),
.A2(n_276),
.B1(n_295),
.B2(n_28),
.Y(n_468)
);

AOI22x1_ASAP7_75t_L g469 ( 
.A1(n_398),
.A2(n_345),
.B1(n_344),
.B2(n_340),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_389),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_389),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_393),
.B(n_206),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_370),
.A2(n_345),
.B1(n_344),
.B2(n_340),
.Y(n_473)
);

OAI22xp33_ASAP7_75t_L g474 ( 
.A1(n_393),
.A2(n_207),
.B1(n_336),
.B2(n_335),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_382),
.A2(n_337),
.B1(n_336),
.B2(n_335),
.Y(n_475)
);

OAI22xp33_ASAP7_75t_SL g476 ( 
.A1(n_398),
.A2(n_337),
.B1(n_331),
.B2(n_330),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_406),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_350),
.Y(n_478)
);

OAI22xp33_ASAP7_75t_L g479 ( 
.A1(n_393),
.A2(n_331),
.B1(n_330),
.B2(n_328),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_399),
.B(n_207),
.Y(n_480)
);

OAI22xp33_ASAP7_75t_L g481 ( 
.A1(n_399),
.A2(n_208),
.B1(n_216),
.B2(n_223),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_394),
.Y(n_482)
);

OAI22xp33_ASAP7_75t_R g483 ( 
.A1(n_365),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_399),
.B(n_208),
.Y(n_484)
);

AO22x2_ASAP7_75t_L g485 ( 
.A1(n_398),
.A2(n_349),
.B1(n_374),
.B2(n_351),
.Y(n_485)
);

OAI22xp33_ASAP7_75t_SL g486 ( 
.A1(n_367),
.A2(n_401),
.B1(n_412),
.B2(n_407),
.Y(n_486)
);

OAI22xp33_ASAP7_75t_L g487 ( 
.A1(n_402),
.A2(n_216),
.B1(n_223),
.B2(n_226),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_403),
.A2(n_328),
.B1(n_281),
.B2(n_226),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_403),
.A2(n_281),
.B1(n_325),
.B2(n_315),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_389),
.B(n_245),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_406),
.Y(n_491)
);

AO22x2_ASAP7_75t_L g492 ( 
.A1(n_349),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_406),
.Y(n_493)
);

AO22x2_ASAP7_75t_L g494 ( 
.A1(n_351),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_421),
.A2(n_327),
.B1(n_314),
.B2(n_313),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_408),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_387),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_408),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_394),
.Y(n_500)
);

OAI22xp33_ASAP7_75t_SL g501 ( 
.A1(n_419),
.A2(n_312),
.B1(n_311),
.B2(n_309),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_SL g502 ( 
.A(n_373),
.B(n_248),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_408),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_421),
.B(n_387),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_493),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_R g506 ( 
.A(n_504),
.B(n_423),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_443),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_498),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_454),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_493),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_458),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_436),
.B(n_441),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_465),
.B(n_423),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_477),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_438),
.B(n_359),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_491),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_460),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_478),
.Y(n_518)
);

BUFx6f_ASAP7_75t_SL g519 ( 
.A(n_437),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_495),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_497),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_414),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_499),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_503),
.Y(n_524)
);

INVxp33_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_464),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_467),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_482),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_500),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_437),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_485),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_462),
.B(n_414),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_478),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_478),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_438),
.B(n_468),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_462),
.B(n_414),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_450),
.B(n_409),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_466),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_448),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_444),
.B(n_379),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_472),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_468),
.B(n_384),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_435),
.B(n_439),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_457),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_480),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_484),
.B(n_414),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_490),
.B(n_409),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_453),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_460),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_453),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_459),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_459),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_470),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_470),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_469),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_471),
.Y(n_556)
);

NAND2x1p5_ASAP7_75t_L g557 ( 
.A(n_463),
.B(n_357),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_471),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_486),
.B(n_434),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_486),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_494),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_437),
.B(n_423),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_494),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_492),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_492),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_502),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_476),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_476),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_496),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_531),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_549),
.B(n_434),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_517),
.B(n_545),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_532),
.B(n_451),
.Y(n_573)
);

AND2x2_ASAP7_75t_SL g574 ( 
.A(n_548),
.B(n_561),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_532),
.B(n_451),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_513),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_531),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_507),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_536),
.B(n_427),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_518),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_562),
.B(n_423),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_545),
.B(n_434),
.Y(n_582)
);

INVxp33_ASAP7_75t_L g583 ( 
.A(n_540),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_536),
.B(n_374),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_509),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_509),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_560),
.B(n_374),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_513),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_522),
.B(n_385),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_522),
.B(n_385),
.Y(n_590)
);

BUFx4f_ASAP7_75t_L g591 ( 
.A(n_548),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_541),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_550),
.B(n_546),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_507),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_546),
.B(n_434),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_529),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_562),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_562),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_514),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_514),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_529),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_559),
.B(n_501),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_513),
.B(n_474),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_553),
.B(n_501),
.Y(n_604)
);

NAND2x1p5_ASAP7_75t_L g605 ( 
.A(n_561),
.B(n_357),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_543),
.B(n_385),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_543),
.B(n_428),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_567),
.B(n_428),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_567),
.B(n_428),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_518),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_516),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_553),
.B(n_449),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_555),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_518),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_540),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_563),
.B(n_428),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_518),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_537),
.B(n_479),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_547),
.B(n_481),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_568),
.B(n_432),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_518),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_563),
.B(n_432),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_516),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_520),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_520),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_521),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_521),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_568),
.B(n_432),
.Y(n_628)
);

AND2x2_ASAP7_75t_SL g629 ( 
.A(n_564),
.B(n_432),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_566),
.B(n_449),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_555),
.B(n_475),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_523),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_523),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_506),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_508),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_557),
.B(n_456),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_564),
.B(n_373),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_524),
.Y(n_638)
);

NAND3xp33_ASAP7_75t_SL g639 ( 
.A(n_569),
.B(n_452),
.C(n_489),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_557),
.B(n_488),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_508),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_519),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_519),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_551),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_524),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_526),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_526),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_527),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_527),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_557),
.A2(n_431),
.B(n_425),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_528),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_565),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_528),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_566),
.B(n_456),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_565),
.B(n_366),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_511),
.B(n_473),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_635),
.Y(n_657)
);

INVxp67_ASAP7_75t_SL g658 ( 
.A(n_597),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_597),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_577),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_570),
.Y(n_661)
);

BUFx5_ASAP7_75t_L g662 ( 
.A(n_577),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_615),
.B(n_512),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_584),
.B(n_552),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_584),
.B(n_554),
.Y(n_665)
);

AND2x6_ASAP7_75t_L g666 ( 
.A(n_581),
.B(n_519),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_598),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_577),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_570),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_578),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_652),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_574),
.B(n_569),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_635),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_618),
.B(n_556),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_577),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_621),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_642),
.B(n_643),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_615),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_574),
.B(n_530),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_621),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_592),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_642),
.B(n_643),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_606),
.B(n_558),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_578),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_652),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_578),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_642),
.B(n_544),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_578),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_621),
.Y(n_689)
);

BUFx12f_ASAP7_75t_L g690 ( 
.A(n_642),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_606),
.B(n_461),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_594),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_642),
.B(n_643),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_642),
.B(n_643),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_574),
.B(n_512),
.Y(n_695)
);

BUFx4f_ASAP7_75t_L g696 ( 
.A(n_574),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_573),
.B(n_535),
.Y(n_697)
);

INVx6_ASAP7_75t_L g698 ( 
.A(n_643),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_606),
.B(n_461),
.Y(n_699)
);

INVx6_ASAP7_75t_L g700 ( 
.A(n_643),
.Y(n_700)
);

BUFx8_ASAP7_75t_L g701 ( 
.A(n_579),
.Y(n_701)
);

OR2x6_ASAP7_75t_SL g702 ( 
.A(n_619),
.B(n_535),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_585),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_621),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_573),
.B(n_542),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_585),
.Y(n_706)
);

NAND2x1_ASAP7_75t_SL g707 ( 
.A(n_634),
.B(n_573),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_598),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_585),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_619),
.B(n_487),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_575),
.B(n_542),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_586),
.Y(n_712)
);

CKINVDCx8_ASAP7_75t_R g713 ( 
.A(n_581),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_586),
.Y(n_714)
);

AND2x2_ASAP7_75t_SL g715 ( 
.A(n_591),
.B(n_420),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_621),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_607),
.B(n_409),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_586),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_599),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_599),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_641),
.B(n_525),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_607),
.B(n_409),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_621),
.Y(n_723)
);

AND2x6_ASAP7_75t_L g724 ( 
.A(n_581),
.B(n_533),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_591),
.B(n_505),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_576),
.B(n_539),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_575),
.B(n_447),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_641),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_594),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_599),
.Y(n_730)
);

AO21x2_ASAP7_75t_L g731 ( 
.A1(n_650),
.A2(n_534),
.B(n_533),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_607),
.B(n_416),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_SL g733 ( 
.A(n_634),
.B(n_538),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_592),
.Y(n_734)
);

NAND2x1p5_ASAP7_75t_L g735 ( 
.A(n_591),
.B(n_510),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_572),
.B(n_416),
.Y(n_736)
);

NAND2x2_ASAP7_75t_L g737 ( 
.A(n_603),
.B(n_483),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_581),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_591),
.Y(n_739)
);

NOR2x1_ASAP7_75t_SL g740 ( 
.A(n_621),
.B(n_534),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_572),
.B(n_629),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_575),
.B(n_366),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_621),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_629),
.B(n_416),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_581),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_600),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_600),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_576),
.B(n_588),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_600),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_621),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_596),
.Y(n_751)
);

INVx3_ASAP7_75t_SL g752 ( 
.A(n_673),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_738),
.Y(n_753)
);

INVxp67_ASAP7_75t_SL g754 ( 
.A(n_660),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_703),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_660),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_670),
.Y(n_757)
);

INVx8_ASAP7_75t_L g758 ( 
.A(n_666),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_728),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_689),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_663),
.B(n_640),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_689),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_690),
.Y(n_763)
);

NAND2x1p5_ASAP7_75t_L g764 ( 
.A(n_660),
.B(n_668),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_728),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_706),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_689),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_709),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_738),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_670),
.Y(n_770)
);

INVx3_ASAP7_75t_SL g771 ( 
.A(n_673),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_690),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_659),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_698),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_742),
.B(n_579),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_712),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_668),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_657),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_678),
.Y(n_779)
);

INVx8_ASAP7_75t_L g780 ( 
.A(n_666),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_659),
.Y(n_781)
);

CKINVDCx16_ASAP7_75t_R g782 ( 
.A(n_657),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_714),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_695),
.A2(n_697),
.B1(n_672),
.B2(n_705),
.Y(n_784)
);

BUFx12f_ASAP7_75t_L g785 ( 
.A(n_701),
.Y(n_785)
);

NAND2x1p5_ASAP7_75t_L g786 ( 
.A(n_668),
.B(n_591),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_689),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_681),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_675),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_718),
.Y(n_790)
);

BUFx12f_ASAP7_75t_L g791 ( 
.A(n_701),
.Y(n_791)
);

CKINVDCx6p67_ASAP7_75t_R g792 ( 
.A(n_666),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_684),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_719),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_701),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_675),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_720),
.Y(n_797)
);

INVx3_ASAP7_75t_SL g798 ( 
.A(n_666),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_684),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_730),
.Y(n_800)
);

BUFx8_ASAP7_75t_L g801 ( 
.A(n_666),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_746),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_667),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_734),
.Y(n_804)
);

INVx3_ASAP7_75t_SL g805 ( 
.A(n_666),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_667),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_675),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_686),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_747),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_745),
.B(n_576),
.Y(n_810)
);

BUFx4_ASAP7_75t_SL g811 ( 
.A(n_663),
.Y(n_811)
);

CKINVDCx14_ASAP7_75t_R g812 ( 
.A(n_721),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_726),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_726),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_662),
.B(n_713),
.Y(n_815)
);

CKINVDCx16_ASAP7_75t_R g816 ( 
.A(n_727),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_745),
.B(n_576),
.Y(n_817)
);

BUFx12f_ASAP7_75t_L g818 ( 
.A(n_726),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_710),
.B(n_583),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_749),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_708),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_708),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_696),
.B(n_629),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_661),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_669),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_689),
.Y(n_826)
);

BUFx12f_ASAP7_75t_L g827 ( 
.A(n_677),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_677),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_696),
.B(n_629),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_736),
.A2(n_650),
.B(n_625),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_686),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_696),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_688),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_727),
.B(n_579),
.Y(n_834)
);

BUFx4f_ASAP7_75t_L g835 ( 
.A(n_724),
.Y(n_835)
);

INVxp67_ASAP7_75t_SL g836 ( 
.A(n_662),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_750),
.Y(n_837)
);

INVx8_ASAP7_75t_L g838 ( 
.A(n_724),
.Y(n_838)
);

NAND2x1p5_ASAP7_75t_L g839 ( 
.A(n_739),
.B(n_633),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_677),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_750),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_688),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_682),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_698),
.Y(n_844)
);

AND2x2_ASAP7_75t_SL g845 ( 
.A(n_715),
.B(n_602),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_824),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_824),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_827),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_845),
.A2(n_695),
.B1(n_697),
.B2(n_705),
.Y(n_849)
);

CKINVDCx11_ASAP7_75t_R g850 ( 
.A(n_795),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_825),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_825),
.Y(n_852)
);

BUFx2_ASAP7_75t_SL g853 ( 
.A(n_763),
.Y(n_853)
);

BUFx4f_ASAP7_75t_SL g854 ( 
.A(n_785),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_845),
.A2(n_711),
.B1(n_440),
.B2(n_442),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_773),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_845),
.A2(n_639),
.B1(n_737),
.B2(n_583),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_755),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_757),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_773),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_782),
.Y(n_861)
);

INVx6_ASAP7_75t_L g862 ( 
.A(n_827),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_781),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_812),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_757),
.Y(n_865)
);

CKINVDCx14_ASAP7_75t_R g866 ( 
.A(n_778),
.Y(n_866)
);

BUFx10_ASAP7_75t_L g867 ( 
.A(n_778),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_770),
.Y(n_868)
);

CKINVDCx6p67_ASAP7_75t_R g869 ( 
.A(n_752),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_755),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_835),
.A2(n_715),
.B1(n_665),
.B2(n_664),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_835),
.A2(n_644),
.B1(n_683),
.B2(n_741),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_834),
.A2(n_711),
.B1(n_672),
.B2(n_737),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_SL g874 ( 
.A1(n_816),
.A2(n_702),
.B1(n_733),
.B2(n_679),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_834),
.A2(n_602),
.B1(n_639),
.B2(n_630),
.Y(n_875)
);

INVx1_ASAP7_75t_SL g876 ( 
.A(n_759),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_835),
.A2(n_644),
.B1(n_713),
.B2(n_674),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_788),
.A2(n_804),
.B1(n_775),
.B2(n_819),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_766),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_SL g880 ( 
.A1(n_765),
.A2(n_515),
.B(n_604),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_766),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_779),
.A2(n_744),
.B1(n_691),
.B2(n_699),
.Y(n_882)
);

BUFx8_ASAP7_75t_L g883 ( 
.A(n_785),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_768),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_SL g885 ( 
.A1(n_836),
.A2(n_739),
.B(n_693),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_784),
.A2(n_654),
.B1(n_630),
.B2(n_636),
.Y(n_886)
);

AO22x1_ASAP7_75t_L g887 ( 
.A1(n_801),
.A2(n_679),
.B1(n_640),
.B2(n_654),
.Y(n_887)
);

CKINVDCx6p67_ASAP7_75t_R g888 ( 
.A(n_752),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_768),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_761),
.A2(n_636),
.B1(n_445),
.B2(n_515),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_761),
.A2(n_445),
.B1(n_446),
.B2(n_702),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_781),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_776),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_770),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_776),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_783),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_752),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_783),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_793),
.Y(n_899)
);

INVx8_ASAP7_75t_L g900 ( 
.A(n_838),
.Y(n_900)
);

BUFx8_ASAP7_75t_L g901 ( 
.A(n_791),
.Y(n_901)
);

INVx1_ASAP7_75t_SL g902 ( 
.A(n_771),
.Y(n_902)
);

INVx6_ASAP7_75t_L g903 ( 
.A(n_801),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_782),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_818),
.A2(n_631),
.B1(n_604),
.B2(n_612),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_793),
.Y(n_906)
);

INVx8_ASAP7_75t_L g907 ( 
.A(n_838),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_SL g908 ( 
.A1(n_816),
.A2(n_605),
.B1(n_603),
.B2(n_582),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_803),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_821),
.A2(n_658),
.B1(n_722),
.B2(n_717),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_818),
.A2(n_612),
.B1(n_605),
.B2(n_364),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_790),
.Y(n_912)
);

BUFx8_ASAP7_75t_L g913 ( 
.A(n_791),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_813),
.A2(n_605),
.B1(n_395),
.B2(n_388),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_803),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_771),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_821),
.A2(n_732),
.B1(n_588),
.B2(n_576),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_790),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_794),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_794),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_799),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_797),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_814),
.A2(n_605),
.B1(n_623),
.B2(n_611),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_811),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_771),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_797),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_799),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_838),
.Y(n_928)
);

BUFx4f_ASAP7_75t_SL g929 ( 
.A(n_806),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_823),
.A2(n_605),
.B1(n_623),
.B2(n_611),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_822),
.B(n_707),
.Y(n_931)
);

OAI22xp33_ASAP7_75t_L g932 ( 
.A1(n_838),
.A2(n_685),
.B1(n_671),
.B2(n_656),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_806),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_822),
.B(n_655),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_800),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_823),
.A2(n_623),
.B1(n_627),
.B2(n_611),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_829),
.A2(n_623),
.B1(n_627),
.B2(n_611),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_SL g938 ( 
.A1(n_829),
.A2(n_581),
.B(n_404),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_SL g939 ( 
.A1(n_838),
.A2(n_582),
.B1(n_571),
.B2(n_662),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_753),
.Y(n_940)
);

OAI22xp33_ASAP7_75t_R g941 ( 
.A1(n_800),
.A2(n_410),
.B1(n_38),
.B2(n_35),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_SL g942 ( 
.A1(n_801),
.A2(n_571),
.B1(n_662),
.B2(n_698),
.Y(n_942)
);

INVx6_ASAP7_75t_L g943 ( 
.A(n_801),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_808),
.Y(n_944)
);

INVx4_ASAP7_75t_L g945 ( 
.A(n_828),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_763),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_753),
.B(n_593),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_810),
.A2(n_632),
.B1(n_645),
.B2(n_627),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_810),
.A2(n_632),
.B1(n_645),
.B2(n_627),
.Y(n_949)
);

CKINVDCx11_ASAP7_75t_R g950 ( 
.A(n_772),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_808),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_769),
.B(n_655),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_772),
.Y(n_953)
);

CKINVDCx11_ASAP7_75t_R g954 ( 
.A(n_760),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_SL g955 ( 
.A1(n_810),
.A2(n_595),
.B(n_748),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_954),
.Y(n_956)
);

OAI22xp33_ASAP7_75t_L g957 ( 
.A1(n_857),
.A2(n_769),
.B1(n_832),
.B2(n_805),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_855),
.A2(n_810),
.B1(n_817),
.B2(n_786),
.Y(n_958)
);

OAI22xp33_ASAP7_75t_L g959 ( 
.A1(n_938),
.A2(n_832),
.B1(n_798),
.B2(n_805),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_855),
.A2(n_595),
.B1(n_817),
.B2(n_780),
.Y(n_960)
);

OAI21xp33_ASAP7_75t_L g961 ( 
.A1(n_875),
.A2(n_809),
.B(n_802),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_856),
.B(n_828),
.Y(n_962)
);

OAI22xp33_ASAP7_75t_L g963 ( 
.A1(n_880),
.A2(n_805),
.B1(n_798),
.B2(n_840),
.Y(n_963)
);

AND2x2_ASAP7_75t_SL g964 ( 
.A(n_930),
.B(n_682),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_858),
.B(n_802),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_856),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_890),
.A2(n_817),
.B1(n_780),
.B2(n_758),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_SL g968 ( 
.A1(n_882),
.A2(n_780),
.B1(n_758),
.B2(n_682),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_954),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_940),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_SL g971 ( 
.A1(n_877),
.A2(n_780),
.B1(n_758),
.B2(n_693),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_890),
.A2(n_817),
.B1(n_780),
.B2(n_758),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_859),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_849),
.A2(n_874),
.B1(n_891),
.B2(n_941),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_929),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_875),
.B(n_809),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_873),
.A2(n_786),
.B1(n_820),
.B2(n_840),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_876),
.B(n_400),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_910),
.A2(n_830),
.B(n_725),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_878),
.B(n_820),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_903),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_SL g982 ( 
.A1(n_873),
.A2(n_694),
.B(n_693),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_871),
.A2(n_786),
.B1(n_843),
.B2(n_756),
.Y(n_983)
);

CKINVDCx14_ASAP7_75t_R g984 ( 
.A(n_850),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_849),
.A2(n_758),
.B1(n_792),
.B2(n_798),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_870),
.B(n_731),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_859),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_900),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_947),
.B(n_886),
.Y(n_989)
);

CKINVDCx16_ASAP7_75t_R g990 ( 
.A(n_861),
.Y(n_990)
);

OAI222xp33_ASAP7_75t_L g991 ( 
.A1(n_891),
.A2(n_593),
.B1(n_656),
.B2(n_842),
.C1(n_831),
.C2(n_833),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_931),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_886),
.B(n_831),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_908),
.A2(n_792),
.B1(n_687),
.B2(n_843),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_850),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_902),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_945),
.B(n_826),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_903),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_905),
.A2(n_833),
.B1(n_694),
.B2(n_624),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_SL g1000 ( 
.A1(n_872),
.A2(n_694),
.B1(n_700),
.B2(n_698),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_905),
.A2(n_911),
.B1(n_914),
.B2(n_932),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_911),
.A2(n_807),
.B1(n_754),
.B2(n_748),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_914),
.A2(n_624),
.B1(n_626),
.B2(n_625),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_879),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_SL g1005 ( 
.A1(n_955),
.A2(n_609),
.B(n_608),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_881),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_860),
.B(n_842),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_930),
.A2(n_624),
.B1(n_626),
.B2(n_625),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_903),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_864),
.B(n_400),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_948),
.A2(n_748),
.B1(n_588),
.B2(n_764),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_923),
.A2(n_626),
.B1(n_638),
.B2(n_648),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_948),
.A2(n_588),
.B1(n_764),
.B2(n_777),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_884),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_889),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_865),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_923),
.A2(n_638),
.B1(n_649),
.B2(n_648),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_893),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_939),
.A2(n_638),
.B1(n_649),
.B2(n_648),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_SL g1020 ( 
.A1(n_866),
.A2(n_609),
.B(n_608),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_895),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_865),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_883),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_896),
.B(n_731),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_863),
.Y(n_1025)
);

CKINVDCx11_ASAP7_75t_R g1026 ( 
.A(n_904),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_900),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_862),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_898),
.Y(n_1029)
);

OAI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_949),
.A2(n_392),
.B(n_410),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_952),
.A2(n_648),
.B1(n_651),
.B2(n_649),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_943),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_SL g1033 ( 
.A1(n_866),
.A2(n_400),
.B1(n_735),
.B2(n_700),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_892),
.Y(n_1034)
);

BUFx12f_ASAP7_75t_L g1035 ( 
.A(n_883),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_943),
.Y(n_1036)
);

AOI222xp33_ASAP7_75t_L g1037 ( 
.A1(n_887),
.A2(n_628),
.B1(n_620),
.B2(n_609),
.C1(n_608),
.C2(n_637),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_912),
.B(n_731),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_909),
.B(n_777),
.Y(n_1039)
);

BUFx4f_ASAP7_75t_SL g1040 ( 
.A(n_883),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_915),
.B(n_777),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_943),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_868),
.Y(n_1043)
);

OAI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_924),
.A2(n_588),
.B1(n_700),
.B2(n_735),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_SL g1045 ( 
.A1(n_848),
.A2(n_628),
.B(n_620),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_934),
.A2(n_649),
.B1(n_653),
.B2(n_651),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_974),
.A2(n_917),
.B1(n_937),
.B2(n_936),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_970),
.B(n_933),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1004),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_1001),
.A2(n_942),
.B1(n_894),
.B2(n_899),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_986),
.B(n_918),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_980),
.B(n_846),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_960),
.A2(n_894),
.B1(n_899),
.B2(n_868),
.Y(n_1053)
);

AOI222xp33_ASAP7_75t_L g1054 ( 
.A1(n_991),
.A2(n_392),
.B1(n_628),
.B2(n_620),
.C1(n_851),
.C2(n_847),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_SL g1055 ( 
.A1(n_958),
.A2(n_862),
.B1(n_852),
.B2(n_853),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_963),
.A2(n_921),
.B1(n_927),
.B2(n_906),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_SL g1057 ( 
.A1(n_964),
.A2(n_862),
.B1(n_920),
.B2(n_919),
.Y(n_1057)
);

AOI221xp5_ASAP7_75t_L g1058 ( 
.A1(n_961),
.A2(n_369),
.B1(n_375),
.B2(n_376),
.C(n_381),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_SL g1059 ( 
.A1(n_964),
.A2(n_922),
.B1(n_935),
.B2(n_926),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_967),
.A2(n_906),
.B1(n_927),
.B2(n_921),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_SL g1061 ( 
.A1(n_964),
.A2(n_848),
.B1(n_913),
.B2(n_901),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_972),
.A2(n_951),
.B1(n_944),
.B2(n_936),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1005),
.A2(n_949),
.B1(n_916),
.B2(n_888),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_986),
.B(n_937),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_SL g1065 ( 
.A1(n_976),
.A2(n_901),
.B1(n_913),
.B2(n_854),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1037),
.A2(n_944),
.B1(n_951),
.B2(n_946),
.Y(n_1066)
);

OAI221xp5_ASAP7_75t_L g1067 ( 
.A1(n_1020),
.A2(n_953),
.B1(n_369),
.B2(n_375),
.C(n_376),
.Y(n_1067)
);

AOI221xp5_ASAP7_75t_L g1068 ( 
.A1(n_961),
.A2(n_989),
.B1(n_978),
.B2(n_381),
.C(n_1010),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_959),
.A2(n_950),
.B1(n_725),
.B2(n_653),
.Y(n_1069)
);

OAI221xp5_ASAP7_75t_SL g1070 ( 
.A1(n_1045),
.A2(n_392),
.B1(n_869),
.B2(n_637),
.C(n_885),
.Y(n_1070)
);

AND2x2_ASAP7_75t_SL g1071 ( 
.A(n_956),
.B(n_928),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_992),
.A2(n_950),
.B1(n_653),
.B2(n_651),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_968),
.A2(n_653),
.B1(n_651),
.B2(n_815),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_977),
.A2(n_700),
.B1(n_692),
.B2(n_751),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1024),
.B(n_826),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_SL g1076 ( 
.A1(n_993),
.A2(n_913),
.B1(n_901),
.B2(n_900),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_SL g1077 ( 
.A1(n_1033),
.A2(n_907),
.B1(n_945),
.B2(n_928),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_957),
.A2(n_729),
.B1(n_692),
.B2(n_596),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_982),
.A2(n_925),
.B1(n_897),
.B2(n_764),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_997),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_999),
.A2(n_601),
.B1(n_596),
.B2(n_907),
.Y(n_1081)
);

OAI222xp33_ASAP7_75t_L g1082 ( 
.A1(n_994),
.A2(n_587),
.B1(n_613),
.B2(n_601),
.C1(n_596),
.C2(n_844),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1004),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_965),
.B(n_789),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_SL g1085 ( 
.A1(n_1003),
.A2(n_839),
.B(n_622),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1008),
.A2(n_839),
.B1(n_789),
.B2(n_796),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1024),
.A2(n_601),
.B1(n_907),
.B2(n_646),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_SL g1088 ( 
.A1(n_983),
.A2(n_844),
.B(n_774),
.Y(n_1088)
);

AO22x1_ASAP7_75t_L g1089 ( 
.A1(n_956),
.A2(n_826),
.B1(n_837),
.B2(n_774),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1038),
.A2(n_601),
.B1(n_646),
.B2(n_724),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1038),
.A2(n_646),
.B1(n_724),
.B2(n_662),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_SL g1092 ( 
.A1(n_979),
.A2(n_662),
.B1(n_587),
.B2(n_408),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1006),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_985),
.A2(n_646),
.B1(n_724),
.B2(n_662),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_SL g1095 ( 
.A1(n_1028),
.A2(n_587),
.B1(n_415),
.B2(n_411),
.Y(n_1095)
);

OAI221xp5_ASAP7_75t_SL g1096 ( 
.A1(n_1030),
.A2(n_637),
.B1(n_590),
.B2(n_589),
.C(n_613),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1030),
.A2(n_646),
.B1(n_724),
.B2(n_633),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1006),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1035),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1014),
.Y(n_1100)
);

OA21x2_ASAP7_75t_L g1101 ( 
.A1(n_1014),
.A2(n_613),
.B(n_356),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1012),
.A2(n_646),
.B1(n_633),
.B2(n_415),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1017),
.A2(n_646),
.B1(n_633),
.B2(n_415),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1031),
.A2(n_646),
.B1(n_633),
.B2(n_415),
.Y(n_1104)
);

OAI21xp33_ASAP7_75t_L g1105 ( 
.A1(n_965),
.A2(n_411),
.B(n_415),
.Y(n_1105)
);

OA222x2_ASAP7_75t_L g1106 ( 
.A1(n_1007),
.A2(n_796),
.B1(n_789),
.B2(n_837),
.C1(n_647),
.C2(n_617),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1046),
.A2(n_646),
.B1(n_633),
.B2(n_411),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_1025),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_971),
.A2(n_633),
.B1(n_411),
.B2(n_647),
.Y(n_1109)
);

AOI221xp5_ASAP7_75t_SL g1110 ( 
.A1(n_996),
.A2(n_424),
.B1(n_433),
.B2(n_411),
.C(n_41),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1075),
.B(n_1051),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_L g1112 ( 
.A(n_1068),
.B(n_1034),
.C(n_1039),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1108),
.B(n_966),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1075),
.B(n_1015),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1052),
.B(n_1051),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_1071),
.B(n_956),
.Y(n_1116)
);

NOR3xp33_ASAP7_75t_L g1117 ( 
.A(n_1070),
.B(n_966),
.C(n_1041),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1096),
.A2(n_990),
.B1(n_1000),
.B2(n_984),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1049),
.B(n_1015),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1049),
.B(n_1018),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1066),
.A2(n_1002),
.B1(n_962),
.B2(n_987),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1048),
.B(n_1083),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_SL g1123 ( 
.A1(n_1063),
.A2(n_969),
.B(n_1040),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1093),
.B(n_1021),
.Y(n_1124)
);

NAND4xp25_ASAP7_75t_L g1125 ( 
.A(n_1067),
.B(n_975),
.C(n_1021),
.D(n_1029),
.Y(n_1125)
);

OAI221xp5_ASAP7_75t_L g1126 ( 
.A1(n_1110),
.A2(n_1028),
.B1(n_1029),
.B2(n_1042),
.C(n_1019),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1047),
.A2(n_1085),
.B1(n_1059),
.B2(n_1069),
.Y(n_1127)
);

AND4x1_ASAP7_75t_L g1128 ( 
.A(n_1088),
.B(n_1035),
.C(n_1023),
.D(n_1026),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1093),
.B(n_969),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1098),
.B(n_969),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1047),
.A2(n_1011),
.B1(n_1013),
.B2(n_990),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_L g1132 ( 
.A(n_1072),
.B(n_411),
.C(n_1026),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1098),
.B(n_962),
.Y(n_1133)
);

NAND3xp33_ASAP7_75t_L g1134 ( 
.A(n_1054),
.B(n_995),
.C(n_962),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1085),
.A2(n_1057),
.B1(n_1061),
.B2(n_1055),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1100),
.B(n_997),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1076),
.B(n_1042),
.Y(n_1137)
);

NAND4xp25_ASAP7_75t_L g1138 ( 
.A(n_1079),
.B(n_975),
.C(n_416),
.D(n_997),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1100),
.B(n_998),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_L g1140 ( 
.A(n_1092),
.B(n_995),
.C(n_981),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1064),
.B(n_1080),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_L g1142 ( 
.A(n_1058),
.B(n_981),
.C(n_998),
.Y(n_1142)
);

OAI221xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1088),
.A2(n_1044),
.B1(n_1036),
.B2(n_1032),
.C(n_1009),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1065),
.B(n_981),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1064),
.B(n_973),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_L g1146 ( 
.A(n_1097),
.B(n_1009),
.C(n_998),
.Y(n_1146)
);

NOR3xp33_ASAP7_75t_SL g1147 ( 
.A(n_1099),
.B(n_867),
.C(n_1023),
.Y(n_1147)
);

AOI221xp5_ASAP7_75t_L g1148 ( 
.A1(n_1084),
.A2(n_424),
.B1(n_433),
.B2(n_260),
.C(n_262),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_L g1149 ( 
.A(n_1105),
.B(n_1036),
.C(n_1032),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1080),
.B(n_1032),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_L g1151 ( 
.A(n_1089),
.B(n_1036),
.C(n_796),
.Y(n_1151)
);

OAI221xp5_ASAP7_75t_L g1152 ( 
.A1(n_1073),
.A2(n_250),
.B1(n_305),
.B2(n_254),
.C(n_264),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1089),
.B(n_973),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1086),
.B(n_987),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_SL g1155 ( 
.A1(n_1106),
.A2(n_988),
.B1(n_1027),
.B2(n_1022),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1050),
.B(n_1016),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1074),
.B(n_1016),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1060),
.A2(n_1043),
.B1(n_1022),
.B2(n_633),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1111),
.B(n_1106),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1119),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1113),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1127),
.A2(n_1105),
.B1(n_1077),
.B2(n_1056),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1115),
.B(n_1101),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_L g1164 ( 
.A(n_1155),
.B(n_1087),
.C(n_1078),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_SL g1165 ( 
.A1(n_1135),
.A2(n_1101),
.B1(n_1099),
.B2(n_988),
.Y(n_1165)
);

NAND4xp75_ASAP7_75t_L g1166 ( 
.A(n_1131),
.B(n_1101),
.C(n_1082),
.D(n_1043),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1118),
.A2(n_433),
.B1(n_424),
.B2(n_291),
.C(n_293),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_1111),
.B(n_1101),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1141),
.B(n_1091),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1114),
.B(n_1053),
.Y(n_1170)
);

AND2x2_ASAP7_75t_SL g1171 ( 
.A(n_1128),
.B(n_988),
.Y(n_1171)
);

NAND4xp75_ASAP7_75t_L g1172 ( 
.A(n_1137),
.B(n_1144),
.C(n_1131),
.D(n_1116),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1141),
.B(n_867),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1128),
.B(n_988),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1114),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1136),
.B(n_1090),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1136),
.B(n_1094),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_L g1178 ( 
.A(n_1138),
.B(n_1095),
.C(n_837),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1129),
.B(n_1109),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1129),
.B(n_760),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_1112),
.B(n_1081),
.C(n_1062),
.Y(n_1181)
);

NOR3xp33_ASAP7_75t_L g1182 ( 
.A(n_1125),
.B(n_647),
.C(n_617),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1120),
.Y(n_1183)
);

NAND4xp75_ASAP7_75t_L g1184 ( 
.A(n_1153),
.B(n_422),
.C(n_348),
.D(n_356),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1120),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1122),
.B(n_1102),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1117),
.B(n_1104),
.C(n_1107),
.Y(n_1187)
);

NAND4xp75_ASAP7_75t_L g1188 ( 
.A(n_1147),
.B(n_1027),
.C(n_988),
.D(n_589),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1134),
.A2(n_424),
.B1(n_433),
.B2(n_299),
.C(n_300),
.Y(n_1189)
);

NAND4xp75_ASAP7_75t_L g1190 ( 
.A(n_1156),
.B(n_422),
.C(n_348),
.D(n_356),
.Y(n_1190)
);

AOI221xp5_ASAP7_75t_L g1191 ( 
.A1(n_1134),
.A2(n_433),
.B1(n_282),
.B2(n_303),
.C(n_304),
.Y(n_1191)
);

XNOR2xp5_ASAP7_75t_L g1192 ( 
.A(n_1130),
.B(n_36),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1124),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1145),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1132),
.A2(n_1103),
.B1(n_633),
.B2(n_273),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1133),
.B(n_1139),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1150),
.B(n_38),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1154),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1157),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_L g1200 ( 
.A(n_1151),
.B(n_1027),
.C(n_762),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1146),
.Y(n_1201)
);

OAI211xp5_ASAP7_75t_SL g1202 ( 
.A1(n_1123),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_1202)
);

NAND4xp25_ASAP7_75t_L g1203 ( 
.A(n_1126),
.B(n_40),
.C(n_42),
.D(n_44),
.Y(n_1203)
);

NOR3xp33_ASAP7_75t_SL g1204 ( 
.A(n_1143),
.B(n_266),
.C(n_44),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1140),
.A2(n_839),
.B(n_377),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1146),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1121),
.B(n_46),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1149),
.B(n_46),
.Y(n_1208)
);

XNOR2x2_ASAP7_75t_L g1209 ( 
.A(n_1192),
.B(n_1149),
.Y(n_1209)
);

AO22x2_ASAP7_75t_L g1210 ( 
.A1(n_1199),
.A2(n_1142),
.B1(n_1158),
.B2(n_1148),
.Y(n_1210)
);

XNOR2xp5_ASAP7_75t_L g1211 ( 
.A(n_1192),
.B(n_1172),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1206),
.A2(n_1152),
.B1(n_405),
.B2(n_386),
.Y(n_1212)
);

XNOR2xp5_ASAP7_75t_L g1213 ( 
.A(n_1171),
.B(n_47),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1162),
.A2(n_1027),
.B1(n_841),
.B2(n_787),
.Y(n_1214)
);

XNOR2x2_ASAP7_75t_L g1215 ( 
.A(n_1166),
.B(n_48),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1201),
.B(n_49),
.Y(n_1216)
);

NOR3xp33_ASAP7_75t_L g1217 ( 
.A(n_1203),
.B(n_50),
.C(n_53),
.Y(n_1217)
);

OA22x2_ASAP7_75t_L g1218 ( 
.A1(n_1159),
.A2(n_655),
.B1(n_647),
.B2(n_704),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1175),
.B(n_50),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1166),
.A2(n_273),
.B1(n_655),
.B2(n_767),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1171),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1198),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1165),
.A2(n_273),
.B1(n_655),
.B2(n_767),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1168),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1159),
.B(n_760),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1193),
.Y(n_1226)
);

NAND4xp75_ASAP7_75t_SL g1227 ( 
.A(n_1174),
.B(n_1188),
.C(n_1173),
.D(n_1202),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1168),
.Y(n_1228)
);

XOR2x2_ASAP7_75t_L g1229 ( 
.A(n_1207),
.B(n_54),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1161),
.B(n_56),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1204),
.A2(n_841),
.B1(n_787),
.B2(n_767),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1173),
.B(n_56),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1196),
.B(n_57),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1208),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1174),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1160),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1181),
.A2(n_1164),
.B1(n_1207),
.B2(n_1187),
.Y(n_1237)
);

XNOR2xp5_ASAP7_75t_L g1238 ( 
.A(n_1211),
.B(n_1188),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1219),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1226),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1224),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1222),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1233),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_1213),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1221),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1221),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1236),
.Y(n_1247)
);

AO22x2_ASAP7_75t_L g1248 ( 
.A1(n_1234),
.A2(n_1170),
.B1(n_1163),
.B2(n_1186),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_1216),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1230),
.Y(n_1250)
);

XOR2x2_ASAP7_75t_L g1251 ( 
.A(n_1229),
.B(n_1189),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1224),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1228),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1234),
.Y(n_1254)
);

XOR2x2_ASAP7_75t_L g1255 ( 
.A(n_1229),
.B(n_1191),
.Y(n_1255)
);

XOR2xp5_ASAP7_75t_L g1256 ( 
.A(n_1209),
.B(n_1197),
.Y(n_1256)
);

INVx5_ASAP7_75t_L g1257 ( 
.A(n_1235),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1228),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1225),
.Y(n_1259)
);

AO22x2_ASAP7_75t_L g1260 ( 
.A1(n_1217),
.A2(n_1200),
.B1(n_1169),
.B2(n_1176),
.Y(n_1260)
);

XNOR2x2_ASAP7_75t_L g1261 ( 
.A(n_1215),
.B(n_1167),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1218),
.Y(n_1262)
);

AOI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1217),
.A2(n_1182),
.B1(n_1176),
.B2(n_1177),
.Y(n_1263)
);

OA22x2_ASAP7_75t_L g1264 ( 
.A1(n_1256),
.A2(n_1220),
.B1(n_1223),
.B2(n_1214),
.Y(n_1264)
);

CKINVDCx16_ASAP7_75t_R g1265 ( 
.A(n_1238),
.Y(n_1265)
);

AO22x2_ASAP7_75t_L g1266 ( 
.A1(n_1256),
.A2(n_1227),
.B1(n_1237),
.B2(n_1210),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_1260),
.Y(n_1267)
);

AO22x2_ASAP7_75t_L g1268 ( 
.A1(n_1249),
.A2(n_1210),
.B1(n_1194),
.B2(n_1179),
.Y(n_1268)
);

OA22x2_ASAP7_75t_L g1269 ( 
.A1(n_1263),
.A2(n_1177),
.B1(n_1194),
.B2(n_1205),
.Y(n_1269)
);

INVx5_ASAP7_75t_L g1270 ( 
.A(n_1257),
.Y(n_1270)
);

OA22x2_ASAP7_75t_L g1271 ( 
.A1(n_1250),
.A2(n_1179),
.B1(n_1183),
.B2(n_1185),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1260),
.A2(n_1210),
.B1(n_1212),
.B2(n_1232),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1247),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1260),
.A2(n_1180),
.B1(n_1231),
.B2(n_1195),
.Y(n_1274)
);

INVx4_ASAP7_75t_R g1275 ( 
.A(n_1239),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1244),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1245),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1240),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1254),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1243),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1242),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1258),
.Y(n_1282)
);

OA22x2_ASAP7_75t_L g1283 ( 
.A1(n_1262),
.A2(n_1180),
.B1(n_1178),
.B2(n_1190),
.Y(n_1283)
);

XOR2x2_ASAP7_75t_L g1284 ( 
.A(n_1251),
.B(n_1184),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1241),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1252),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1273),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1273),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1278),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1277),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1278),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1266),
.A2(n_1255),
.B1(n_1251),
.B2(n_1248),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1281),
.Y(n_1293)
);

OAI322xp33_ASAP7_75t_L g1294 ( 
.A1(n_1267),
.A2(n_1261),
.A3(n_1246),
.B1(n_1253),
.B2(n_1252),
.C1(n_1248),
.C2(n_1259),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1281),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1272),
.A2(n_1257),
.B1(n_1248),
.B2(n_1253),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1279),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1266),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1275),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1282),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1268),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1276),
.Y(n_1302)
);

OAI322xp33_ASAP7_75t_L g1303 ( 
.A1(n_1265),
.A2(n_1274),
.A3(n_1269),
.B1(n_1271),
.B2(n_1264),
.C1(n_1280),
.C2(n_1283),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1285),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1286),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1284),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1270),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1270),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1270),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1273),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1292),
.A2(n_1257),
.B1(n_841),
.B2(n_787),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1302),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1287),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_SL g1314 ( 
.A1(n_1299),
.A2(n_1257),
.B(n_60),
.C(n_61),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1287),
.Y(n_1315)
);

OA22x2_ASAP7_75t_L g1316 ( 
.A1(n_1296),
.A2(n_58),
.B1(n_61),
.B2(n_63),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1290),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1290),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_SL g1319 ( 
.A1(n_1307),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1298),
.A2(n_273),
.B1(n_647),
.B2(n_377),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1293),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1298),
.A2(n_841),
.B1(n_787),
.B2(n_767),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1293),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1295),
.Y(n_1324)
);

BUFx4_ASAP7_75t_R g1325 ( 
.A(n_1306),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1295),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1306),
.A2(n_273),
.B1(n_377),
.B2(n_762),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1300),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1297),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1309),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1309),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1300),
.Y(n_1332)
);

OA22x2_ASAP7_75t_L g1333 ( 
.A1(n_1301),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1288),
.Y(n_1334)
);

OA22x2_ASAP7_75t_SL g1335 ( 
.A1(n_1308),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1289),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1291),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1310),
.Y(n_1338)
);

OA22x2_ASAP7_75t_L g1339 ( 
.A1(n_1308),
.A2(n_71),
.B1(n_72),
.B2(n_616),
.Y(n_1339)
);

NAND4xp75_ASAP7_75t_L g1340 ( 
.A(n_1294),
.B(n_1303),
.C(n_1304),
.D(n_1305),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1325),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1340),
.A2(n_762),
.B1(n_760),
.B2(n_743),
.Y(n_1342)
);

INVxp67_ASAP7_75t_L g1343 ( 
.A(n_1317),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1329),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1335),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1311),
.A2(n_377),
.B1(n_405),
.B2(n_386),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1316),
.A2(n_762),
.B1(n_743),
.B2(n_676),
.Y(n_1347)
);

OA22x2_ASAP7_75t_L g1348 ( 
.A1(n_1311),
.A2(n_622),
.B1(n_616),
.B2(n_610),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1313),
.Y(n_1349)
);

AOI221xp5_ASAP7_75t_L g1350 ( 
.A1(n_1319),
.A2(n_405),
.B1(n_386),
.B2(n_622),
.C(n_616),
.Y(n_1350)
);

INVxp33_ASAP7_75t_SL g1351 ( 
.A(n_1318),
.Y(n_1351)
);

OA22x2_ASAP7_75t_L g1352 ( 
.A1(n_1330),
.A2(n_622),
.B1(n_616),
.B2(n_610),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1315),
.Y(n_1353)
);

INVxp67_ASAP7_75t_L g1354 ( 
.A(n_1339),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1314),
.A2(n_622),
.B(n_589),
.C(n_590),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1321),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1323),
.Y(n_1357)
);

AOI31xp33_ASAP7_75t_L g1358 ( 
.A1(n_1331),
.A2(n_590),
.A3(n_762),
.B(n_740),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1335),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1334),
.Y(n_1360)
);

AND4x1_ASAP7_75t_L g1361 ( 
.A(n_1327),
.B(n_81),
.C(n_82),
.D(n_86),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1324),
.Y(n_1362)
);

A2O1A1Ixp33_ASAP7_75t_SL g1363 ( 
.A1(n_1326),
.A2(n_617),
.B(n_610),
.C(n_426),
.Y(n_1363)
);

AO22x2_ASAP7_75t_L g1364 ( 
.A1(n_1336),
.A2(n_723),
.B1(n_716),
.B2(n_704),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1328),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1333),
.A2(n_377),
.B1(n_386),
.B2(n_405),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1332),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1337),
.A2(n_426),
.B(n_363),
.C(n_413),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1338),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1320),
.A2(n_377),
.B1(n_350),
.B2(n_380),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1322),
.Y(n_1371)
);

OAI22x1_ASAP7_75t_L g1372 ( 
.A1(n_1312),
.A2(n_723),
.B1(n_363),
.B2(n_617),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1325),
.Y(n_1373)
);

AO22x1_ASAP7_75t_L g1374 ( 
.A1(n_1342),
.A2(n_1345),
.B1(n_1359),
.B2(n_1373),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1342),
.A2(n_743),
.B1(n_680),
.B2(n_676),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1360),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1341),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1352),
.Y(n_1378)
);

NOR2x1_ASAP7_75t_L g1379 ( 
.A(n_1344),
.B(n_750),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1352),
.Y(n_1380)
);

AOI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1354),
.A2(n_743),
.B1(n_680),
.B2(n_676),
.Y(n_1381)
);

NOR4xp25_ASAP7_75t_L g1382 ( 
.A(n_1343),
.B(n_617),
.C(n_610),
.D(n_92),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1371),
.A2(n_350),
.B1(n_380),
.B2(n_352),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1349),
.Y(n_1384)
);

OA22x2_ASAP7_75t_L g1385 ( 
.A1(n_1369),
.A2(n_610),
.B1(n_89),
.B2(n_94),
.Y(n_1385)
);

AO22x2_ASAP7_75t_L g1386 ( 
.A1(n_1353),
.A2(n_1365),
.B1(n_1356),
.B2(n_1362),
.Y(n_1386)
);

AO22x2_ASAP7_75t_L g1387 ( 
.A1(n_1357),
.A2(n_614),
.B1(n_580),
.B2(n_99),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1347),
.A2(n_680),
.B1(n_352),
.B2(n_380),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1350),
.A2(n_352),
.B1(n_380),
.B2(n_383),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1372),
.Y(n_1390)
);

OA22x2_ASAP7_75t_L g1391 ( 
.A1(n_1367),
.A2(n_87),
.B1(n_98),
.B2(n_100),
.Y(n_1391)
);

NOR2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1351),
.B(n_750),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1355),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1348),
.A2(n_352),
.B1(n_383),
.B2(n_580),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1366),
.A2(n_383),
.B1(n_750),
.B2(n_580),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_SL g1396 ( 
.A1(n_1346),
.A2(n_1358),
.B1(n_1348),
.B2(n_1370),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1361),
.Y(n_1397)
);

NOR2xp67_ASAP7_75t_L g1398 ( 
.A(n_1363),
.B(n_103),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1364),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1368),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1342),
.A2(n_614),
.B1(n_418),
.B2(n_417),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1342),
.A2(n_614),
.B1(n_418),
.B2(n_417),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1360),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1360),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1377),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1386),
.Y(n_1406)
);

NOR3xp33_ASAP7_75t_SL g1407 ( 
.A(n_1376),
.B(n_104),
.C(n_105),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1393),
.A2(n_418),
.B1(n_417),
.B2(n_378),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1386),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1403),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1404),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1378),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1391),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1384),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1387),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1387),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1397),
.A2(n_418),
.B1(n_417),
.B2(n_378),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1380),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1374),
.B(n_106),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1374),
.B(n_1399),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1400),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1382),
.B(n_378),
.Y(n_1422)
);

NOR3xp33_ASAP7_75t_L g1423 ( 
.A(n_1396),
.B(n_108),
.C(n_109),
.Y(n_1423)
);

AND3x4_ASAP7_75t_L g1424 ( 
.A(n_1379),
.B(n_1398),
.C(n_1390),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1385),
.A2(n_378),
.B1(n_121),
.B2(n_122),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1392),
.B(n_114),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1381),
.B(n_124),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1389),
.Y(n_1428)
);

NOR2x1_ASAP7_75t_L g1429 ( 
.A(n_1394),
.B(n_125),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1395),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1388),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1383),
.Y(n_1432)
);

INVxp67_ASAP7_75t_SL g1433 ( 
.A(n_1401),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1402),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1409),
.A2(n_1375),
.B1(n_130),
.B2(n_132),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1405),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1406),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1412),
.A2(n_1408),
.B1(n_1410),
.B2(n_1411),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1420),
.Y(n_1439)
);

OA22x2_ASAP7_75t_L g1440 ( 
.A1(n_1418),
.A2(n_128),
.B1(n_133),
.B2(n_134),
.Y(n_1440)
);

AO22x2_ASAP7_75t_L g1441 ( 
.A1(n_1423),
.A2(n_138),
.B1(n_139),
.B2(n_141),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1421),
.Y(n_1442)
);

NOR2xp67_ASAP7_75t_L g1443 ( 
.A(n_1414),
.B(n_142),
.Y(n_1443)
);

NAND3xp33_ASAP7_75t_L g1444 ( 
.A(n_1423),
.B(n_144),
.C(n_145),
.Y(n_1444)
);

AND4x1_ASAP7_75t_L g1445 ( 
.A(n_1407),
.B(n_152),
.C(n_153),
.D(n_155),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1424),
.Y(n_1446)
);

NOR3xp33_ASAP7_75t_L g1447 ( 
.A(n_1419),
.B(n_156),
.C(n_158),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1413),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1433),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1415),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1416),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1434),
.Y(n_1452)
);

NOR2x1_ASAP7_75t_L g1453 ( 
.A(n_1422),
.B(n_165),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1425),
.A2(n_166),
.B1(n_169),
.B2(n_170),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1446),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1449),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1439),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1439),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1446),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1437),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1436),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1448),
.A2(n_1425),
.B1(n_1417),
.B2(n_1429),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1450),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1442),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1452),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1443),
.B(n_1431),
.Y(n_1466)
);

INVxp67_ASAP7_75t_SL g1467 ( 
.A(n_1453),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1441),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1441),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1440),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1451),
.Y(n_1471)
);

OAI22x1_ASAP7_75t_L g1472 ( 
.A1(n_1455),
.A2(n_1454),
.B1(n_1435),
.B2(n_1445),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1456),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1456),
.A2(n_1438),
.B1(n_1444),
.B2(n_1430),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1465),
.Y(n_1475)
);

AO22x2_ASAP7_75t_L g1476 ( 
.A1(n_1457),
.A2(n_1447),
.B1(n_1428),
.B2(n_1432),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1457),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1467),
.A2(n_1426),
.B1(n_1427),
.B2(n_185),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1459),
.B(n_171),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1459),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1461),
.A2(n_194),
.B1(n_195),
.B2(n_201),
.Y(n_1481)
);

OAI22x1_ASAP7_75t_L g1482 ( 
.A1(n_1463),
.A2(n_1471),
.B1(n_1470),
.B2(n_1462),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1473),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1479),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1477),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1476),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1475),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1476),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1485),
.A2(n_1480),
.B1(n_1460),
.B2(n_1458),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1485),
.A2(n_1482),
.B1(n_1472),
.B2(n_1470),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1483),
.A2(n_1464),
.B1(n_1478),
.B2(n_1474),
.Y(n_1491)
);

OAI22xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1488),
.A2(n_1464),
.B1(n_1466),
.B2(n_1468),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1490),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1489),
.Y(n_1494)
);

AO22x2_ASAP7_75t_L g1495 ( 
.A1(n_1493),
.A2(n_1486),
.B1(n_1491),
.B2(n_1484),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1495),
.Y(n_1496)
);

AOI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1496),
.A2(n_1492),
.B1(n_1464),
.B2(n_1494),
.C(n_1487),
.Y(n_1497)
);

AOI211xp5_ASAP7_75t_L g1498 ( 
.A1(n_1497),
.A2(n_1469),
.B(n_1468),
.C(n_1481),
.Y(n_1498)
);


endmodule