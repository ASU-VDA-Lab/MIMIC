module real_jpeg_4479_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_1),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_1),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_89)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_1),
.A2(n_124),
.B1(n_155),
.B2(n_159),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_1),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_1),
.A2(n_65),
.B1(n_94),
.B2(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_2),
.A2(n_62),
.B1(n_65),
.B2(n_67),
.Y(n_61)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_2),
.A2(n_45),
.B1(n_67),
.B2(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_4),
.Y(n_137)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_5),
.Y(n_173)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_5),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_5),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_5),
.B(n_9),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_6),
.A2(n_77),
.B1(n_80),
.B2(n_81),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_6),
.A2(n_80),
.B1(n_167),
.B2(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_7),
.Y(n_101)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_7),
.Y(n_117)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_8),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_9),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_9),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_9),
.A2(n_57),
.B1(n_91),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_9),
.A2(n_57),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_9),
.A2(n_57),
.B1(n_77),
.B2(n_185),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_9),
.A2(n_227),
.B(n_228),
.C(n_232),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_9),
.B(n_22),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_9),
.B(n_263),
.C(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_9),
.B(n_153),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_9),
.B(n_148),
.C(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_9),
.B(n_96),
.Y(n_300)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_10),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_10),
.Y(n_93)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_10),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_11),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_211),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_210),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_189),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_15),
.B(n_189),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_162),
.C(n_175),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_16),
.B(n_162),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_87),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_17),
.B(n_88),
.C(n_161),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_60),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_18),
.A2(n_60),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_18),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_18),
.A2(n_223),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_19),
.A2(n_20),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_47),
.B1(n_52),
.B2(n_59),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_21),
.B(n_52),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_21),
.A2(n_47),
.B1(n_52),
.B2(n_59),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_21),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_21),
.A2(n_52),
.B(n_59),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_34),
.Y(n_21)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_28),
.B2(n_32),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_38),
.Y(n_202)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_39),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_39),
.Y(n_140)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_40),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_40),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_57),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_59),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_60),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_68),
.B1(n_75),
.B2(n_83),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_61),
.A2(n_180),
.B(n_183),
.Y(n_179)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_64),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_64),
.Y(n_266)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_68),
.B(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_69),
.B(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_69),
.A2(n_184),
.B1(n_235),
.B2(n_238),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_69),
.A2(n_184),
.B1(n_235),
.B2(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_74),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_76),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_77),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_121),
.B1(n_160),
.B2(n_161),
.Y(n_87)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_88),
.B(n_203),
.C(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_88),
.A2(n_160),
.B1(n_203),
.B2(n_301),
.Y(n_326)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_95),
.B1(n_118),
.B2(n_120),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_89),
.A2(n_95),
.B1(n_118),
.B2(n_120),
.Y(n_188)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_93),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_95),
.A2(n_118),
.B(n_120),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_108),
.Y(n_95)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_102),
.B2(n_105),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_99),
.Y(n_227)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_101),
.Y(n_229)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_113),
.B2(n_115),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_121),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_121),
.A2(n_161),
.B1(n_177),
.B2(n_178),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_121),
.B(n_177),
.C(n_280),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_121),
.A2(n_161),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_121),
.B(n_219),
.C(n_312),
.Y(n_330)
);

AO22x2_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_128),
.B1(n_153),
.B2(n_154),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_122),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

INVx6_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_129),
.B(n_130),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_129),
.A2(n_130),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_145),
.Y(n_129)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

AOI22x1_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_133),
.B1(n_138),
.B2(n_141),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g283 ( 
.A(n_147),
.Y(n_283)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_170),
.B2(n_174),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_170),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_168),
.B(n_169),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_168),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_170),
.A2(n_174),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_171),
.B(n_184),
.Y(n_286)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_186),
.C(n_188),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_177),
.A2(n_178),
.B1(n_259),
.B2(n_267),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_177),
.B(n_267),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_179),
.Y(n_328)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_188),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_188),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_188),
.A2(n_219),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_208),
.B2(n_209),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_197),
.B1(n_198),
.B2(n_207),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_203),
.B(n_206),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_203),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_203),
.A2(n_297),
.B1(n_298),
.B2(n_301),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_203),
.Y(n_301)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_208),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_239),
.B(n_338),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_214),
.B(n_216),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.C(n_224),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_217),
.B(n_221),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_223),
.B(n_234),
.C(n_273),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_223),
.B(n_293),
.C(n_295),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_224),
.B(n_322),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_225),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_233),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_226),
.A2(n_233),
.B1(n_234),
.B2(n_318),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_226),
.Y(n_318)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_234),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_234),
.B(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_254),
.Y(n_255)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_320),
.B(n_336),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_305),
.B(n_319),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_290),
.B(n_304),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_277),
.B(n_289),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_269),
.B(n_276),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_256),
.B(n_268),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_253),
.B(n_255),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_251),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_251),
.A2(n_257),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_258),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_257),
.B(n_299),
.C(n_301),
.Y(n_315)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_275),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_275),
.Y(n_276)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_279),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_288),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_286),
.B2(n_287),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_287),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_303),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_303),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_295),
.B1(n_296),
.B2(n_302),
.Y(n_291)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_307),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_315),
.C(n_316),
.Y(n_332)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_323),
.B(n_331),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_323),
.C(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.C(n_329),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_334),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_327),
.A2(n_329),
.B1(n_330),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);


endmodule