module fake_netlist_6_1008_n_803 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_803);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_803;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_758;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_631;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_608;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_508;
wire n_361;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g159 ( 
.A(n_42),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_35),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_130),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_1),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_13),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_146),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_11),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_95),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_8),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_38),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g172 ( 
.A(n_12),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_92),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_15),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_46),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_18),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_12),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_124),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_114),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_97),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_51),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_82),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_73),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_30),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_70),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_54),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_58),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_3),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_27),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_74),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_85),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_101),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_87),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_44),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_53),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_111),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_147),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_27),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_6),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_136),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_14),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_90),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_49),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_102),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_104),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_2),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_141),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_110),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_167),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g221 ( 
.A(n_162),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_163),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_199),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_164),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_207),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_168),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_173),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_0),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_175),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_180),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_181),
.B(n_0),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_182),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_183),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_159),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_214),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_185),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_160),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_160),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_181),
.B(n_1),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_161),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_171),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_172),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_186),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_161),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_172),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_189),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_172),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_L g258 ( 
.A(n_164),
.B(n_2),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_178),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_179),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_184),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_227),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_176),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_226),
.B(n_176),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_195),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_232),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_233),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_235),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_222),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_218),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_229),
.B(n_176),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_218),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_236),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_238),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_239),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_259),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_234),
.B(n_166),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_242),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_237),
.B(n_166),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_221),
.B(n_213),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_213),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_247),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_248),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_248),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_250),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_250),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_240),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_246),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_253),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_223),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_225),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_230),
.B(n_215),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_256),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_230),
.B(n_215),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_219),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_231),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_245),
.Y(n_310)
);

NAND2xp33_ASAP7_75t_SL g311 ( 
.A(n_245),
.B(n_206),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_231),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_271),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_285),
.Y(n_314)
);

NAND2xp33_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_188),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

INVx4_ASAP7_75t_SL g318 ( 
.A(n_289),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_294),
.B(n_188),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_265),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_267),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_241),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_263),
.Y(n_324)
);

AND2x2_ASAP7_75t_SL g325 ( 
.A(n_287),
.B(n_188),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

AND2x2_ASAP7_75t_SL g327 ( 
.A(n_287),
.B(n_188),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_285),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_274),
.Y(n_329)
);

BUFx4f_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_294),
.B(n_241),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_270),
.B(n_194),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_252),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_263),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_266),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_263),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_266),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_294),
.B(n_187),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_272),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_269),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_269),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_269),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_278),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_286),
.B(n_255),
.Y(n_347)
);

AO22x2_ASAP7_75t_L g348 ( 
.A1(n_303),
.A2(n_203),
.B1(n_210),
.B2(n_196),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_278),
.Y(n_349)
);

NAND3x1_ASAP7_75t_L g350 ( 
.A(n_295),
.B(n_190),
.C(n_201),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_276),
.Y(n_351)
);

NAND2x1p5_ASAP7_75t_L g352 ( 
.A(n_293),
.B(n_205),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_285),
.B(n_257),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_278),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_295),
.B(n_216),
.Y(n_355)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_276),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_277),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_281),
.B(n_198),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_277),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_277),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_262),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_282),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_281),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_290),
.B(n_200),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_262),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_281),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_264),
.B(n_202),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_293),
.B(n_204),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_293),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_290),
.A2(n_212),
.B1(n_211),
.B2(n_208),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_291),
.A2(n_307),
.B1(n_305),
.B2(n_279),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_292),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_264),
.B(n_28),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_292),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_293),
.B(n_206),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_303),
.B(n_3),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_279),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_291),
.B(n_29),
.Y(n_378)
);

NAND3xp33_ASAP7_75t_SL g379 ( 
.A(n_375),
.B(n_311),
.C(n_280),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_372),
.B(n_296),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_296),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_297),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_334),
.B(n_305),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_334),
.B(n_307),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_331),
.B(n_297),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_325),
.B(n_308),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_325),
.B(n_308),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_301),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_313),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_336),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_327),
.A2(n_301),
.B1(n_302),
.B2(n_309),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_330),
.A2(n_302),
.B(n_312),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_347),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_327),
.B(n_377),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_309),
.Y(n_397)
);

O2A1O1Ixp5_ASAP7_75t_L g398 ( 
.A1(n_340),
.A2(n_312),
.B(n_268),
.C(n_304),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_304),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_373),
.B(n_275),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_373),
.A2(n_310),
.B1(n_275),
.B2(n_280),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_317),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_356),
.A2(n_378),
.B1(n_328),
.B2(n_321),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_364),
.B(n_283),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_320),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_SL g408 ( 
.A(n_369),
.B(n_310),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_318),
.B(n_283),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_318),
.B(n_300),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_318),
.B(n_306),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_353),
.B(n_31),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_330),
.A2(n_299),
.B(n_298),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_353),
.B(n_333),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_323),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_361),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_371),
.B(n_323),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_322),
.B(n_326),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_336),
.Y(n_419)
);

O2A1O1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_340),
.A2(n_315),
.B(n_368),
.C(n_319),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_330),
.A2(n_284),
.B(n_273),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_316),
.B(n_347),
.Y(n_422)
);

NAND2xp33_ASAP7_75t_L g423 ( 
.A(n_352),
.B(n_345),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_336),
.Y(n_424)
);

NAND2xp33_ASAP7_75t_L g425 ( 
.A(n_352),
.B(n_32),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_369),
.B(n_33),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_369),
.B(n_34),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_365),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_329),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_328),
.B(n_349),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_367),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_365),
.Y(n_432)
);

NOR2x1p5_ASAP7_75t_L g433 ( 
.A(n_376),
.B(n_4),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_368),
.B(n_4),
.Y(n_435)
);

AND2x4_ASAP7_75t_SL g436 ( 
.A(n_367),
.B(n_36),
.Y(n_436)
);

NOR2x1p5_ASAP7_75t_L g437 ( 
.A(n_341),
.B(n_5),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_354),
.B(n_37),
.Y(n_438)
);

NOR3x1_ASAP7_75t_L g439 ( 
.A(n_375),
.B(n_319),
.C(n_350),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_355),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_338),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_338),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_343),
.A2(n_346),
.B1(n_351),
.B2(n_359),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_343),
.B(n_39),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_343),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_339),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_339),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_314),
.B(n_40),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_383),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_R g450 ( 
.A(n_389),
.B(n_341),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_415),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_413),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_384),
.B(n_314),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_314),
.Y(n_455)
);

NAND2x1_ASAP7_75t_L g456 ( 
.A(n_394),
.B(n_400),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_399),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_381),
.B(n_357),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_381),
.B(n_360),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_416),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_428),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_406),
.B(n_362),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_390),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_390),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_428),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_R g468 ( 
.A(n_379),
.B(n_362),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_422),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_421),
.Y(n_470)
);

AO221x1_ASAP7_75t_L g471 ( 
.A1(n_404),
.A2(n_348),
.B1(n_350),
.B2(n_343),
.C(n_346),
.Y(n_471)
);

INVx5_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_382),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_397),
.B(n_363),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

BUFx8_ASAP7_75t_L g476 ( 
.A(n_382),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_432),
.Y(n_477)
);

BUFx12f_ASAP7_75t_SL g478 ( 
.A(n_382),
.Y(n_478)
);

CKINVDCx8_ASAP7_75t_R g479 ( 
.A(n_385),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_431),
.B(n_367),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_385),
.B(n_370),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_397),
.B(n_342),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_401),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_400),
.B(n_342),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_380),
.B(n_344),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_396),
.B(n_344),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_436),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_392),
.B(n_358),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_441),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_441),
.Y(n_490)
);

A2O1A1Ixp33_ASAP7_75t_L g491 ( 
.A1(n_435),
.A2(n_358),
.B(n_332),
.C(n_366),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_434),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_388),
.B(n_366),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_388),
.A2(n_351),
.B1(n_346),
.B2(n_315),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_390),
.Y(n_496)
);

NAND3xp33_ASAP7_75t_SL g497 ( 
.A(n_403),
.B(n_348),
.C(n_335),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_429),
.Y(n_498)
);

BUFx4f_ASAP7_75t_L g499 ( 
.A(n_436),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_434),
.B(n_346),
.Y(n_500)
);

AND3x1_ASAP7_75t_SL g501 ( 
.A(n_437),
.B(n_348),
.C(n_8),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_442),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_395),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_442),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_472),
.B(n_412),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_481),
.A2(n_455),
.B(n_454),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_427),
.B(n_426),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_484),
.A2(n_448),
.B(n_438),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_386),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_469),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_449),
.B(n_386),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_472),
.A2(n_423),
.B(n_424),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_465),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_464),
.B(n_402),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_486),
.A2(n_430),
.B(n_420),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_472),
.A2(n_423),
.B(n_424),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_472),
.A2(n_424),
.B(n_419),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_455),
.A2(n_387),
.B(n_405),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_449),
.A2(n_391),
.B1(n_387),
.B2(n_402),
.Y(n_519)
);

AOI21x1_ASAP7_75t_L g520 ( 
.A1(n_493),
.A2(n_408),
.B(n_446),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_473),
.B(n_418),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_484),
.A2(n_445),
.B(n_447),
.Y(n_522)
);

AOI211x1_ASAP7_75t_L g523 ( 
.A1(n_497),
.A2(n_444),
.B(n_409),
.C(n_410),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_488),
.A2(n_395),
.B(n_425),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_456),
.A2(n_395),
.B(n_425),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_483),
.B(n_435),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_503),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_454),
.A2(n_395),
.B(n_443),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_503),
.A2(n_445),
.B(n_444),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_458),
.B(n_433),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_489),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_459),
.B(n_418),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_476),
.Y(n_533)
);

A2O1A1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_459),
.A2(n_440),
.B(n_398),
.C(n_418),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_461),
.B(n_439),
.Y(n_535)
);

O2A1O1Ixp5_ASAP7_75t_L g536 ( 
.A1(n_491),
.A2(n_440),
.B(n_447),
.C(n_446),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_476),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_486),
.A2(n_411),
.B(n_337),
.Y(n_538)
);

AOI221x1_ASAP7_75t_L g539 ( 
.A1(n_474),
.A2(n_351),
.B1(n_337),
.B2(n_335),
.C(n_324),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_451),
.B(n_351),
.Y(n_540)
);

OA21x2_ASAP7_75t_L g541 ( 
.A1(n_482),
.A2(n_324),
.B(n_83),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_461),
.B(n_7),
.Y(n_542)
);

AO31x2_ASAP7_75t_L g543 ( 
.A1(n_482),
.A2(n_9),
.A3(n_10),
.B(n_11),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_487),
.B(n_9),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_474),
.A2(n_84),
.B(n_156),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_485),
.B(n_495),
.Y(n_546)
);

OA22x2_ASAP7_75t_L g547 ( 
.A1(n_471),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_485),
.A2(n_89),
.B(n_154),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_503),
.A2(n_86),
.B(n_152),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_531),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_510),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_527),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_531),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_532),
.B(n_452),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_535),
.A2(n_499),
.B1(n_470),
.B2(n_453),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_514),
.B(n_457),
.Y(n_556)
);

AO21x2_ASAP7_75t_L g557 ( 
.A1(n_520),
.A2(n_494),
.B(n_477),
.Y(n_557)
);

O2A1O1Ixp33_ASAP7_75t_SL g558 ( 
.A1(n_534),
.A2(n_460),
.B(n_462),
.C(n_463),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_533),
.Y(n_559)
);

OA21x2_ASAP7_75t_L g560 ( 
.A1(n_539),
.A2(n_467),
.B(n_502),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_522),
.A2(n_504),
.B(n_490),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_509),
.A2(n_480),
.B1(n_499),
.B2(n_492),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_521),
.B(n_492),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_540),
.Y(n_564)
);

NAND3xp33_ASAP7_75t_L g565 ( 
.A(n_526),
.B(n_480),
.C(n_498),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_547),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_536),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_521),
.Y(n_568)
);

OAI21x1_ASAP7_75t_L g569 ( 
.A1(n_524),
.A2(n_536),
.B(n_525),
.Y(n_569)
);

NAND2x1p5_ASAP7_75t_L g570 ( 
.A(n_527),
.B(n_492),
.Y(n_570)
);

O2A1O1Ixp33_ASAP7_75t_SL g571 ( 
.A1(n_534),
.A2(n_496),
.B(n_475),
.C(n_501),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_547),
.Y(n_572)
);

AO31x2_ASAP7_75t_L g573 ( 
.A1(n_519),
.A2(n_466),
.A3(n_465),
.B(n_500),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_515),
.A2(n_496),
.B(n_475),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_533),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_509),
.A2(n_478),
.B1(n_468),
.B2(n_500),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_521),
.Y(n_577)
);

OAI21x1_ASAP7_75t_L g578 ( 
.A1(n_515),
.A2(n_503),
.B(n_466),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_546),
.B(n_450),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_530),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_508),
.A2(n_81),
.B(n_151),
.Y(n_581)
);

NOR2x1_ASAP7_75t_L g582 ( 
.A(n_513),
.B(n_41),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_512),
.A2(n_91),
.B(n_150),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_527),
.Y(n_584)
);

CKINVDCx8_ASAP7_75t_R g585 ( 
.A(n_527),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_513),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_542),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_537),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_511),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_516),
.A2(n_80),
.B(n_149),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_543),
.Y(n_591)
);

OAI21x1_ASAP7_75t_L g592 ( 
.A1(n_528),
.A2(n_79),
.B(n_148),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_589),
.B(n_506),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_SL g594 ( 
.A(n_579),
.B(n_548),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_564),
.B(n_544),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_585),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_553),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_576),
.A2(n_523),
.B1(n_518),
.B2(n_537),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_587),
.B(n_538),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_592),
.B(n_505),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_550),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_556),
.B(n_543),
.Y(n_602)
);

NAND2x1_ASAP7_75t_L g603 ( 
.A(n_582),
.B(n_529),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_555),
.A2(n_505),
.B1(n_549),
.B2(n_541),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_565),
.A2(n_541),
.B1(n_545),
.B2(n_517),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_592),
.B(n_545),
.Y(n_606)
);

BUFx4_ASAP7_75t_R g607 ( 
.A(n_588),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_550),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_556),
.B(n_543),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_558),
.A2(n_541),
.B(n_507),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_563),
.B(n_543),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_554),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_566),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_554),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_572),
.B(n_158),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_560),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_568),
.B(n_19),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_568),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_618)
);

O2A1O1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_571),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_552),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_577),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g622 ( 
.A1(n_569),
.A2(n_23),
.B(n_24),
.Y(n_622)
);

OAI221xp5_ASAP7_75t_L g623 ( 
.A1(n_580),
.A2(n_25),
.B1(n_26),
.B2(n_43),
.C(n_45),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_577),
.B(n_99),
.Y(n_624)
);

A2O1A1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_567),
.A2(n_25),
.B(n_26),
.C(n_47),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_563),
.B(n_48),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_562),
.B(n_50),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_585),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_591),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_586),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_586),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_563),
.B(n_567),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_551),
.B(n_52),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_551),
.B(n_571),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_586),
.B(n_145),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_573),
.B(n_55),
.Y(n_636)
);

OAI22xp33_ASAP7_75t_L g637 ( 
.A1(n_559),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_560),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_586),
.B(n_60),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_559),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_588),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_601),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_623),
.A2(n_575),
.B1(n_557),
.B2(n_583),
.Y(n_643)
);

OAI222xp33_ASAP7_75t_L g644 ( 
.A1(n_618),
.A2(n_575),
.B1(n_570),
.B2(n_558),
.C1(n_573),
.C2(n_590),
.Y(n_644)
);

AOI222xp33_ASAP7_75t_L g645 ( 
.A1(n_613),
.A2(n_590),
.B1(n_583),
.B2(n_584),
.C1(n_552),
.C2(n_581),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_594),
.A2(n_557),
.B1(n_552),
.B2(n_584),
.Y(n_646)
);

OAI211xp5_ASAP7_75t_L g647 ( 
.A1(n_621),
.A2(n_581),
.B(n_584),
.C(n_552),
.Y(n_647)
);

INVx5_ASAP7_75t_SL g648 ( 
.A(n_600),
.Y(n_648)
);

AOI211xp5_ASAP7_75t_L g649 ( 
.A1(n_637),
.A2(n_584),
.B(n_574),
.C(n_578),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_629),
.Y(n_650)
);

AOI221xp5_ASAP7_75t_L g651 ( 
.A1(n_619),
.A2(n_557),
.B1(n_570),
.B2(n_573),
.C(n_561),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_594),
.A2(n_560),
.B1(n_574),
.B2(n_578),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_612),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_593),
.B(n_573),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_598),
.A2(n_561),
.B1(n_65),
.B2(n_67),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_601),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_610),
.A2(n_64),
.B(n_68),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_627),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_627),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_611),
.B(n_78),
.Y(n_660)
);

OAI22xp33_ASAP7_75t_L g661 ( 
.A1(n_640),
.A2(n_595),
.B1(n_599),
.B2(n_628),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_597),
.Y(n_662)
);

OA21x2_ASAP7_75t_L g663 ( 
.A1(n_622),
.A2(n_93),
.B(n_94),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_628),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_634),
.A2(n_96),
.B1(n_98),
.B2(n_100),
.Y(n_665)
);

AND2x2_ASAP7_75t_SL g666 ( 
.A(n_636),
.B(n_607),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_593),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_615),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_602),
.B(n_112),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_614),
.B(n_115),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_617),
.B(n_116),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_609),
.B(n_144),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_616),
.Y(n_673)
);

AOI221xp5_ASAP7_75t_SL g674 ( 
.A1(n_625),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.C(n_120),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_615),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_675)
);

AOI221xp5_ASAP7_75t_L g676 ( 
.A1(n_625),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.C(n_128),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_607),
.Y(n_677)
);

OR2x6_ASAP7_75t_L g678 ( 
.A(n_600),
.B(n_129),
.Y(n_678)
);

OAI211xp5_ASAP7_75t_SL g679 ( 
.A1(n_633),
.A2(n_132),
.B(n_134),
.C(n_135),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_654),
.B(n_616),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_676),
.A2(n_636),
.B1(n_640),
.B2(n_641),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_673),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_650),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_642),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_662),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_653),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_678),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_648),
.B(n_638),
.Y(n_688)
);

INVxp67_ASAP7_75t_SL g689 ( 
.A(n_642),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_656),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_648),
.B(n_606),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_648),
.B(n_606),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_656),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_648),
.B(n_606),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_678),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_652),
.B(n_606),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_646),
.B(n_600),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_677),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_663),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_678),
.B(n_600),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_651),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_678),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_664),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_663),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_677),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_669),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_683),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_687),
.B(n_666),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_703),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_683),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_687),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_681),
.A2(n_666),
.B1(n_677),
.B2(n_659),
.Y(n_712)
);

AND2x2_ASAP7_75t_SL g713 ( 
.A(n_687),
.B(n_701),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_701),
.B(n_674),
.C(n_671),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_688),
.B(n_700),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_703),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_688),
.B(n_663),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_683),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_707),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_711),
.B(n_680),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_716),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_715),
.B(n_706),
.Y(n_722)
);

OAI21xp33_ASAP7_75t_L g723 ( 
.A1(n_714),
.A2(n_681),
.B(n_706),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_709),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_715),
.B(n_700),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_711),
.B(n_713),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_713),
.B(n_717),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_722),
.B(n_717),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_720),
.B(n_710),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_723),
.B(n_686),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_719),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_726),
.B(n_686),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_719),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_731),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_730),
.B(n_727),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_732),
.B(n_727),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_728),
.B(n_725),
.Y(n_737)
);

AND4x1_ASAP7_75t_L g738 ( 
.A(n_733),
.B(n_649),
.C(n_702),
.D(n_695),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_SL g739 ( 
.A1(n_735),
.A2(n_712),
.B1(n_721),
.B2(n_687),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_734),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_737),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_735),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_741),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_742),
.B(n_736),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_R g745 ( 
.A(n_743),
.B(n_741),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_744),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_SL g747 ( 
.A(n_743),
.B(n_739),
.Y(n_747)
);

NAND4xp25_ASAP7_75t_L g748 ( 
.A(n_746),
.B(n_740),
.C(n_708),
.D(n_664),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_747),
.B(n_729),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_745),
.Y(n_750)
);

NOR3x1_ASAP7_75t_L g751 ( 
.A(n_746),
.B(n_703),
.C(n_738),
.Y(n_751)
);

NOR3xp33_ASAP7_75t_SL g752 ( 
.A(n_745),
.B(n_661),
.C(n_721),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_745),
.B(n_671),
.C(n_658),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_SL g754 ( 
.A(n_752),
.B(n_675),
.C(n_668),
.Y(n_754)
);

OAI211xp5_ASAP7_75t_L g755 ( 
.A1(n_750),
.A2(n_667),
.B(n_655),
.C(n_643),
.Y(n_755)
);

AND4x1_ASAP7_75t_L g756 ( 
.A(n_753),
.B(n_626),
.C(n_657),
.D(n_702),
.Y(n_756)
);

NAND4xp75_ASAP7_75t_L g757 ( 
.A(n_751),
.B(n_660),
.C(n_670),
.D(n_626),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_749),
.A2(n_687),
.B1(n_724),
.B2(n_698),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_748),
.A2(n_665),
.B(n_679),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_750),
.A2(n_699),
.B(n_635),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_757),
.B(n_725),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_754),
.A2(n_687),
.B1(n_695),
.B2(n_698),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_758),
.A2(n_687),
.B1(n_698),
.B2(n_705),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_756),
.Y(n_764)
);

AOI221xp5_ASAP7_75t_L g765 ( 
.A1(n_760),
.A2(n_704),
.B1(n_699),
.B2(n_644),
.C(n_647),
.Y(n_765)
);

AOI21xp33_ASAP7_75t_SL g766 ( 
.A1(n_755),
.A2(n_596),
.B(n_669),
.Y(n_766)
);

OAI21xp33_ASAP7_75t_L g767 ( 
.A1(n_759),
.A2(n_705),
.B(n_700),
.Y(n_767)
);

AOI221x1_ASAP7_75t_L g768 ( 
.A1(n_758),
.A2(n_639),
.B1(n_596),
.B2(n_624),
.C(n_631),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_764),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_767),
.A2(n_705),
.B1(n_709),
.B2(n_704),
.Y(n_770)
);

NOR3xp33_ASAP7_75t_L g771 ( 
.A(n_766),
.B(n_596),
.C(n_672),
.Y(n_771)
);

XNOR2xp5_ASAP7_75t_L g772 ( 
.A(n_762),
.B(n_660),
.Y(n_772)
);

O2A1O1Ixp5_ASAP7_75t_L g773 ( 
.A1(n_763),
.A2(n_704),
.B(n_699),
.C(n_603),
.Y(n_773)
);

NOR2xp67_ASAP7_75t_SL g774 ( 
.A(n_761),
.B(n_624),
.Y(n_774)
);

AOI322xp5_ASAP7_75t_L g775 ( 
.A1(n_765),
.A2(n_704),
.A3(n_696),
.B1(n_697),
.B2(n_716),
.C1(n_604),
.C2(n_694),
.Y(n_775)
);

AOI222xp33_ASAP7_75t_L g776 ( 
.A1(n_768),
.A2(n_704),
.B1(n_696),
.B2(n_697),
.C1(n_685),
.C2(n_605),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_764),
.B(n_696),
.Y(n_777)
);

AOI32xp33_ASAP7_75t_L g778 ( 
.A1(n_769),
.A2(n_620),
.A3(n_697),
.B1(n_672),
.B2(n_694),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_777),
.B(n_685),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_SL g780 ( 
.A(n_771),
.B(n_645),
.C(n_620),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_SL g781 ( 
.A(n_775),
.B(n_620),
.C(n_692),
.Y(n_781)
);

XOR2xp5_ASAP7_75t_L g782 ( 
.A(n_772),
.B(n_140),
.Y(n_782)
);

OAI222xp33_ASAP7_75t_L g783 ( 
.A1(n_774),
.A2(n_692),
.B1(n_691),
.B2(n_630),
.C1(n_694),
.C2(n_710),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_SL g784 ( 
.A(n_776),
.B(n_691),
.C(n_692),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_770),
.A2(n_718),
.B1(n_707),
.B2(n_688),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_773),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_L g787 ( 
.A(n_786),
.B(n_718),
.C(n_691),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_782),
.A2(n_785),
.B1(n_778),
.B2(n_779),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_779),
.B(n_693),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_781),
.Y(n_790)
);

CKINVDCx16_ASAP7_75t_R g791 ( 
.A(n_784),
.Y(n_791)
);

OAI221xp5_ASAP7_75t_L g792 ( 
.A1(n_780),
.A2(n_783),
.B1(n_680),
.B2(n_689),
.C(n_690),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_782),
.Y(n_793)
);

INVx1_ASAP7_75t_SL g794 ( 
.A(n_793),
.Y(n_794)
);

AO22x2_ASAP7_75t_L g795 ( 
.A1(n_790),
.A2(n_693),
.B1(n_690),
.B2(n_684),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_791),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_796),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_797),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_798),
.A2(n_794),
.B1(n_787),
.B2(n_788),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_799),
.A2(n_798),
.B1(n_792),
.B2(n_795),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_800),
.B(n_789),
.Y(n_801)
);

OAI221xp5_ASAP7_75t_L g802 ( 
.A1(n_801),
.A2(n_142),
.B1(n_143),
.B2(n_608),
.C(n_689),
.Y(n_802)
);

AOI211xp5_ASAP7_75t_L g803 ( 
.A1(n_802),
.A2(n_684),
.B(n_682),
.C(n_632),
.Y(n_803)
);


endmodule