module fake_netlist_1_5532_n_520 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_520);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_520;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g73 ( .A(n_27), .Y(n_73) );
BUFx3_ASAP7_75t_L g74 ( .A(n_42), .Y(n_74) );
CKINVDCx20_ASAP7_75t_R g75 ( .A(n_51), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_41), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_69), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_44), .Y(n_78) );
BUFx6f_ASAP7_75t_L g79 ( .A(n_43), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_59), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_13), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_11), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_53), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_32), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_62), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_64), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_72), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_26), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_28), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_35), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_66), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_15), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_1), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_14), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_10), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_2), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_25), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_3), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_47), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_34), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_61), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_58), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_12), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_52), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_7), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_87), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_76), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_87), .Y(n_108) );
AND2x4_ASAP7_75t_L g109 ( .A(n_94), .B(n_82), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_76), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_79), .Y(n_111) );
INVx3_ASAP7_75t_L g112 ( .A(n_94), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_92), .B(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_80), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_79), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_83), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_82), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_93), .B(n_0), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_83), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_84), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_98), .B(n_1), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_84), .Y(n_123) );
NAND2xp33_ASAP7_75t_SL g124 ( .A(n_90), .B(n_2), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_79), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_73), .B(n_3), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_85), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_85), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_109), .B(n_98), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_118), .B(n_91), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_109), .B(n_103), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_107), .B(n_97), .Y(n_132) );
INVx4_ASAP7_75t_L g133 ( .A(n_122), .Y(n_133) );
AO22x2_ASAP7_75t_L g134 ( .A1(n_122), .A2(n_86), .B1(n_99), .B2(n_102), .Y(n_134) );
INVx4_ASAP7_75t_L g135 ( .A(n_122), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_122), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_107), .B(n_86), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_106), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_112), .Y(n_139) );
INVx4_ASAP7_75t_L g140 ( .A(n_109), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_106), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_110), .B(n_99), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_109), .B(n_103), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_112), .B(n_105), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g146 ( .A(n_110), .B(n_101), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_108), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_112), .B(n_95), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_114), .B(n_102), .Y(n_149) );
BUFx2_ASAP7_75t_L g150 ( .A(n_126), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_114), .B(n_96), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_111), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_115), .B(n_117), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_115), .B(n_101), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_133), .B(n_126), .Y(n_155) );
INVx5_ASAP7_75t_L g156 ( .A(n_153), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_146), .B(n_117), .Y(n_157) );
BUFx4f_ASAP7_75t_L g158 ( .A(n_153), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_139), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_150), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_146), .B(n_128), .Y(n_161) );
INVx2_ASAP7_75t_SL g162 ( .A(n_153), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_139), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
NAND3xp33_ASAP7_75t_L g167 ( .A(n_133), .B(n_128), .C(n_127), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
INVxp67_ASAP7_75t_L g169 ( .A(n_150), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_131), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_133), .B(n_135), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_146), .B(n_120), .Y(n_172) );
AOI21xp33_ASAP7_75t_L g173 ( .A1(n_134), .A2(n_127), .B(n_120), .Y(n_173) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_134), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
CKINVDCx6p67_ASAP7_75t_R g179 ( .A(n_153), .Y(n_179) );
CKINVDCx11_ASAP7_75t_R g180 ( .A(n_131), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_135), .B(n_78), .Y(n_181) );
BUFx12f_ASAP7_75t_SL g182 ( .A(n_140), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_135), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_140), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_129), .B(n_121), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_154), .B(n_121), .Y(n_187) );
NAND3xp33_ASAP7_75t_L g188 ( .A(n_173), .B(n_130), .C(n_140), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_179), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_157), .B(n_154), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_175), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_163), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_176), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_174), .A2(n_134), .B1(n_154), .B2(n_151), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_176), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_186), .B(n_134), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_175), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_163), .Y(n_198) );
INVx1_ASAP7_75t_SL g199 ( .A(n_180), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_157), .B(n_154), .Y(n_201) );
BUFx2_ASAP7_75t_L g202 ( .A(n_182), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_173), .A2(n_134), .B1(n_151), .B2(n_131), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_186), .B(n_151), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_179), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_176), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_177), .Y(n_207) );
INVxp67_ASAP7_75t_SL g208 ( .A(n_164), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_178), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_156), .B(n_140), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_161), .A2(n_142), .B1(n_149), .B2(n_137), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_164), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_178), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_177), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_182), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_178), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_186), .B(n_151), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_184), .Y(n_218) );
NAND3xp33_ASAP7_75t_L g219 ( .A(n_167), .B(n_155), .C(n_161), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_164), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g221 ( .A1(n_199), .A2(n_170), .B1(n_169), .B2(n_160), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_194), .A2(n_172), .B1(n_187), .B2(n_186), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_219), .A2(n_167), .B(n_172), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_SL g224 ( .A1(n_211), .A2(n_137), .B(n_142), .C(n_149), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_218), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_218), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_192), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_196), .A2(n_182), .B1(n_185), .B2(n_184), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_211), .A2(n_187), .B(n_132), .C(n_113), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_192), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_199), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_205), .B(n_175), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_190), .A2(n_171), .B(n_181), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_198), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_198), .Y(n_235) );
OAI21xp33_ASAP7_75t_SL g236 ( .A1(n_194), .A2(n_132), .B(n_159), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_207), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_196), .A2(n_185), .B1(n_184), .B2(n_124), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_193), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_207), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_193), .Y(n_241) );
OR2x6_ASAP7_75t_L g242 ( .A(n_196), .B(n_164), .Y(n_242) );
NOR2xp33_ASAP7_75t_R g243 ( .A(n_202), .B(n_75), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_193), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_204), .B(n_175), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_222), .A2(n_203), .B1(n_190), .B2(n_201), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_225), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_225), .B(n_204), .Y(n_248) );
INVx4_ASAP7_75t_L g249 ( .A(n_242), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_226), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_221), .A2(n_204), .B1(n_217), .B2(n_203), .Y(n_251) );
NOR2xp67_ASAP7_75t_L g252 ( .A(n_226), .B(n_205), .Y(n_252) );
OAI21xp33_ASAP7_75t_L g253 ( .A1(n_238), .A2(n_188), .B(n_217), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_239), .B(n_217), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_239), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_241), .B(n_201), .Y(n_256) );
BUFx12f_ASAP7_75t_L g257 ( .A(n_242), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_241), .B(n_216), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_229), .A2(n_188), .B1(n_205), .B2(n_77), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_244), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_236), .A2(n_81), .B1(n_219), .B2(n_100), .Y(n_261) );
OAI221xp5_ASAP7_75t_L g262 ( .A1(n_231), .A2(n_119), .B1(n_215), .B2(n_202), .C(n_123), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_227), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_232), .Y(n_264) );
AOI21xp33_ASAP7_75t_L g265 ( .A1(n_232), .A2(n_215), .B(n_214), .Y(n_265) );
NAND2xp33_ASAP7_75t_R g266 ( .A(n_256), .B(n_243), .Y(n_266) );
BUFx2_ASAP7_75t_L g267 ( .A(n_249), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_256), .B(n_244), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_261), .A2(n_228), .B1(n_234), .B2(n_240), .Y(n_269) );
AOI221xp5_ASAP7_75t_L g270 ( .A1(n_262), .A2(n_224), .B1(n_129), .B2(n_245), .C(n_131), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_263), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_261), .A2(n_242), .B1(n_227), .B2(n_240), .Y(n_272) );
INVx8_ASAP7_75t_L g273 ( .A(n_257), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_247), .B(n_230), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_248), .B(n_245), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_263), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_258), .B(n_230), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_255), .A2(n_237), .B(n_235), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_255), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_247), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_246), .A2(n_237), .B1(n_235), .B2(n_234), .Y(n_281) );
OAI21x1_ASAP7_75t_L g282 ( .A1(n_260), .A2(n_223), .B(n_233), .Y(n_282) );
NAND4xp25_ASAP7_75t_SL g283 ( .A(n_251), .B(n_123), .C(n_138), .D(n_141), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_250), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_260), .A2(n_206), .B(n_195), .Y(n_285) );
AOI222xp33_ASAP7_75t_L g286 ( .A1(n_248), .A2(n_143), .B1(n_148), .B2(n_144), .C1(n_214), .C2(n_147), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_259), .A2(n_242), .B1(n_205), .B2(n_189), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_283), .A2(n_257), .B1(n_253), .B2(n_249), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_271), .B(n_249), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_279), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_271), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_276), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_276), .B(n_250), .Y(n_293) );
AOI211xp5_ASAP7_75t_L g294 ( .A1(n_272), .A2(n_265), .B(n_143), .C(n_104), .Y(n_294) );
OAI322xp33_ASAP7_75t_L g295 ( .A1(n_266), .A2(n_284), .A3(n_280), .B1(n_274), .B2(n_275), .C1(n_254), .C2(n_141), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_282), .A2(n_252), .B(n_258), .Y(n_296) );
INVxp67_ASAP7_75t_R g297 ( .A(n_277), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_280), .B(n_254), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_268), .B(n_264), .Y(n_299) );
AO22x1_ASAP7_75t_L g300 ( .A1(n_267), .A2(n_264), .B1(n_232), .B2(n_78), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_284), .B(n_264), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_268), .B(n_264), .Y(n_302) );
INVxp67_ASAP7_75t_L g303 ( .A(n_277), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_279), .B(n_264), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_279), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_278), .B(n_252), .Y(n_306) );
NAND3xp33_ASAP7_75t_L g307 ( .A(n_270), .B(n_79), .C(n_74), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_274), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_278), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_269), .A2(n_232), .B1(n_216), .B2(n_195), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_282), .Y(n_311) );
NOR3xp33_ASAP7_75t_SL g312 ( .A(n_287), .B(n_88), .C(n_138), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_285), .Y(n_313) );
AOI331xp33_ASAP7_75t_L g314 ( .A1(n_281), .A2(n_145), .A3(n_147), .B1(n_6), .B2(n_7), .B3(n_8), .C1(n_9), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_286), .B(n_79), .C(n_74), .Y(n_315) );
OAI33xp33_ASAP7_75t_L g316 ( .A1(n_286), .A2(n_145), .A3(n_88), .B1(n_6), .B2(n_8), .B3(n_9), .Y(n_316) );
AO21x2_ASAP7_75t_L g317 ( .A1(n_285), .A2(n_144), .B(n_148), .Y(n_317) );
OAI221xp5_ASAP7_75t_L g318 ( .A1(n_267), .A2(n_89), .B1(n_197), .B2(n_191), .C(n_168), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_273), .A2(n_148), .B1(n_144), .B2(n_143), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_273), .B(n_89), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_320), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_303), .B(n_273), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_308), .B(n_273), .Y(n_323) );
OAI33xp33_ASAP7_75t_L g324 ( .A1(n_291), .A2(n_4), .A3(n_5), .B1(n_10), .B2(n_11), .B3(n_12), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_290), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_293), .Y(n_326) );
NAND3xp33_ASAP7_75t_L g327 ( .A(n_300), .B(n_111), .C(n_116), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_293), .B(n_291), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_292), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_292), .B(n_273), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_306), .B(n_111), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_299), .B(n_111), .Y(n_332) );
NAND4xp25_ASAP7_75t_L g333 ( .A(n_294), .B(n_148), .C(n_144), .D(n_143), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_306), .B(n_111), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_299), .B(n_116), .Y(n_335) );
INVxp67_ASAP7_75t_L g336 ( .A(n_320), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_301), .B(n_4), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_293), .Y(n_338) );
NOR3xp33_ASAP7_75t_L g339 ( .A(n_316), .B(n_197), .C(n_191), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_298), .B(n_5), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_295), .A2(n_197), .B(n_191), .C(n_159), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_302), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_290), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_302), .B(n_116), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_305), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_304), .Y(n_346) );
OAI31xp33_ASAP7_75t_L g347 ( .A1(n_315), .A2(n_189), .A3(n_159), .B(n_168), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_298), .B(n_13), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_304), .B(n_116), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_301), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_297), .B(n_116), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_314), .B(n_289), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_297), .B(n_125), .Y(n_353) );
BUFx3_ASAP7_75t_L g354 ( .A(n_289), .Y(n_354) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_312), .A2(n_189), .B(n_158), .C(n_195), .Y(n_355) );
OAI221xp5_ASAP7_75t_L g356 ( .A1(n_288), .A2(n_125), .B1(n_197), .B2(n_166), .C(n_168), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_305), .B(n_125), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_307), .A2(n_213), .B(n_206), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_289), .B(n_14), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_309), .Y(n_360) );
NAND3xp33_ASAP7_75t_L g361 ( .A(n_300), .B(n_125), .C(n_213), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_309), .B(n_15), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_310), .B(n_16), .Y(n_363) );
OAI31xp33_ASAP7_75t_SL g364 ( .A1(n_318), .A2(n_16), .A3(n_17), .B(n_18), .Y(n_364) );
OAI221xp5_ASAP7_75t_L g365 ( .A1(n_319), .A2(n_125), .B1(n_165), .B2(n_166), .C(n_191), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_313), .B(n_17), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_313), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_329), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_350), .B(n_311), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_328), .B(n_311), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_338), .B(n_317), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_326), .B(n_317), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_346), .B(n_296), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_360), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_366), .B(n_317), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_360), .Y(n_376) );
OAI211xp5_ASAP7_75t_SL g377 ( .A1(n_352), .A2(n_152), .B(n_18), .C(n_191), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_342), .B(n_332), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_321), .B(n_296), .Y(n_379) );
NOR2xp67_ASAP7_75t_L g380 ( .A(n_361), .B(n_327), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_354), .B(n_213), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_331), .Y(n_382) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_330), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_362), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_366), .B(n_209), .Y(n_385) );
INVx1_ASAP7_75t_SL g386 ( .A(n_330), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_332), .B(n_209), .Y(n_387) );
XNOR2xp5_ASAP7_75t_L g388 ( .A(n_323), .B(n_19), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_351), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_354), .B(n_209), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_362), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_325), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_352), .B(n_20), .Y(n_393) );
NAND2xp33_ASAP7_75t_SL g394 ( .A(n_337), .B(n_205), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_335), .B(n_21), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_331), .B(n_220), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_337), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_336), .B(n_206), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_331), .B(n_220), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_335), .Y(n_400) );
NOR4xp25_ASAP7_75t_L g401 ( .A(n_340), .B(n_166), .C(n_165), .D(n_152), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_359), .A2(n_165), .B1(n_208), .B2(n_185), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_344), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_344), .B(n_22), .Y(n_404) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_334), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_325), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g407 ( .A1(n_355), .A2(n_208), .B(n_158), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_348), .B(n_23), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_322), .B(n_24), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_334), .B(n_322), .Y(n_410) );
OAI21xp33_ASAP7_75t_L g411 ( .A1(n_364), .A2(n_152), .B(n_30), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_343), .B(n_29), .Y(n_412) );
NOR2x1_ASAP7_75t_L g413 ( .A(n_351), .B(n_220), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_349), .B(n_31), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_343), .B(n_33), .Y(n_415) );
INVx1_ASAP7_75t_SL g416 ( .A(n_353), .Y(n_416) );
NAND2x2_ASAP7_75t_L g417 ( .A(n_363), .B(n_36), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_349), .B(n_37), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_386), .B(n_345), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_377), .A2(n_393), .B1(n_394), .B2(n_411), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_378), .B(n_334), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_368), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_393), .A2(n_324), .B1(n_333), .B2(n_339), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_383), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_397), .B(n_367), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_378), .B(n_345), .Y(n_426) );
CKINVDCx16_ASAP7_75t_R g427 ( .A(n_388), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_381), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_384), .B(n_349), .Y(n_429) );
OAI21xp33_ASAP7_75t_L g430 ( .A1(n_401), .A2(n_353), .B(n_355), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_391), .B(n_357), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_369), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_410), .B(n_357), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_370), .Y(n_434) );
NAND2xp33_ASAP7_75t_SL g435 ( .A(n_382), .B(n_358), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_389), .B(n_356), .Y(n_436) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_394), .A2(n_347), .B(n_341), .C(n_365), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_405), .B(n_38), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_372), .B(n_152), .C(n_212), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_374), .Y(n_440) );
NAND3xp33_ASAP7_75t_L g441 ( .A(n_371), .B(n_220), .C(n_212), .Y(n_441) );
XNOR2xp5_ASAP7_75t_L g442 ( .A(n_400), .B(n_403), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_373), .B(n_39), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_376), .Y(n_444) );
XOR2x2_ASAP7_75t_L g445 ( .A(n_409), .B(n_40), .Y(n_445) );
NOR3xp33_ASAP7_75t_SL g446 ( .A(n_409), .B(n_210), .C(n_46), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_375), .B(n_45), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_373), .B(n_48), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_390), .Y(n_449) );
OAI33xp33_ASAP7_75t_L g450 ( .A1(n_408), .A2(n_49), .A3(n_50), .B1(n_54), .B2(n_55), .B3(n_56), .Y(n_450) );
AOI32xp33_ASAP7_75t_L g451 ( .A1(n_416), .A2(n_183), .A3(n_60), .B1(n_63), .B2(n_65), .Y(n_451) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_379), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_392), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_392), .B(n_57), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_406), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_406), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_413), .B(n_67), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_385), .B(n_68), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_380), .A2(n_158), .B(n_153), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_398), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_417), .A2(n_153), .B1(n_183), .B2(n_220), .Y(n_461) );
OAI22xp33_ASAP7_75t_L g462 ( .A1(n_417), .A2(n_179), .B1(n_212), .B2(n_220), .Y(n_462) );
NAND2x1_ASAP7_75t_L g463 ( .A(n_412), .B(n_220), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_387), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_396), .A2(n_158), .B(n_212), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_395), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g467 ( .A(n_396), .B(n_212), .C(n_200), .Y(n_467) );
AOI31xp33_ASAP7_75t_L g468 ( .A1(n_399), .A2(n_395), .A3(n_407), .B(n_402), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_399), .B(n_70), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_412), .B(n_71), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_404), .A2(n_183), .B1(n_200), .B2(n_212), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_414), .A2(n_200), .B(n_212), .C(n_183), .Y(n_472) );
OAI211xp5_ASAP7_75t_L g473 ( .A1(n_418), .A2(n_200), .B(n_156), .C(n_164), .Y(n_473) );
OAI21xp33_ASAP7_75t_L g474 ( .A1(n_415), .A2(n_200), .B(n_162), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_368), .Y(n_475) );
NOR2x1_ASAP7_75t_SL g476 ( .A(n_396), .B(n_200), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_397), .B(n_162), .Y(n_477) );
INVx2_ASAP7_75t_SL g478 ( .A(n_378), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_368), .Y(n_479) );
NAND3xp33_ASAP7_75t_L g480 ( .A(n_393), .B(n_156), .C(n_162), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_368), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_368), .Y(n_482) );
NAND2xp33_ASAP7_75t_L g483 ( .A(n_411), .B(n_156), .Y(n_483) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_468), .A2(n_434), .B1(n_452), .B2(n_432), .C(n_424), .Y(n_484) );
AOI211xp5_ASAP7_75t_L g485 ( .A1(n_462), .A2(n_436), .B(n_483), .C(n_430), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_427), .Y(n_486) );
NAND2xp33_ASAP7_75t_SL g487 ( .A(n_466), .B(n_442), .Y(n_487) );
NAND3xp33_ASAP7_75t_SL g488 ( .A(n_420), .B(n_451), .C(n_423), .Y(n_488) );
NAND4xp75_ASAP7_75t_L g489 ( .A(n_420), .B(n_423), .C(n_461), .D(n_446), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_482), .Y(n_490) );
OAI21xp33_ASAP7_75t_L g491 ( .A1(n_478), .A2(n_421), .B(n_429), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_449), .B(n_428), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_445), .A2(n_464), .B1(n_435), .B2(n_450), .Y(n_493) );
OAI32xp33_ASAP7_75t_L g494 ( .A1(n_430), .A2(n_426), .A3(n_419), .B1(n_448), .B2(n_475), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_460), .B(n_479), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_481), .Y(n_496) );
OAI321xp33_ASAP7_75t_L g497 ( .A1(n_462), .A2(n_431), .A3(n_459), .B1(n_437), .B2(n_447), .C(n_425), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_453), .Y(n_498) );
AOI31xp33_ASAP7_75t_L g499 ( .A1(n_480), .A2(n_438), .A3(n_443), .B(n_457), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_498), .Y(n_500) );
NAND3xp33_ASAP7_75t_SL g501 ( .A(n_493), .B(n_473), .C(n_465), .Y(n_501) );
AOI211xp5_ASAP7_75t_L g502 ( .A1(n_488), .A2(n_443), .B(n_438), .C(n_422), .Y(n_502) );
OAI21xp5_ASAP7_75t_SL g503 ( .A1(n_493), .A2(n_470), .B(n_473), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_490), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_494), .A2(n_472), .B(n_458), .C(n_469), .Y(n_505) );
AOI211xp5_ASAP7_75t_L g506 ( .A1(n_497), .A2(n_439), .B(n_474), .C(n_472), .Y(n_506) );
OAI31xp33_ASAP7_75t_L g507 ( .A1(n_487), .A2(n_453), .A3(n_467), .B(n_433), .Y(n_507) );
NAND5xp2_ASAP7_75t_L g508 ( .A(n_503), .B(n_485), .C(n_484), .D(n_489), .E(n_491), .Y(n_508) );
OAI221xp5_ASAP7_75t_L g509 ( .A1(n_507), .A2(n_486), .B1(n_499), .B2(n_496), .C(n_492), .Y(n_509) );
OAI22x1_ASAP7_75t_L g510 ( .A1(n_504), .A2(n_498), .B1(n_495), .B2(n_471), .Y(n_510) );
NAND3xp33_ASAP7_75t_SL g511 ( .A(n_502), .B(n_463), .C(n_454), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_509), .B(n_501), .C(n_505), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_510), .Y(n_513) );
AOI221x1_ASAP7_75t_L g514 ( .A1(n_508), .A2(n_500), .B1(n_505), .B2(n_477), .C(n_440), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_513), .Y(n_515) );
AOI211xp5_ASAP7_75t_L g516 ( .A1(n_512), .A2(n_511), .B(n_506), .C(n_441), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_515), .A2(n_514), .B(n_476), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_517), .Y(n_518) );
BUFx2_ASAP7_75t_L g519 ( .A(n_518), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g520 ( .A1(n_519), .A2(n_516), .B1(n_456), .B2(n_455), .C(n_444), .Y(n_520) );
endmodule