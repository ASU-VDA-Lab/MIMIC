module fake_jpeg_24507_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_1),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_29),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_44),
.Y(n_60)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_30),
.B1(n_26),
.B2(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_18),
.B(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_46),
.B(n_32),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_47),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_20),
.C(n_24),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_22),
.C(n_19),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_59),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_34),
.B1(n_30),
.B2(n_20),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_70),
.B1(n_20),
.B2(n_24),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_66),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_30),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_71),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_37),
.B(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_27),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_25),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_34),
.B1(n_43),
.B2(n_42),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_83),
.B1(n_86),
.B2(n_88),
.Y(n_116)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_80),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_92),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_85),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_24),
.B1(n_45),
.B2(n_29),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_26),
.B1(n_22),
.B2(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_93),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_77),
.B(n_75),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_38),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_25),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_68),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_73),
.B(n_11),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

HAxp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_28),
.CON(n_110),
.SN(n_110)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_120),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_69),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_58),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_92),
.B(n_15),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_115),
.B(n_14),
.Y(n_137)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_75),
.A2(n_68),
.A3(n_49),
.B1(n_50),
.B2(n_55),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_83),
.A2(n_49),
.B1(n_55),
.B2(n_63),
.Y(n_119)
);

AO22x1_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_48),
.B1(n_57),
.B2(n_78),
.Y(n_131)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_126),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_90),
.C(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_137),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_80),
.B(n_91),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_107),
.B(n_106),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_131),
.A2(n_57),
.B1(n_58),
.B2(n_103),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_91),
.C(n_68),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_69),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_139),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_95),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_103),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_147),
.B1(n_151),
.B2(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_146),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_152),
.Y(n_161)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

OAI22x1_ASAP7_75t_SL g147 ( 
.A1(n_126),
.A2(n_116),
.B1(n_99),
.B2(n_101),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_127),
.B(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_154),
.A2(n_133),
.B1(n_122),
.B2(n_114),
.Y(n_167)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_155),
.B(n_157),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_120),
.B(n_116),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_125),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_104),
.A3(n_100),
.B1(n_108),
.B2(n_120),
.C1(n_105),
.C2(n_101),
.Y(n_157)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_124),
.Y(n_158)
);

AOI321xp33_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_149),
.A3(n_141),
.B1(n_154),
.B2(n_146),
.C(n_131),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_125),
.A3(n_129),
.B1(n_121),
.B2(n_136),
.C1(n_135),
.C2(n_100),
.Y(n_162)
);

AOI31xp33_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_156),
.A3(n_145),
.B(n_153),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_48),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_144),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_123),
.C(n_133),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_170),
.C(n_61),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_132),
.C(n_115),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_171),
.A2(n_174),
.B(n_168),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_149),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_177),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_131),
.B(n_61),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_160),
.B(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_179),
.B(n_180),
.Y(n_181)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_166),
.B(n_163),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_185),
.B(n_14),
.Y(n_191)
);

AOI221xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_87),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_169),
.B1(n_161),
.B2(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_177),
.C(n_179),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_190),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_184),
.A2(n_178),
.B1(n_174),
.B2(n_172),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_192),
.B(n_1),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g193 ( 
.A1(n_189),
.A2(n_181),
.A3(n_186),
.B1(n_87),
.B2(n_4),
.C1(n_5),
.C2(n_1),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_196),
.C(n_2),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_192),
.A2(n_2),
.B(n_3),
.Y(n_196)
);

AO21x2_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_6),
.B(n_7),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_3),
.C(n_5),
.Y(n_199)
);

AOI221xp5_ASAP7_75t_L g201 ( 
.A1(n_199),
.A2(n_6),
.B1(n_8),
.B2(n_198),
.C(n_196),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_201),
.Y(n_202)
);


endmodule