module fake_jpeg_3170_n_104 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_43),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_38),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_48),
.B1(n_40),
.B2(n_29),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_33),
.B1(n_37),
.B2(n_34),
.Y(n_48)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_40),
.B1(n_51),
.B2(n_52),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_60),
.B1(n_62),
.B2(n_2),
.Y(n_73)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_32),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_33),
.B1(n_38),
.B2(n_31),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_46),
.B(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_72),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_66),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_71),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_1),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_3),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_3),
.B(n_4),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_6),
.B(n_11),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_4),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_79),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_82),
.Y(n_85)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_87),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_17),
.C(n_25),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_90),
.C(n_91),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_19),
.C(n_9),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_12),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_94),
.C(n_85),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_93),
.B(n_88),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_89),
.B1(n_95),
.B2(n_74),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

AOI31xp67_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_76),
.A3(n_16),
.B(n_20),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_15),
.B1(n_21),
.B2(n_23),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_24),
.Y(n_104)
);


endmodule