module fake_netlist_1_8094_n_14 (n_1, n_2, n_0, n_14);
input n_1;
input n_2;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
AND2x4_ASAP7_75t_L g3 ( .A(n_0), .B(n_1), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_1), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_6) );
OAI21x1_ASAP7_75t_L g7 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_6), .B(n_3), .Y(n_9) );
AOI21xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_8), .B(n_6), .Y(n_10) );
OR2x2_ASAP7_75t_L g11 ( .A(n_9), .B(n_3), .Y(n_11) );
OAI211xp5_ASAP7_75t_SL g12 ( .A1(n_11), .A2(n_8), .B(n_2), .C(n_9), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
AOI22xp33_ASAP7_75t_SL g14 ( .A1(n_13), .A2(n_2), .B1(n_10), .B2(n_9), .Y(n_14) );
endmodule