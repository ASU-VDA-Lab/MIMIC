module real_jpeg_5544_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_249;
wire n_288;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_295;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx8_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_1),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_1),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_1),
.B(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_2),
.Y(n_114)
);

NAND2x1p5_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_3),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_3),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_3),
.B(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_3),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_3),
.B(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_3),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_4),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_5),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_5),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_5),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_5),
.B(n_79),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_5),
.B(n_129),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_5),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_5),
.B(n_215),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_5),
.B(n_254),
.Y(n_253)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_7),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_7),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_7),
.Y(n_199)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_7),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_8),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_8),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_8),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_8),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_8),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_9),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_9),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_9),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_9),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_9),
.B(n_49),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_10),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_10),
.B(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_11),
.Y(n_173)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_13),
.Y(n_109)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_13),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_14),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_14),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_14),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_14),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_14),
.B(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_14),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_14),
.B(n_79),
.Y(n_257)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_15),
.Y(n_215)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_16),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_16),
.B(n_40),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_16),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_16),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_17),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_17),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_17),
.B(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_183),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_182),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_153),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_22),
.B(n_153),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_92),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_61),
.C(n_72),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_24),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_43),
.C(n_50),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_25),
.A2(n_26),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_27),
.B(n_33),
.C(n_42),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_28),
.B(n_246),
.Y(n_245)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_31),
.Y(n_234)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_31),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_37),
.B2(n_42),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_44),
.B(n_51),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_45),
.B(n_48),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_47),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_49),
.Y(n_129)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJx2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.C(n_58),
.Y(n_51)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_52),
.B(n_54),
.CI(n_58),
.CON(n_270),
.SN(n_270)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_57),
.Y(n_219)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_57),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_57),
.Y(n_255)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_61),
.B(n_72),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_67),
.C(n_70),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_82),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_74),
.B(n_78),
.C(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_82),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.C(n_90),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_83),
.B(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_86),
.A2(n_90),
.B1(n_91),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_86),
.Y(n_178)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_88),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_89),
.Y(n_246)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_120),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_111),
.Y(n_119)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_113),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_140),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_135),
.C(n_139),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_122),
.A2(n_123),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_128),
.C(n_150),
.Y(n_149)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_133),
.Y(n_193)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_136),
.B(n_138),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_139),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_143),
.B1(n_151),
.B2(n_152),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_149),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_179),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_155),
.B(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_157),
.B(n_179),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_174),
.C(n_175),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_158),
.B(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_166),
.C(n_171),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_159),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_160),
.A2(n_161),
.B1(n_164),
.B2(n_165),
.Y(n_247)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_167),
.B(n_172),
.Y(n_267)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_174),
.Y(n_287)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

AOI21x1_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_291),
.B(n_295),
.Y(n_183)
);

OAI21x1_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_278),
.B(n_290),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_263),
.B(n_277),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_238),
.B(n_262),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_221),
.B(n_237),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_201),
.B(n_220),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_197),
.B(n_200),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_195),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_194),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_203),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_211),
.B2(n_212),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_214),
.C(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_208),
.Y(n_229)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_236),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_236),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_230),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_229),
.C(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_227),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_230),
.Y(n_296)
);

FAx1_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.CI(n_235),
.CON(n_230),
.SN(n_230)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_250),
.C(n_251),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_241),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_249),
.C(n_252),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_245),
.C(n_247),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_258),
.C(n_260),
.Y(n_275)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_257),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_258),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_276),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_276),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_268),
.C(n_289),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_273),
.C(n_274),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_270),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_288),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_288),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_285),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_282),
.C(n_285),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_292),
.B(n_294),
.Y(n_295)
);


endmodule