module fake_jpeg_12198_n_446 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_446);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_446;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_41),
.Y(n_47)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_47),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_27),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_53),
.Y(n_103)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_70),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_23),
.Y(n_70)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx4f_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_27),
.B(n_16),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_91),
.Y(n_93)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_0),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_17),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_82),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_0),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_89),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_90),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_41),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_46),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_109),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_21),
.B1(n_18),
.B2(n_32),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_97),
.A2(n_100),
.B1(n_135),
.B2(n_137),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_37),
.B1(n_45),
.B2(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_34),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_104),
.B(n_115),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_63),
.A2(n_46),
.B1(n_21),
.B2(n_37),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_105),
.A2(n_117),
.B1(n_119),
.B2(n_25),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_21),
.C(n_32),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_86),
.B1(n_66),
.B2(n_78),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_45),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_52),
.A2(n_44),
.B1(n_43),
.B2(n_42),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_54),
.A2(n_34),
.B1(n_33),
.B2(n_20),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_47),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_123),
.B(n_130),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_38),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_59),
.A2(n_44),
.B1(n_43),
.B2(n_42),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_71),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_87),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_58),
.A2(n_38),
.B1(n_43),
.B2(n_42),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_62),
.A2(n_44),
.B1(n_39),
.B2(n_28),
.Y(n_137)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_148),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_92),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_149),
.B(n_165),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_150),
.B(n_168),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_151),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_83),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_152),
.B(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_105),
.A2(n_68),
.B1(n_65),
.B2(n_88),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_158),
.A2(n_180),
.B1(n_181),
.B2(n_186),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_69),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_159),
.B(n_161),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_103),
.B(n_75),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_87),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_162),
.Y(n_215)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_39),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_164),
.B(n_184),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_39),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_166),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_124),
.A2(n_134),
.B(n_97),
.C(n_106),
.Y(n_167)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_125),
.A3(n_139),
.B1(n_145),
.B2(n_122),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_95),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_67),
.B1(n_74),
.B2(n_72),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_SL g204 ( 
.A1(n_169),
.A2(n_141),
.B(n_107),
.C(n_110),
.Y(n_204)
);

HAxp5_ASAP7_75t_SL g170 ( 
.A(n_143),
.B(n_60),
.CON(n_170),
.SN(n_170)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_118),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_172),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_80),
.B1(n_28),
.B2(n_25),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_173),
.A2(n_128),
.B1(n_145),
.B2(n_122),
.Y(n_202)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_106),
.B(n_25),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_141),
.C(n_7),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_28),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_177),
.B(n_178),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_24),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_133),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_24),
.B1(n_142),
.B2(n_114),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_0),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_182),
.B(n_192),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_98),
.B(n_2),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_98),
.Y(n_185)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_142),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_3),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_5),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_191),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_242)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_193),
.Y(n_235)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_194),
.Y(n_211)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_197),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_118),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_114),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_10),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_201),
.B(n_169),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_202),
.A2(n_210),
.B1(n_228),
.B2(n_190),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_204),
.A2(n_229),
.B1(n_152),
.B2(n_173),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_165),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_195),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_147),
.A2(n_125),
.B(n_141),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_207),
.B(n_214),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_150),
.A2(n_107),
.B1(n_129),
.B2(n_110),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_177),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_176),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_171),
.A2(n_129),
.B1(n_146),
.B2(n_8),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_157),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_160),
.A2(n_146),
.B1(n_7),
.B2(n_8),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_190),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_147),
.B(n_6),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_233),
.C(n_241),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_147),
.B(n_6),
.C(n_8),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_237),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_149),
.B(n_162),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_182),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_244),
.B(n_245),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_218),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_246),
.B(n_252),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_187),
.B1(n_171),
.B2(n_178),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_247),
.A2(n_251),
.B1(n_259),
.B2(n_264),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_248),
.A2(n_254),
.B1(n_258),
.B2(n_263),
.Y(n_289)
);

AO21x1_ASAP7_75t_L g312 ( 
.A1(n_249),
.A2(n_253),
.B(n_257),
.Y(n_312)
);

OAI32xp33_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_167),
.A3(n_187),
.B1(n_162),
.B2(n_179),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_261),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_176),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_216),
.A2(n_169),
.B1(n_174),
.B2(n_193),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_255),
.Y(n_310)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_210),
.A2(n_154),
.B1(n_156),
.B2(n_185),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_215),
.A2(n_169),
.B1(n_148),
.B2(n_185),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_192),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_269),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_225),
.B(n_153),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_262),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_216),
.A2(n_194),
.B1(n_196),
.B2(n_155),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_215),
.A2(n_191),
.B1(n_183),
.B2(n_166),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_229),
.A2(n_175),
.B1(n_170),
.B2(n_168),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_265),
.A2(n_272),
.B1(n_277),
.B2(n_243),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_227),
.B(n_163),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_270),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_216),
.A2(n_172),
.B1(n_197),
.B2(n_14),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_267),
.A2(n_275),
.B(n_266),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_241),
.B(n_11),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_226),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_213),
.B(n_12),
.Y(n_273)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_211),
.Y(n_275)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_212),
.Y(n_276)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_203),
.A2(n_12),
.B1(n_15),
.B2(n_220),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_221),
.B(n_230),
.Y(n_278)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_231),
.B(n_207),
.C(n_233),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_279),
.B(n_269),
.C(n_283),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_230),
.B(n_201),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_280),
.A2(n_247),
.B(n_253),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_223),
.B(n_214),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_274),
.Y(n_290)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_223),
.B(n_200),
.C(n_206),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_200),
.C(n_206),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_257),
.A2(n_224),
.B(n_204),
.Y(n_284)
);

OAI21xp33_ASAP7_75t_SL g327 ( 
.A1(n_284),
.A2(n_295),
.B(n_316),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_287),
.B(n_288),
.C(n_292),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_204),
.C(n_235),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_290),
.B(n_297),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_204),
.C(n_211),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_248),
.A2(n_204),
.B1(n_202),
.B2(n_217),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_293),
.A2(n_294),
.B1(n_298),
.B2(n_306),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_257),
.A2(n_212),
.B(n_199),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_199),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_304),
.C(n_313),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_254),
.A2(n_217),
.B1(n_208),
.B2(n_236),
.Y(n_298)
);

AO22x1_ASAP7_75t_L g299 ( 
.A1(n_249),
.A2(n_209),
.B1(n_232),
.B2(n_208),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_299),
.B(n_311),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_245),
.B(n_279),
.C(n_281),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_280),
.A2(n_217),
.B1(n_236),
.B2(n_240),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_260),
.A2(n_240),
.B1(n_209),
.B2(n_232),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_307),
.A2(n_318),
.B1(n_310),
.B2(n_289),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_252),
.B(n_244),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_255),
.Y(n_314)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_314),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_270),
.A2(n_261),
.B(n_250),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_315),
.B(n_311),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_265),
.C(n_256),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_293),
.A2(n_259),
.B1(n_275),
.B2(n_264),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_319),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_262),
.Y(n_320)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_320),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_282),
.Y(n_321)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_268),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_322),
.B(n_324),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_323),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_276),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_285),
.A2(n_277),
.B1(n_251),
.B2(n_263),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_328),
.A2(n_338),
.B1(n_347),
.B2(n_304),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_330),
.Y(n_350)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_314),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_331),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_345),
.C(n_286),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_300),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_335),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_307),
.Y(n_335)
);

HAxp5_ASAP7_75t_SL g336 ( 
.A(n_316),
.B(n_267),
.CON(n_336),
.SN(n_336)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_336),
.B(n_340),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_285),
.A2(n_276),
.B1(n_292),
.B2(n_312),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_339),
.A2(n_337),
.B(n_343),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_301),
.B(n_313),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_287),
.B(n_306),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_341),
.B(n_343),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_329),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_291),
.B(n_315),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_346),
.Y(n_358)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_296),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_312),
.A2(n_288),
.B1(n_284),
.B2(n_299),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_349),
.A2(n_353),
.B1(n_359),
.B2(n_365),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_328),
.A2(n_299),
.B1(n_317),
.B2(n_309),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_321),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_329),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_338),
.A2(n_309),
.B1(n_305),
.B2(n_290),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_335),
.A2(n_323),
.B1(n_332),
.B2(n_337),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_361),
.A2(n_366),
.B1(n_368),
.B2(n_330),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_331),
.C(n_344),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_364),
.A2(n_365),
.B(n_355),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_347),
.A2(n_301),
.B1(n_295),
.B2(n_286),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_327),
.A2(n_341),
.B1(n_333),
.B2(n_320),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_334),
.A2(n_323),
.B1(n_332),
.B2(n_339),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_345),
.B(n_325),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_370),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_325),
.B(n_326),
.Y(n_370)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_371),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_367),
.B(n_326),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_372),
.B(n_378),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_342),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_379),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_357),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_376),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_358),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_346),
.Y(n_380)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_380),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_358),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_385),
.Y(n_397)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_363),
.Y(n_382)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_382),
.Y(n_401)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_383),
.Y(n_398)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_363),
.Y(n_384)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_384),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_360),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_330),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_391),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_388),
.A2(n_348),
.B1(n_356),
.B2(n_351),
.Y(n_395)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_389),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_354),
.B(n_350),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_390),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_385),
.A2(n_368),
.B1(n_349),
.B2(n_361),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_394),
.A2(n_405),
.B1(n_386),
.B2(n_373),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_395),
.A2(n_359),
.B1(n_373),
.B2(n_381),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_389),
.A2(n_353),
.B1(n_356),
.B2(n_351),
.Y(n_405)
);

BUFx24_ASAP7_75t_SL g406 ( 
.A(n_391),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_406),
.B(n_374),
.Y(n_412)
);

AOI21x1_ASAP7_75t_L g408 ( 
.A1(n_400),
.A2(n_364),
.B(n_355),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_409),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_387),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_379),
.C(n_377),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_410),
.B(n_413),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_411),
.A2(n_352),
.B1(n_398),
.B2(n_404),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_412),
.B(n_402),
.Y(n_420)
);

OAI21x1_ASAP7_75t_SL g413 ( 
.A1(n_397),
.A2(n_390),
.B(n_376),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_395),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_415),
.Y(n_428)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_392),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_416),
.B(n_418),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_402),
.A2(n_386),
.B1(n_407),
.B2(n_403),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_417),
.A2(n_407),
.B(n_371),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_377),
.C(n_362),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_397),
.B(n_366),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_419),
.B(n_401),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_384),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_422),
.A2(n_414),
.B(n_417),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_423),
.B(n_424),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_418),
.B(n_382),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_425),
.B(n_410),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_429),
.B(n_431),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_422),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_427),
.B(n_419),
.C(n_409),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_432),
.B(n_434),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_396),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_433),
.B(n_421),
.C(n_426),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_435),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_436),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_440),
.A2(n_437),
.B(n_438),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_441),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_439),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_443),
.A2(n_442),
.B1(n_398),
.B2(n_426),
.Y(n_444)
);

AOI221xp5_ASAP7_75t_L g445 ( 
.A1(n_444),
.A2(n_423),
.B1(n_352),
.B2(n_396),
.C(n_383),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_375),
.Y(n_446)
);


endmodule