module fake_jpeg_27679_n_273 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_38;
wire n_26;
wire n_28;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_33),
.Y(n_48)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_38),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_23),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_42),
.B(n_19),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_26),
.B1(n_32),
.B2(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_24),
.B1(n_32),
.B2(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_26),
.B1(n_24),
.B2(n_32),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_26),
.B1(n_19),
.B2(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_33),
.A2(n_19),
.B1(n_18),
.B2(n_27),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_16),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_30),
.B1(n_29),
.B2(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_29),
.B1(n_16),
.B2(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_25),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_36),
.Y(n_63)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_63),
.B(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_58),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_68),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_73),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_37),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_89),
.C(n_37),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_18),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_23),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_54),
.B(n_29),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_22),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_34),
.B1(n_39),
.B2(n_37),
.Y(n_87)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_41),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_37),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_103),
.Y(n_123)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g137 ( 
.A(n_96),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_98),
.Y(n_128)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_112),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_64),
.B(n_37),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_88),
.B(n_87),
.Y(n_136)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_61),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_15),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_0),
.Y(n_141)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_116),
.B(n_118),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_86),
.B1(n_74),
.B2(n_83),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_119),
.B1(n_125),
.B2(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_69),
.B1(n_89),
.B2(n_67),
.Y(n_119)
);

AOI22x1_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_81),
.B1(n_87),
.B2(n_71),
.Y(n_120)
);

OA21x2_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_121),
.B(n_87),
.Y(n_152)
);

AO21x1_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_81),
.B(n_87),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_130),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_136),
.B(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_63),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_124),
.B(n_127),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_65),
.B1(n_68),
.B2(n_82),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_80),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_132),
.Y(n_163)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_103),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_71),
.B1(n_61),
.B2(n_78),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_45),
.B1(n_34),
.B2(n_48),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_79),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_85),
.B1(n_70),
.B2(n_75),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_84),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_21),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_94),
.B(n_21),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_141),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_145),
.A2(n_20),
.B(n_16),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_120),
.A2(n_111),
.B1(n_95),
.B2(n_99),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_146),
.A2(n_152),
.B1(n_59),
.B2(n_20),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_110),
.B1(n_99),
.B2(n_111),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_148),
.A2(n_149),
.B1(n_164),
.B2(n_48),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_109),
.B1(n_77),
.B2(n_108),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_77),
.C(n_97),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_166),
.C(n_167),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_159),
.B1(n_118),
.B2(n_128),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_107),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_1),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_168),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_72),
.B(n_108),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_171),
.B(n_90),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_136),
.B1(n_121),
.B2(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_97),
.B1(n_96),
.B2(n_104),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_107),
.C(n_113),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_113),
.C(n_37),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_104),
.B(n_96),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_112),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_90),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_145),
.B(n_132),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_176),
.B(n_158),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_177),
.Y(n_208)
);

HAxp5_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_134),
.CON(n_176),
.SN(n_176)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_185),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_182),
.B1(n_189),
.B2(n_168),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_146),
.A2(n_62),
.B1(n_112),
.B2(n_59),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_190),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_152),
.A2(n_34),
.B1(n_76),
.B2(n_90),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_152),
.Y(n_209)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_194),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_28),
.C(n_2),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_156),
.C(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_144),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_197),
.A2(n_210),
.B1(n_189),
.B2(n_163),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_198),
.B(n_200),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_185),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_183),
.B(n_3),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_150),
.C(n_166),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_215),
.C(n_193),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_147),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_211),
.Y(n_225)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_209),
.A2(n_186),
.B(n_175),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_162),
.B1(n_147),
.B2(n_149),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_179),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_148),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_212),
.B(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_213),
.B(n_216),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_165),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_165),
.C(n_163),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_187),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_215),
.A2(n_176),
.B1(n_182),
.B2(n_195),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_228),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_230),
.C(n_231),
.Y(n_232)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

BUFx12_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

NOR3xp33_ASAP7_75t_SL g230 ( 
.A(n_202),
.B(n_178),
.C(n_195),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_206),
.C(n_205),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_235),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_212),
.C(n_211),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_198),
.C(n_208),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_240),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_183),
.C(n_207),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_230),
.B(n_2),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_242),
.A2(n_221),
.B1(n_5),
.B2(n_6),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_2),
.C(n_4),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_219),
.B1(n_231),
.B2(n_220),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_246),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_237),
.A2(n_217),
.B(n_229),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_248),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_227),
.B1(n_229),
.B2(n_6),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_227),
.B1(n_5),
.B2(n_6),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_252),
.B(n_247),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_238),
.C(n_240),
.Y(n_254)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_253),
.C(n_244),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_4),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_258),
.B(n_260),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_239),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_235),
.B(n_8),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_261),
.A2(n_264),
.B(n_259),
.C(n_257),
.Y(n_266)
);

NOR2x1_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_14),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_9),
.C(n_10),
.Y(n_267)
);

OAI321xp33_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_262),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.C(n_9),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_263),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_270),
.B(n_13),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_11),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_272),
.B(n_12),
.Y(n_273)
);


endmodule