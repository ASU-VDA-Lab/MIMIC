module fake_netlist_1_6929_n_1224 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1224);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1224;
wire n_1173;
wire n_663;
wire n_791;
wire n_707;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_1198;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_1202;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_1196;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_1211;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_564;
wire n_353;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_1175;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_1177;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_1185;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_1217;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1197;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_476;
wire n_617;
wire n_384;
wire n_1200;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_1201;
wire n_1191;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_1194;
wire n_694;
wire n_301;
wire n_1179;
wire n_922;
wire n_465;
wire n_796;
wire n_1216;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1215;
wire n_286;
wire n_1174;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1078;
wire n_1097;
wire n_572;
wire n_1017;
wire n_324;
wire n_1016;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1169;
wire n_1204;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_1042;
wire n_1060;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_1222;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_1183;
wire n_567;
wire n_809;
wire n_888;
wire n_1188;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1011;
wire n_1025;
wire n_1132;
wire n_880;
wire n_1101;
wire n_1159;
wire n_630;
wire n_1155;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_1180;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_769;
wire n_624;
wire n_426;
wire n_725;
wire n_818;
wire n_844;
wire n_1160;
wire n_1184;
wire n_274;
wire n_1018;
wire n_1195;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_533;
wire n_506;
wire n_490;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_1171;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_1212;
wire n_696;
wire n_735;
wire n_771;
wire n_1091;
wire n_1203;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_1220;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_805;
wire n_729;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_1186;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_1157;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_1206;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_1178;
wire n_1209;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1218;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_1041;
wire n_578;
wire n_926;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1210;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_875;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_1214;
wire n_996;
wire n_1176;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_666;
wire n_423;
wire n_342;
wire n_621;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_1181;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_716;
wire n_357;
wire n_653;
wire n_899;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_1199;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_1221;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_1170;
wire n_419;
wire n_1193;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_1208;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_912;
wire n_620;
wire n_841;
wire n_947;
wire n_924;
wire n_1043;
wire n_1141;
wire n_378;
wire n_582;
wire n_1213;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_1189;
wire n_923;
wire n_1205;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_1172;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_1182;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_1223;
wire n_774;
wire n_1207;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_1187;
wire n_742;
wire n_1120;
wire n_1219;
wire n_585;
wire n_913;
wire n_845;
wire n_1190;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1146;
wire n_287;
wire n_1108;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_1192;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
wire n_269;
INVx1_ASAP7_75t_L g264 ( .A(n_24), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_184), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_87), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_203), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_240), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_172), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_24), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_162), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_12), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_197), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_47), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_135), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_150), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_263), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_35), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_53), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_84), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_56), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_183), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_105), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_15), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_257), .Y(n_285) );
INVxp67_ASAP7_75t_L g286 ( .A(n_237), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_13), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_51), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_222), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_110), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_206), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_189), .Y(n_292) );
INVxp67_ASAP7_75t_SL g293 ( .A(n_108), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_218), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_100), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_148), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_179), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_221), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_11), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_64), .Y(n_300) );
INVxp67_ASAP7_75t_SL g301 ( .A(n_173), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_59), .Y(n_302) );
INVxp33_ASAP7_75t_SL g303 ( .A(n_243), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_232), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_98), .Y(n_305) );
INVx1_ASAP7_75t_SL g306 ( .A(n_164), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_86), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_39), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_194), .Y(n_309) );
INVxp33_ASAP7_75t_L g310 ( .A(n_65), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_72), .Y(n_311) );
INVxp33_ASAP7_75t_SL g312 ( .A(n_177), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_242), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_71), .Y(n_314) );
CKINVDCx16_ASAP7_75t_R g315 ( .A(n_181), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_163), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_216), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_43), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_85), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_256), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_42), .Y(n_321) );
INVxp33_ASAP7_75t_SL g322 ( .A(n_182), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_174), .Y(n_323) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_45), .Y(n_324) );
INVxp67_ASAP7_75t_L g325 ( .A(n_193), .Y(n_325) );
BUFx2_ASAP7_75t_SL g326 ( .A(n_90), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_33), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_255), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_19), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_9), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_228), .Y(n_331) );
INVxp33_ASAP7_75t_L g332 ( .A(n_230), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_234), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_45), .Y(n_334) );
CKINVDCx14_ASAP7_75t_R g335 ( .A(n_125), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_54), .Y(n_336) );
INVxp33_ASAP7_75t_SL g337 ( .A(n_77), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_202), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_138), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_205), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_55), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_123), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_9), .Y(n_343) );
INVxp67_ASAP7_75t_L g344 ( .A(n_8), .Y(n_344) );
CKINVDCx16_ASAP7_75t_R g345 ( .A(n_159), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_213), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_251), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_68), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_258), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_20), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_145), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_168), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_115), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_137), .Y(n_354) );
CKINVDCx14_ASAP7_75t_R g355 ( .A(n_191), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_208), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_12), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_19), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_196), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_112), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_25), .Y(n_361) );
INVxp67_ASAP7_75t_SL g362 ( .A(n_47), .Y(n_362) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_126), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_244), .Y(n_364) );
CKINVDCx16_ASAP7_75t_R g365 ( .A(n_199), .Y(n_365) );
INVxp33_ASAP7_75t_SL g366 ( .A(n_175), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_36), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_64), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_130), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_169), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_259), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_209), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_212), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_8), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_109), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_102), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_142), .Y(n_377) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_156), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_78), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_40), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_74), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_29), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_250), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_176), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_11), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_253), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_188), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_80), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_77), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_55), .Y(n_390) );
BUFx2_ASAP7_75t_SL g391 ( .A(n_235), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_20), .Y(n_392) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_161), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_220), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_94), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_118), .Y(n_396) );
INVxp67_ASAP7_75t_L g397 ( .A(n_97), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_146), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_151), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_57), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_171), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_300), .B(n_0), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_290), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_300), .B(n_0), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_320), .Y(n_405) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_320), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_331), .B(n_1), .Y(n_407) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_320), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_265), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_265), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_310), .B(n_1), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_320), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_332), .B(n_2), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_284), .Y(n_414) );
INVxp67_ASAP7_75t_L g415 ( .A(n_284), .Y(n_415) );
INVx4_ASAP7_75t_L g416 ( .A(n_321), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_344), .B(n_2), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_266), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_321), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_264), .B(n_3), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_320), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_274), .B(n_288), .Y(n_422) );
INVx3_ASAP7_75t_L g423 ( .A(n_290), .Y(n_423) );
INVx3_ASAP7_75t_L g424 ( .A(n_309), .Y(n_424) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_354), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_354), .Y(n_426) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_354), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_315), .B(n_3), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_343), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_264), .B(n_4), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_345), .B(n_4), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_266), .Y(n_432) );
BUFx8_ASAP7_75t_L g433 ( .A(n_354), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_282), .Y(n_434) );
INVx4_ASAP7_75t_L g435 ( .A(n_416), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_405), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_403), .Y(n_437) );
AND2x2_ASAP7_75t_SL g438 ( .A(n_402), .B(n_365), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_403), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_405), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_416), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_416), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_418), .B(n_309), .Y(n_443) );
INVxp33_ASAP7_75t_L g444 ( .A(n_402), .Y(n_444) );
NAND3x1_ASAP7_75t_L g445 ( .A(n_402), .B(n_285), .C(n_282), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_403), .Y(n_446) );
INVx2_ASAP7_75t_SL g447 ( .A(n_433), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_403), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_419), .B(n_335), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_405), .Y(n_451) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_419), .Y(n_452) );
OAI221xp5_ASAP7_75t_L g453 ( .A1(n_420), .A2(n_330), .B1(n_362), .B2(n_329), .C(n_324), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_418), .A2(n_381), .B1(n_337), .B2(n_311), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_428), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_404), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_403), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_405), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_418), .B(n_333), .Y(n_459) );
AND2x6_ASAP7_75t_L g460 ( .A(n_404), .B(n_401), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_414), .B(n_415), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_405), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_403), .Y(n_463) );
XOR2x2_ASAP7_75t_L g464 ( .A(n_428), .B(n_337), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_405), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_429), .B(n_343), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_405), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_429), .B(n_355), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_431), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_423), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_405), .Y(n_471) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_405), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_423), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_414), .B(n_274), .Y(n_474) );
AND3x4_ASAP7_75t_L g475 ( .A(n_422), .B(n_357), .C(n_288), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_423), .Y(n_476) );
INVx4_ASAP7_75t_L g477 ( .A(n_416), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_423), .Y(n_478) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_406), .Y(n_479) );
AND3x1_ASAP7_75t_SL g480 ( .A(n_453), .B(n_279), .C(n_278), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_461), .B(n_415), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_447), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_438), .A2(n_413), .B1(n_431), .B2(n_404), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_469), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_449), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_461), .A2(n_434), .B(n_432), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_452), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_452), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_469), .Y(n_489) );
INVx4_ASAP7_75t_L g490 ( .A(n_447), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_437), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_466), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_466), .Y(n_493) );
NAND2xp33_ASAP7_75t_L g494 ( .A(n_460), .B(n_431), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_456), .Y(n_495) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_447), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_438), .A2(n_413), .B1(n_411), .B2(n_407), .Y(n_497) );
INVx3_ASAP7_75t_L g498 ( .A(n_460), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_450), .B(n_413), .Y(n_499) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_460), .Y(n_500) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_460), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_450), .B(n_411), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_437), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_438), .A2(n_407), .B1(n_417), .B2(n_311), .Y(n_504) );
BUFx8_ASAP7_75t_L g505 ( .A(n_460), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_444), .B(n_409), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_435), .B(n_432), .Y(n_507) );
INVx3_ASAP7_75t_L g508 ( .A(n_460), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_468), .B(n_409), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_466), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_439), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_444), .B(n_410), .Y(n_512) );
NAND2x2_ASAP7_75t_L g513 ( .A(n_464), .B(n_420), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_438), .A2(n_417), .B1(n_368), .B2(n_390), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_468), .B(n_410), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_439), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_460), .A2(n_368), .B1(n_390), .B2(n_270), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_456), .A2(n_280), .B1(n_328), .B2(n_295), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_466), .B(n_432), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_466), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_446), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_468), .B(n_270), .Y(n_522) );
OR2x6_ASAP7_75t_L g523 ( .A(n_454), .B(n_430), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_446), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_460), .B(n_422), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_454), .B(n_430), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_460), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_448), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_448), .Y(n_529) );
BUFx2_ASAP7_75t_L g530 ( .A(n_455), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_457), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_457), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_464), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_463), .Y(n_534) );
OR2x6_ASAP7_75t_L g535 ( .A(n_445), .B(n_422), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_464), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_475), .Y(n_537) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_463), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_470), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_474), .B(n_434), .Y(n_540) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_470), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_475), .A2(n_434), .B1(n_312), .B2(n_322), .Y(n_542) );
INVx5_ASAP7_75t_L g543 ( .A(n_435), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_473), .Y(n_544) );
BUFx3_ASAP7_75t_L g545 ( .A(n_475), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_474), .B(n_416), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_473), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_474), .B(n_422), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_476), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_474), .B(n_422), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_445), .B(n_416), .Y(n_551) );
NOR2xp67_ASAP7_75t_L g552 ( .A(n_453), .B(n_423), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_475), .Y(n_553) );
BUFx3_ASAP7_75t_L g554 ( .A(n_476), .Y(n_554) );
INVx6_ASAP7_75t_L g555 ( .A(n_435), .Y(n_555) );
AND2x4_ASAP7_75t_L g556 ( .A(n_443), .B(n_272), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_478), .Y(n_557) );
CKINVDCx8_ASAP7_75t_R g558 ( .A(n_445), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_478), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_441), .Y(n_560) );
INVx3_ASAP7_75t_L g561 ( .A(n_435), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_441), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_443), .B(n_272), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_525), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_483), .A2(n_312), .B1(n_322), .B2(n_303), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_499), .B(n_459), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_505), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_502), .B(n_459), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_484), .B(n_423), .Y(n_569) );
BUFx3_ASAP7_75t_L g570 ( .A(n_505), .Y(n_570) );
OR2x6_ASAP7_75t_L g571 ( .A(n_500), .B(n_326), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_525), .B(n_281), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_484), .B(n_424), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_525), .B(n_281), .Y(n_574) );
BUFx2_ASAP7_75t_L g575 ( .A(n_505), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_487), .B(n_287), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_533), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_535), .A2(n_366), .B1(n_303), .B2(n_318), .Y(n_578) );
INVx3_ASAP7_75t_L g579 ( .A(n_500), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_492), .Y(n_580) );
BUFx2_ASAP7_75t_L g581 ( .A(n_500), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_493), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_560), .Y(n_583) );
AOI222xp33_ASAP7_75t_L g584 ( .A1(n_536), .A2(n_361), .B1(n_400), .B2(n_287), .C1(n_392), .C2(n_299), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_560), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_535), .A2(n_366), .B1(n_327), .B2(n_334), .Y(n_586) );
INVx6_ASAP7_75t_L g587 ( .A(n_543), .Y(n_587) );
BUFx3_ASAP7_75t_L g588 ( .A(n_500), .Y(n_588) );
OAI22xp5_ASAP7_75t_SL g589 ( .A1(n_536), .A2(n_339), .B1(n_342), .B2(n_316), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_501), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_481), .B(n_316), .Y(n_591) );
NOR2x1_ASAP7_75t_SL g592 ( .A(n_501), .B(n_326), .Y(n_592) );
BUFx12f_ASAP7_75t_L g593 ( .A(n_530), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_489), .B(n_424), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_510), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_562), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_562), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_L g598 ( .A1(n_489), .A2(n_336), .B(n_341), .C(n_314), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_520), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_523), .A2(n_342), .B1(n_359), .B2(n_339), .Y(n_600) );
BUFx8_ASAP7_75t_L g601 ( .A(n_501), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_491), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_501), .Y(n_603) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_527), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_491), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_495), .B(n_435), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_535), .A2(n_350), .B1(n_358), .B2(n_348), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_523), .A2(n_380), .B1(n_382), .B2(n_374), .Y(n_608) );
BUFx3_ASAP7_75t_L g609 ( .A(n_527), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_503), .Y(n_610) );
INVxp67_ASAP7_75t_SL g611 ( .A(n_527), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_481), .B(n_359), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_523), .B(n_299), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_503), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_527), .A2(n_386), .B1(n_387), .B2(n_373), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_511), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_550), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_488), .B(n_302), .Y(n_618) );
BUFx3_ASAP7_75t_L g619 ( .A(n_543), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_526), .B(n_424), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_511), .Y(n_621) );
AOI21xp33_ASAP7_75t_L g622 ( .A1(n_494), .A2(n_386), .B(n_373), .Y(n_622) );
BUFx2_ASAP7_75t_L g623 ( .A(n_545), .Y(n_623) );
INVxp33_ASAP7_75t_L g624 ( .A(n_518), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_494), .A2(n_385), .B1(n_308), .B2(n_361), .Y(n_625) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_482), .Y(n_626) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_482), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_516), .Y(n_628) );
BUFx3_ASAP7_75t_L g629 ( .A(n_543), .Y(n_629) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_490), .Y(n_630) );
BUFx2_ASAP7_75t_L g631 ( .A(n_545), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_558), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_506), .B(n_387), .Y(n_633) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_490), .Y(n_634) );
BUFx3_ASAP7_75t_L g635 ( .A(n_543), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_507), .A2(n_442), .B(n_441), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_509), .A2(n_308), .B(n_388), .C(n_302), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_516), .Y(n_638) );
INVx3_ASAP7_75t_L g639 ( .A(n_498), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_537), .A2(n_389), .B1(n_392), .B2(n_388), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_558), .Y(n_641) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_537), .A2(n_396), .B1(n_391), .B2(n_389), .Y(n_642) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_490), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_522), .Y(n_644) );
BUFx2_ASAP7_75t_L g645 ( .A(n_553), .Y(n_645) );
INVx3_ASAP7_75t_L g646 ( .A(n_498), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_542), .A2(n_396), .B1(n_400), .B2(n_293), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_553), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_506), .B(n_477), .Y(n_649) );
BUFx2_ASAP7_75t_L g650 ( .A(n_508), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_515), .B(n_424), .Y(n_651) );
NAND2x1p5_ASAP7_75t_L g652 ( .A(n_508), .B(n_477), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_548), .Y(n_653) );
BUFx3_ASAP7_75t_L g654 ( .A(n_548), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_529), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_540), .Y(n_656) );
BUFx3_ASAP7_75t_L g657 ( .A(n_555), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_512), .B(n_424), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_529), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_497), .A2(n_301), .B1(n_363), .B2(n_283), .Y(n_660) );
CKINVDCx6p67_ASAP7_75t_R g661 ( .A(n_551), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_534), .Y(n_662) );
BUFx2_ASAP7_75t_L g663 ( .A(n_554), .Y(n_663) );
BUFx2_ASAP7_75t_L g664 ( .A(n_554), .Y(n_664) );
BUFx12f_ASAP7_75t_L g665 ( .A(n_556), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_485), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_512), .B(n_424), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_546), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_519), .B(n_357), .Y(n_669) );
BUFx12f_ASAP7_75t_L g670 ( .A(n_556), .Y(n_670) );
OR2x6_ASAP7_75t_L g671 ( .A(n_552), .B(n_391), .Y(n_671) );
INVx3_ASAP7_75t_L g672 ( .A(n_555), .Y(n_672) );
AO21x1_ASAP7_75t_L g673 ( .A1(n_519), .A2(n_426), .B(n_289), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_521), .Y(n_674) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_496), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_534), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_486), .A2(n_379), .B(n_367), .C(n_286), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_524), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_504), .B(n_477), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_514), .B(n_477), .Y(n_680) );
AND2x6_ASAP7_75t_L g681 ( .A(n_561), .B(n_285), .Y(n_681) );
AND2x4_ASAP7_75t_SL g682 ( .A(n_517), .B(n_367), .Y(n_682) );
A2O1A1Ixp33_ASAP7_75t_L g683 ( .A1(n_528), .A2(n_379), .B(n_291), .C(n_296), .Y(n_683) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_513), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_531), .Y(n_685) );
OAI22xp33_ASAP7_75t_L g686 ( .A1(n_624), .A2(n_513), .B1(n_480), .B2(n_556), .Y(n_686) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_645), .A2(n_563), .B1(n_480), .B2(n_294), .Y(n_687) );
NAND2x1p5_ASAP7_75t_L g688 ( .A(n_570), .B(n_561), .Y(n_688) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_663), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_624), .B(n_507), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_602), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_636), .A2(n_539), .B(n_532), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_645), .A2(n_563), .B1(n_547), .B2(n_557), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_666), .B(n_563), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_677), .A2(n_549), .B(n_559), .C(n_544), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_602), .Y(n_696) );
NOR2xp67_ASAP7_75t_SL g697 ( .A(n_567), .B(n_555), .Y(n_697) );
CKINVDCx5p33_ASAP7_75t_R g698 ( .A(n_593), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_632), .A2(n_294), .B1(n_372), .B2(n_292), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_665), .A2(n_559), .B1(n_544), .B2(n_538), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_600), .A2(n_541), .B(n_538), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_613), .A2(n_538), .B1(n_541), .B2(n_496), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_572), .A2(n_541), .B1(n_538), .B2(n_291), .Y(n_703) );
OAI22xp33_ASAP7_75t_SL g704 ( .A1(n_613), .A2(n_296), .B1(n_297), .B2(n_289), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_644), .B(n_541), .Y(n_705) );
AND2x4_ASAP7_75t_L g706 ( .A(n_564), .B(n_496), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_589), .A2(n_496), .B1(n_371), .B2(n_393), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_651), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_648), .B(n_5), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_584), .B(n_6), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_651), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_569), .Y(n_712) );
CKINVDCx6p67_ASAP7_75t_R g713 ( .A(n_593), .Y(n_713) );
OR2x2_ASAP7_75t_L g714 ( .A(n_572), .B(n_6), .Y(n_714) );
INVx8_ASAP7_75t_L g715 ( .A(n_665), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_684), .B(n_7), .Y(n_716) );
AO31x2_ASAP7_75t_L g717 ( .A1(n_673), .A2(n_426), .A3(n_304), .B(n_305), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_670), .A2(n_304), .B1(n_305), .B2(n_297), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_670), .A2(n_313), .B1(n_360), .B2(n_307), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_654), .A2(n_313), .B1(n_360), .B2(n_307), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_569), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_663), .A2(n_377), .B1(n_397), .B2(n_325), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_572), .B(n_7), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_573), .Y(n_724) );
BUFx6f_ASAP7_75t_L g725 ( .A(n_604), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_574), .A2(n_395), .B1(n_398), .B2(n_364), .Y(n_726) );
OR2x6_ASAP7_75t_L g727 ( .A(n_575), .B(n_364), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_605), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_679), .A2(n_442), .B(n_441), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_573), .Y(n_730) );
OAI21x1_ASAP7_75t_SL g731 ( .A1(n_673), .A2(n_398), .B(n_395), .Y(n_731) );
BUFx2_ASAP7_75t_L g732 ( .A(n_601), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_594), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_608), .B(n_441), .Y(n_734) );
A2O1A1Ixp33_ASAP7_75t_L g735 ( .A1(n_637), .A2(n_401), .B(n_399), .C(n_268), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_594), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_565), .B(n_442), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_654), .B(n_442), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_610), .Y(n_739) );
INVx6_ASAP7_75t_SL g740 ( .A(n_574), .Y(n_740) );
OAI221xp5_ASAP7_75t_L g741 ( .A1(n_660), .A2(n_399), .B1(n_269), .B2(n_271), .C(n_273), .Y(n_741) );
BUFx12f_ASAP7_75t_L g742 ( .A(n_601), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_576), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_664), .A2(n_306), .B1(n_298), .B2(n_275), .Y(n_744) );
BUFx6f_ASAP7_75t_L g745 ( .A(n_604), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_576), .Y(n_746) );
O2A1O1Ixp5_ASAP7_75t_L g747 ( .A1(n_683), .A2(n_369), .B(n_394), .C(n_333), .Y(n_747) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_598), .A2(n_375), .B1(n_276), .B2(n_277), .C(n_317), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_576), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_610), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_618), .Y(n_751) );
AOI211xp5_ASAP7_75t_L g752 ( .A1(n_622), .A2(n_319), .B(n_323), .C(n_267), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_623), .B(n_10), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_680), .A2(n_442), .B(n_440), .Y(n_754) );
OAI22xp33_ASAP7_75t_L g755 ( .A1(n_632), .A2(n_372), .B1(n_292), .B2(n_340), .Y(n_755) );
CKINVDCx14_ASAP7_75t_R g756 ( .A(n_577), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_617), .B(n_338), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_618), .Y(n_758) );
INVx1_ASAP7_75t_SL g759 ( .A(n_664), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_623), .A2(n_347), .B1(n_349), .B2(n_346), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_618), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_674), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_678), .Y(n_763) );
OR2x6_ASAP7_75t_L g764 ( .A(n_575), .B(n_351), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_685), .Y(n_765) );
AOI22xp33_ASAP7_75t_SL g766 ( .A1(n_641), .A2(n_353), .B1(n_356), .B2(n_352), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_656), .B(n_370), .Y(n_767) );
AOI221xp5_ASAP7_75t_L g768 ( .A1(n_620), .A2(n_376), .B1(n_383), .B2(n_384), .C(n_354), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_620), .B(n_13), .Y(n_769) );
AO221x2_ASAP7_75t_L g770 ( .A1(n_615), .A2(n_14), .B1(n_15), .B2(n_16), .C(n_17), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_625), .A2(n_426), .B1(n_378), .B2(n_408), .Y(n_771) );
A2O1A1Ixp33_ASAP7_75t_L g772 ( .A1(n_566), .A2(n_378), .B(n_406), .C(n_408), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_682), .A2(n_378), .B1(n_406), .B2(n_408), .Y(n_773) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_614), .Y(n_774) );
BUFx2_ASAP7_75t_SL g775 ( .A(n_619), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_616), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_631), .B(n_14), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_682), .A2(n_378), .B1(n_406), .B2(n_408), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_631), .B(n_17), .Y(n_779) );
O2A1O1Ixp5_ASAP7_75t_L g780 ( .A1(n_683), .A2(n_436), .B(n_440), .C(n_471), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_580), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_616), .Y(n_782) );
A2O1A1Ixp33_ASAP7_75t_L g783 ( .A1(n_568), .A2(n_378), .B(n_406), .C(n_408), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_668), .A2(n_433), .B1(n_408), .B2(n_412), .Y(n_784) );
O2A1O1Ixp5_ASAP7_75t_L g785 ( .A1(n_658), .A2(n_440), .B(n_451), .C(n_471), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_653), .A2(n_433), .B1(n_408), .B2(n_412), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_621), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g788 ( .A1(n_671), .A2(n_18), .B1(n_21), .B2(n_22), .Y(n_788) );
NAND2x1p5_ASAP7_75t_L g789 ( .A(n_588), .B(n_406), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_647), .B(n_18), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_582), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_640), .B(n_21), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_658), .A2(n_433), .B1(n_408), .B2(n_412), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_567), .Y(n_794) );
OAI22xp33_ASAP7_75t_L g795 ( .A1(n_671), .A2(n_22), .B1(n_23), .B2(n_25), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_578), .B(n_23), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_595), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_586), .A2(n_433), .B1(n_408), .B2(n_412), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_628), .A2(n_406), .B1(n_412), .B2(n_421), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_606), .A2(n_433), .B1(n_412), .B2(n_421), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_628), .A2(n_406), .B1(n_412), .B2(n_421), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_649), .A2(n_451), .B(n_436), .Y(n_802) );
AND2x4_ASAP7_75t_L g803 ( .A(n_619), .B(n_26), .Y(n_803) );
AO21x2_ASAP7_75t_L g804 ( .A1(n_592), .A2(n_451), .B(n_436), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_638), .Y(n_805) );
OAI21x1_ASAP7_75t_L g806 ( .A1(n_638), .A2(n_465), .B(n_462), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_655), .A2(n_406), .B1(n_412), .B2(n_421), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_667), .A2(n_412), .B1(n_421), .B2(n_425), .Y(n_808) );
BUFx3_ASAP7_75t_L g809 ( .A(n_629), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_762), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_686), .A2(n_671), .B1(n_642), .B2(n_667), .Y(n_811) );
OAI221xp5_ASAP7_75t_L g812 ( .A1(n_766), .A2(n_607), .B1(n_612), .B2(n_591), .C(n_633), .Y(n_812) );
AND2x6_ASAP7_75t_L g813 ( .A(n_803), .B(n_604), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g814 ( .A1(n_710), .A2(n_681), .B1(n_571), .B2(n_669), .Y(n_814) );
AOI21xp5_ASAP7_75t_L g815 ( .A1(n_754), .A2(n_659), .B(n_655), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_686), .B(n_661), .Y(n_816) );
AO21x2_ASAP7_75t_L g817 ( .A1(n_731), .A2(n_662), .B(n_659), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_708), .B(n_669), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_774), .Y(n_819) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_774), .Y(n_820) );
OR2x2_ASAP7_75t_L g821 ( .A(n_715), .B(n_662), .Y(n_821) );
INVx3_ASAP7_75t_L g822 ( .A(n_742), .Y(n_822) );
OAI33xp33_ASAP7_75t_L g823 ( .A1(n_788), .A2(n_599), .A3(n_676), .B1(n_596), .B2(n_597), .B3(n_583), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_690), .A2(n_681), .B1(n_661), .B2(n_650), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_727), .A2(n_571), .B1(n_581), .B2(n_627), .Y(n_825) );
OAI21xp33_ASAP7_75t_L g826 ( .A1(n_699), .A2(n_571), .B(n_629), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_796), .A2(n_681), .B1(n_650), .B2(n_672), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_691), .Y(n_828) );
A2O1A1Ixp33_ASAP7_75t_L g829 ( .A1(n_737), .A2(n_635), .B(n_646), .C(n_639), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g830 ( .A1(n_754), .A2(n_585), .B(n_583), .Y(n_830) );
BUFx4f_ASAP7_75t_SL g831 ( .A(n_713), .Y(n_831) );
BUFx8_ASAP7_75t_L g832 ( .A(n_732), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g833 ( .A1(n_727), .A2(n_626), .B1(n_627), .B2(n_581), .Y(n_833) );
BUFx12f_ASAP7_75t_L g834 ( .A(n_698), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_687), .A2(n_681), .B1(n_672), .B2(n_635), .Y(n_835) );
AOI21xp5_ASAP7_75t_L g836 ( .A1(n_692), .A2(n_585), .B(n_675), .Y(n_836) );
AOI221xp5_ASAP7_75t_L g837 ( .A1(n_741), .A2(n_657), .B1(n_639), .B2(n_646), .C(n_611), .Y(n_837) );
AOI21xp33_ASAP7_75t_L g838 ( .A1(n_769), .A2(n_603), .B(n_590), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_763), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_765), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_781), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_696), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_791), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_687), .A2(n_627), .B1(n_626), .B2(n_609), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_797), .Y(n_845) );
OR2x2_ASAP7_75t_L g846 ( .A(n_715), .B(n_657), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_711), .B(n_681), .Y(n_847) );
INVx2_ASAP7_75t_L g848 ( .A(n_728), .Y(n_848) );
INVx3_ASAP7_75t_L g849 ( .A(n_688), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_764), .A2(n_681), .B1(n_639), .B2(n_646), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_714), .Y(n_851) );
OAI21xp5_ASAP7_75t_L g852 ( .A1(n_747), .A2(n_652), .B(n_603), .Y(n_852) );
BUFx3_ASAP7_75t_L g853 ( .A(n_715), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_764), .A2(n_627), .B1(n_626), .B2(n_609), .Y(n_854) );
OAI22xp33_ASAP7_75t_L g855 ( .A1(n_788), .A2(n_626), .B1(n_604), .B2(n_643), .Y(n_855) );
AOI221xp5_ASAP7_75t_L g856 ( .A1(n_748), .A2(n_579), .B1(n_590), .B2(n_652), .C(n_675), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_770), .A2(n_587), .B1(n_579), .B2(n_634), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_739), .Y(n_858) );
OAI211xp5_ASAP7_75t_SL g859 ( .A1(n_748), .A2(n_579), .B(n_465), .C(n_467), .Y(n_859) );
OAI221xp5_ASAP7_75t_SL g860 ( .A1(n_795), .A2(n_26), .B1(n_27), .B2(n_28), .C(n_29), .Y(n_860) );
OR2x6_ASAP7_75t_L g861 ( .A(n_803), .B(n_587), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_712), .B(n_587), .Y(n_862) );
BUFx2_ASAP7_75t_L g863 ( .A(n_740), .Y(n_863) );
AOI22xp33_ASAP7_75t_SL g864 ( .A1(n_770), .A2(n_587), .B1(n_643), .B2(n_634), .Y(n_864) );
AO21x2_ASAP7_75t_L g865 ( .A1(n_772), .A2(n_465), .B(n_462), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_689), .A2(n_643), .B1(n_634), .B2(n_630), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_723), .A2(n_630), .B1(n_675), .B2(n_421), .Y(n_867) );
INVxp67_ASAP7_75t_SL g868 ( .A(n_689), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_790), .A2(n_630), .B1(n_675), .B2(n_421), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_755), .A2(n_675), .B1(n_421), .B2(n_425), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_693), .A2(n_421), .B1(n_425), .B2(n_427), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_709), .A2(n_425), .B1(n_427), .B2(n_471), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_792), .A2(n_427), .B1(n_425), .B2(n_467), .Y(n_873) );
OAI221xp5_ASAP7_75t_L g874 ( .A1(n_766), .A2(n_427), .B1(n_425), .B2(n_467), .C(n_462), .Y(n_874) );
OAI21x1_ASAP7_75t_L g875 ( .A1(n_806), .A2(n_427), .B(n_425), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_721), .B(n_27), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_753), .A2(n_427), .B1(n_425), .B2(n_458), .Y(n_877) );
AOI21xp5_ASAP7_75t_L g878 ( .A1(n_692), .A2(n_427), .B(n_425), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_743), .Y(n_879) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_759), .A2(n_427), .B1(n_472), .B2(n_458), .Y(n_880) );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_704), .A2(n_427), .B1(n_472), .B2(n_458), .C(n_479), .Y(n_881) );
AOI21xp33_ASAP7_75t_L g882 ( .A1(n_752), .A2(n_28), .B(n_30), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g883 ( .A1(n_724), .A2(n_479), .B1(n_472), .B2(n_458), .C(n_34), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_730), .B(n_30), .Y(n_884) );
OAI21x1_ASAP7_75t_L g885 ( .A1(n_785), .A2(n_472), .B(n_458), .Y(n_885) );
OAI221xp5_ASAP7_75t_L g886 ( .A1(n_718), .A2(n_479), .B1(n_472), .B2(n_34), .C(n_35), .Y(n_886) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_699), .B(n_479), .C(n_31), .Y(n_887) );
OA21x2_ASAP7_75t_L g888 ( .A1(n_783), .A2(n_479), .B(n_88), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_716), .B(n_31), .Y(n_889) );
OAI211xp5_ASAP7_75t_SL g890 ( .A1(n_719), .A2(n_32), .B(n_36), .C(n_37), .Y(n_890) );
OAI22xp33_ASAP7_75t_L g891 ( .A1(n_740), .A2(n_37), .B1(n_38), .B2(n_39), .Y(n_891) );
INVx3_ASAP7_75t_L g892 ( .A(n_688), .Y(n_892) );
OAI22xp33_ASAP7_75t_L g893 ( .A1(n_694), .A2(n_38), .B1(n_40), .B2(n_41), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_777), .B(n_41), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_726), .A2(n_42), .B1(n_43), .B2(n_44), .Y(n_895) );
AO21x2_ASAP7_75t_L g896 ( .A1(n_695), .A2(n_89), .B(n_83), .Y(n_896) );
AOI221xp5_ASAP7_75t_L g897 ( .A1(n_733), .A2(n_44), .B1(n_46), .B2(n_48), .C(n_49), .Y(n_897) );
BUFx6f_ASAP7_75t_L g898 ( .A(n_725), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_726), .A2(n_46), .B1(n_48), .B2(n_49), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_746), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_779), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_901) );
AOI21xp33_ASAP7_75t_SL g902 ( .A1(n_744), .A2(n_50), .B(n_52), .Y(n_902) );
BUFx6f_ASAP7_75t_L g903 ( .A(n_725), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_736), .A2(n_56), .B1(n_57), .B2(n_58), .Y(n_904) );
AO21x2_ASAP7_75t_L g905 ( .A1(n_701), .A2(n_92), .B(n_91), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_749), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_906) );
OAI221xp5_ASAP7_75t_L g907 ( .A1(n_735), .A2(n_60), .B1(n_61), .B2(n_62), .C(n_63), .Y(n_907) );
OAI21x1_ASAP7_75t_L g908 ( .A1(n_785), .A2(n_154), .B(n_261), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_703), .A2(n_61), .B1(n_62), .B2(n_63), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_751), .B(n_65), .Y(n_910) );
OAI211xp5_ASAP7_75t_SL g911 ( .A1(n_768), .A2(n_66), .B(n_67), .C(n_68), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_758), .A2(n_761), .B1(n_768), .B2(n_756), .Y(n_912) );
AOI21xp5_ASAP7_75t_L g913 ( .A1(n_802), .A2(n_157), .B(n_260), .Y(n_913) );
BUFx2_ASAP7_75t_L g914 ( .A(n_794), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_703), .A2(n_66), .B1(n_67), .B2(n_69), .Y(n_915) );
OAI21x1_ASAP7_75t_L g916 ( .A1(n_802), .A2(n_158), .B(n_254), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_757), .B(n_69), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_738), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_767), .B(n_760), .Y(n_919) );
OAI322xp33_ASAP7_75t_L g920 ( .A1(n_891), .A2(n_722), .A3(n_707), .B1(n_705), .B2(n_734), .C1(n_771), .C2(n_778), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_816), .A2(n_798), .B1(n_775), .B2(n_793), .Y(n_921) );
OAI221xp5_ASAP7_75t_L g922 ( .A1(n_912), .A2(n_720), .B1(n_793), .B2(n_700), .C(n_784), .Y(n_922) );
OA21x2_ASAP7_75t_L g923 ( .A1(n_878), .A2(n_780), .B(n_808), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_828), .Y(n_924) );
INVx2_ASAP7_75t_L g925 ( .A(n_842), .Y(n_925) );
OAI33xp33_ASAP7_75t_L g926 ( .A1(n_891), .A2(n_773), .A3(n_799), .B1(n_807), .B2(n_801), .B3(n_702), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_848), .Y(n_927) );
INVxp67_ASAP7_75t_SL g928 ( .A(n_868), .Y(n_928) );
OAI221xp5_ASAP7_75t_L g929 ( .A1(n_811), .A2(n_786), .B1(n_800), .B2(n_808), .C(n_809), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_814), .A2(n_697), .B1(n_706), .B2(n_805), .Y(n_930) );
NAND3xp33_ASAP7_75t_L g931 ( .A(n_897), .B(n_706), .C(n_787), .Y(n_931) );
NAND4xp25_ASAP7_75t_L g932 ( .A(n_860), .B(n_729), .C(n_750), .D(n_776), .Y(n_932) );
AOI21xp33_ASAP7_75t_SL g933 ( .A1(n_822), .A2(n_73), .B(n_75), .Y(n_933) );
OR2x2_ASAP7_75t_L g934 ( .A(n_868), .B(n_717), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_851), .B(n_717), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_819), .B(n_782), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_858), .B(n_717), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_820), .B(n_717), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_820), .B(n_789), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_810), .B(n_75), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_861), .B(n_789), .Y(n_941) );
OAI21x1_ASAP7_75t_L g942 ( .A1(n_885), .A2(n_745), .B(n_725), .Y(n_942) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_821), .Y(n_943) );
INVx2_ASAP7_75t_SL g944 ( .A(n_832), .Y(n_944) );
AO21x2_ASAP7_75t_L g945 ( .A1(n_836), .A2(n_804), .B(n_745), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_814), .A2(n_804), .B1(n_78), .B2(n_79), .Y(n_946) );
BUFx3_ASAP7_75t_L g947 ( .A(n_853), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_812), .A2(n_76), .B1(n_79), .B2(n_80), .Y(n_948) );
INVxp67_ASAP7_75t_L g949 ( .A(n_914), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_861), .B(n_76), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_879), .Y(n_951) );
OR2x2_ASAP7_75t_L g952 ( .A(n_839), .B(n_81), .Y(n_952) );
OR2x2_ASAP7_75t_L g953 ( .A(n_840), .B(n_81), .Y(n_953) );
BUFx3_ASAP7_75t_L g954 ( .A(n_831), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_841), .B(n_82), .Y(n_955) );
INVx2_ASAP7_75t_L g956 ( .A(n_900), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_843), .Y(n_957) );
INVx3_ASAP7_75t_L g958 ( .A(n_813), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_845), .B(n_82), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_817), .Y(n_960) );
AOI221xp5_ASAP7_75t_L g961 ( .A1(n_893), .A2(n_93), .B1(n_95), .B2(n_96), .C(n_99), .Y(n_961) );
OAI211xp5_ASAP7_75t_L g962 ( .A1(n_864), .A2(n_101), .B(n_103), .C(n_104), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_864), .B(n_106), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_898), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_919), .A2(n_107), .B1(n_111), .B2(n_113), .Y(n_965) );
INVx2_ASAP7_75t_L g966 ( .A(n_898), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_835), .A2(n_114), .B1(n_116), .B2(n_117), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_876), .Y(n_968) );
OA222x2_ASAP7_75t_L g969 ( .A1(n_822), .A2(n_119), .B1(n_120), .B2(n_121), .C1(n_122), .C2(n_124), .Y(n_969) );
AO21x2_ASAP7_75t_L g970 ( .A1(n_836), .A2(n_127), .B(n_128), .Y(n_970) );
AOI33xp33_ASAP7_75t_L g971 ( .A1(n_893), .A2(n_129), .A3(n_131), .B1(n_132), .B2(n_133), .B3(n_134), .Y(n_971) );
OAI221xp5_ASAP7_75t_L g972 ( .A1(n_882), .A2(n_136), .B1(n_139), .B2(n_140), .C(n_141), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g973 ( .A1(n_813), .A2(n_143), .B1(n_144), .B2(n_147), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_894), .B(n_149), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_817), .Y(n_975) );
OAI221xp5_ASAP7_75t_L g976 ( .A1(n_826), .A2(n_152), .B1(n_153), .B2(n_155), .C(n_160), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_815), .Y(n_977) );
HB1xp67_ASAP7_75t_L g978 ( .A(n_846), .Y(n_978) );
NAND4xp25_ASAP7_75t_L g979 ( .A(n_901), .B(n_165), .C(n_166), .D(n_167), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_911), .A2(n_170), .B1(n_178), .B2(n_180), .Y(n_980) );
INVx2_ASAP7_75t_L g981 ( .A(n_898), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g982 ( .A1(n_857), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_982) );
AND2x4_ASAP7_75t_SL g983 ( .A(n_849), .B(n_262), .Y(n_983) );
BUFx3_ASAP7_75t_L g984 ( .A(n_813), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_911), .A2(n_190), .B1(n_192), .B2(n_195), .Y(n_985) );
OAI221xp5_ASAP7_75t_L g986 ( .A1(n_827), .A2(n_198), .B1(n_200), .B2(n_201), .C(n_204), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_815), .Y(n_987) );
OAI31xp33_ASAP7_75t_L g988 ( .A1(n_890), .A2(n_207), .A3(n_210), .B(n_211), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_830), .Y(n_989) );
OAI211xp5_ASAP7_75t_SL g990 ( .A1(n_918), .A2(n_214), .B(n_215), .C(n_217), .Y(n_990) );
AND2x4_ASAP7_75t_L g991 ( .A(n_849), .B(n_219), .Y(n_991) );
NAND3xp33_ASAP7_75t_L g992 ( .A(n_902), .B(n_223), .C(n_224), .Y(n_992) );
NOR2xp33_ASAP7_75t_L g993 ( .A(n_863), .B(n_225), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_890), .A2(n_226), .B1(n_227), .B2(n_229), .Y(n_994) );
OR2x2_ASAP7_75t_L g995 ( .A(n_818), .B(n_884), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_903), .Y(n_996) );
NAND4xp25_ASAP7_75t_L g997 ( .A(n_889), .B(n_231), .C(n_233), .D(n_236), .Y(n_997) );
OR2x2_ASAP7_75t_L g998 ( .A(n_910), .B(n_238), .Y(n_998) );
OAI221xp5_ASAP7_75t_SL g999 ( .A1(n_907), .A2(n_239), .B1(n_241), .B2(n_245), .C(n_246), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_892), .B(n_247), .Y(n_1000) );
BUFx3_ASAP7_75t_L g1001 ( .A(n_813), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g1002 ( .A1(n_895), .A2(n_248), .B1(n_249), .B2(n_252), .C(n_899), .Y(n_1002) );
OAI221xp5_ASAP7_75t_L g1003 ( .A1(n_917), .A2(n_850), .B1(n_824), .B2(n_886), .C(n_887), .Y(n_1003) );
AOI222xp33_ASAP7_75t_L g1004 ( .A1(n_909), .A2(n_915), .B1(n_823), .B2(n_904), .C1(n_906), .C2(n_813), .Y(n_1004) );
OAI332xp33_ASAP7_75t_SL g1005 ( .A1(n_833), .A2(n_854), .A3(n_855), .B1(n_871), .B2(n_825), .B3(n_866), .C1(n_844), .C2(n_834), .Y(n_1005) );
INVx2_ASAP7_75t_L g1006 ( .A(n_977), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_938), .B(n_896), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_1003), .A2(n_859), .B1(n_881), .B2(n_856), .Y(n_1008) );
OR2x2_ASAP7_75t_L g1009 ( .A(n_928), .B(n_833), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_938), .B(n_903), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1011 ( .A1(n_921), .A2(n_870), .B1(n_847), .B2(n_892), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_937), .B(n_903), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_937), .B(n_865), .Y(n_1013) );
OR2x2_ASAP7_75t_L g1014 ( .A(n_934), .B(n_862), .Y(n_1014) );
OR2x2_ASAP7_75t_L g1015 ( .A(n_934), .B(n_830), .Y(n_1015) );
OAI21x1_ASAP7_75t_L g1016 ( .A1(n_942), .A2(n_908), .B(n_875), .Y(n_1016) );
AOI211xp5_ASAP7_75t_L g1017 ( .A1(n_997), .A2(n_859), .B(n_874), .C(n_913), .Y(n_1017) );
INVx2_ASAP7_75t_L g1018 ( .A(n_977), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_960), .Y(n_1019) );
INVx3_ASAP7_75t_L g1020 ( .A(n_945), .Y(n_1020) );
INVxp67_ASAP7_75t_SL g1021 ( .A(n_943), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_975), .Y(n_1022) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_930), .A2(n_867), .B1(n_869), .B2(n_829), .Y(n_1023) );
INVx2_ASAP7_75t_SL g1024 ( .A(n_939), .Y(n_1024) );
AO21x2_ASAP7_75t_L g1025 ( .A1(n_975), .A2(n_865), .B(n_905), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_957), .B(n_905), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_957), .B(n_852), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_951), .B(n_883), .Y(n_1028) );
INVx2_ASAP7_75t_L g1029 ( .A(n_987), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_935), .Y(n_1030) );
AOI31xp33_ASAP7_75t_L g1031 ( .A1(n_944), .A2(n_913), .A3(n_877), .B(n_837), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_989), .Y(n_1032) );
AOI33xp33_ASAP7_75t_L g1033 ( .A1(n_968), .A2(n_872), .A3(n_873), .B1(n_880), .B2(n_888), .B3(n_838), .Y(n_1033) );
INVx1_ASAP7_75t_SL g1034 ( .A(n_947), .Y(n_1034) );
HB1xp67_ASAP7_75t_L g1035 ( .A(n_978), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_989), .Y(n_1036) );
OAI221xp5_ASAP7_75t_L g1037 ( .A1(n_948), .A2(n_888), .B1(n_916), .B2(n_949), .C(n_946), .Y(n_1037) );
HB1xp67_ASAP7_75t_L g1038 ( .A(n_939), .Y(n_1038) );
AND2x4_ASAP7_75t_L g1039 ( .A(n_945), .B(n_958), .Y(n_1039) );
NAND2xp5_ASAP7_75t_SL g1040 ( .A(n_963), .B(n_958), .Y(n_1040) );
NAND4xp25_ASAP7_75t_L g1041 ( .A(n_952), .B(n_953), .C(n_950), .D(n_940), .Y(n_1041) );
OAI21xp33_ASAP7_75t_L g1042 ( .A1(n_971), .A2(n_979), .B(n_953), .Y(n_1042) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_956), .B(n_952), .Y(n_1043) );
BUFx3_ASAP7_75t_L g1044 ( .A(n_984), .Y(n_1044) );
HB1xp67_ASAP7_75t_L g1045 ( .A(n_936), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_995), .B(n_959), .Y(n_1046) );
INVx2_ASAP7_75t_L g1047 ( .A(n_945), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_922), .A2(n_1004), .B1(n_929), .B2(n_920), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_924), .Y(n_1049) );
AOI221xp5_ASAP7_75t_L g1050 ( .A1(n_933), .A2(n_955), .B1(n_959), .B2(n_995), .C(n_932), .Y(n_1050) );
INVx2_ASAP7_75t_L g1051 ( .A(n_942), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_924), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_925), .B(n_927), .Y(n_1053) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_925), .B(n_927), .Y(n_1054) );
OAI21xp5_ASAP7_75t_L g1055 ( .A1(n_931), .A2(n_992), .B(n_994), .Y(n_1055) );
NOR3xp33_ASAP7_75t_L g1056 ( .A(n_993), .B(n_955), .C(n_999), .Y(n_1056) );
BUFx2_ASAP7_75t_L g1057 ( .A(n_958), .Y(n_1057) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_936), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_964), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_964), .B(n_996), .Y(n_1060) );
BUFx2_ASAP7_75t_L g1061 ( .A(n_1001), .Y(n_1061) );
AOI21x1_ASAP7_75t_L g1062 ( .A1(n_923), .A2(n_962), .B(n_966), .Y(n_1062) );
INVx2_ASAP7_75t_L g1063 ( .A(n_923), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_966), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_981), .Y(n_1065) );
AO21x2_ASAP7_75t_L g1066 ( .A1(n_970), .A2(n_976), .B(n_981), .Y(n_1066) );
AOI33xp33_ASAP7_75t_L g1067 ( .A1(n_974), .A2(n_980), .A3(n_985), .B1(n_983), .B2(n_973), .B3(n_961), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_996), .B(n_941), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_974), .A2(n_983), .B1(n_986), .B2(n_998), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_941), .B(n_923), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1000), .B(n_969), .Y(n_1071) );
OR2x6_ASAP7_75t_L g1072 ( .A(n_991), .B(n_982), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_970), .Y(n_1073) );
HB1xp67_ASAP7_75t_L g1074 ( .A(n_947), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1000), .B(n_970), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1038), .B(n_991), .Y(n_1076) );
INVx1_ASAP7_75t_SL g1077 ( .A(n_1034), .Y(n_1077) );
OR2x2_ASAP7_75t_L g1078 ( .A(n_1045), .B(n_1058), .Y(n_1078) );
INVx2_ASAP7_75t_L g1079 ( .A(n_1054), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1046), .B(n_971), .Y(n_1080) );
INVx2_ASAP7_75t_SL g1081 ( .A(n_1074), .Y(n_1081) );
NAND3xp33_ASAP7_75t_L g1082 ( .A(n_1048), .B(n_988), .C(n_1002), .Y(n_1082) );
NAND2x1_ASAP7_75t_L g1083 ( .A(n_1071), .B(n_967), .Y(n_1083) );
AND2x2_ASAP7_75t_SL g1084 ( .A(n_1071), .B(n_965), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1021), .B(n_954), .Y(n_1085) );
HB1xp67_ASAP7_75t_L g1086 ( .A(n_1006), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_1035), .B(n_1043), .Y(n_1087) );
NOR2x1_ASAP7_75t_SL g1088 ( .A(n_1072), .B(n_1005), .Y(n_1088) );
OAI31xp33_ASAP7_75t_SL g1089 ( .A1(n_1041), .A2(n_990), .A3(n_972), .B(n_926), .Y(n_1089) );
AND2x4_ASAP7_75t_L g1090 ( .A(n_1024), .B(n_1010), .Y(n_1090) );
HB1xp67_ASAP7_75t_L g1091 ( .A(n_1006), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1068), .B(n_1010), .Y(n_1092) );
NOR2xp33_ASAP7_75t_L g1093 ( .A(n_1041), .B(n_1042), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1043), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1049), .Y(n_1095) );
OAI21xp5_ASAP7_75t_SL g1096 ( .A1(n_1056), .A2(n_1050), .B(n_1069), .Y(n_1096) );
INVx1_ASAP7_75t_SL g1097 ( .A(n_1068), .Y(n_1097) );
INVx3_ASAP7_75t_SL g1098 ( .A(n_1072), .Y(n_1098) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1006), .Y(n_1099) );
INVxp67_ASAP7_75t_L g1100 ( .A(n_1032), .Y(n_1100) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_1018), .Y(n_1101) );
AOI331xp33_ASAP7_75t_L g1102 ( .A1(n_1030), .A2(n_1008), .A3(n_1019), .B1(n_1022), .B2(n_1032), .B3(n_1036), .C1(n_1052), .Y(n_1102) );
OR2x6_ASAP7_75t_L g1103 ( .A(n_1072), .B(n_1061), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1012), .B(n_1070), .Y(n_1104) );
A2O1A1Ixp33_ASAP7_75t_L g1105 ( .A1(n_1067), .A2(n_1017), .B(n_1031), .C(n_1040), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1106 ( .A(n_1053), .B(n_1014), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1012), .B(n_1070), .Y(n_1107) );
NAND2x1p5_ASAP7_75t_L g1108 ( .A(n_1044), .B(n_1061), .Y(n_1108) );
OR2x6_ASAP7_75t_L g1109 ( .A(n_1072), .B(n_1009), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1049), .Y(n_1110) );
NOR2xp33_ASAP7_75t_L g1111 ( .A(n_1028), .B(n_1027), .Y(n_1111) );
AOI33xp33_ASAP7_75t_L g1112 ( .A1(n_1027), .A2(n_1022), .A3(n_1019), .B1(n_1007), .B2(n_1075), .B3(n_1013), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1053), .B(n_1060), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1114 ( .A(n_1009), .B(n_1059), .Y(n_1114) );
NOR2xp33_ASAP7_75t_L g1115 ( .A(n_1011), .B(n_1037), .Y(n_1115) );
INVx1_ASAP7_75t_SL g1116 ( .A(n_1044), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1059), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1064), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1064), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1060), .B(n_1065), .Y(n_1120) );
AOI221xp5_ASAP7_75t_SL g1121 ( .A1(n_1023), .A2(n_1055), .B1(n_1075), .B2(n_1007), .C(n_1057), .Y(n_1121) );
OR2x2_ASAP7_75t_L g1122 ( .A(n_1065), .B(n_1015), .Y(n_1122) );
AND2x4_ASAP7_75t_SL g1123 ( .A(n_1072), .B(n_1039), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1036), .Y(n_1124) );
OAI31xp33_ASAP7_75t_L g1125 ( .A1(n_1057), .A2(n_1044), .A3(n_1039), .B(n_1026), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1124), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1104), .B(n_1026), .Y(n_1127) );
AND2x4_ASAP7_75t_L g1128 ( .A(n_1123), .B(n_1039), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1111), .B(n_1029), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1107), .B(n_1039), .Y(n_1130) );
OR2x2_ASAP7_75t_L g1131 ( .A(n_1087), .B(n_1063), .Y(n_1131) );
NAND2x1p5_ASAP7_75t_L g1132 ( .A(n_1116), .B(n_1062), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1078), .Y(n_1133) );
NAND4xp75_ASAP7_75t_SL g1134 ( .A(n_1093), .B(n_1062), .C(n_1033), .D(n_1066), .Y(n_1134) );
NOR2xp33_ASAP7_75t_L g1135 ( .A(n_1077), .B(n_1020), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1086), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1086), .Y(n_1137) );
NAND2x1p5_ASAP7_75t_L g1138 ( .A(n_1081), .B(n_1020), .Y(n_1138) );
NOR2xp67_ASAP7_75t_SL g1139 ( .A(n_1096), .B(n_1020), .Y(n_1139) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1099), .Y(n_1140) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1099), .Y(n_1141) );
NAND4xp75_ASAP7_75t_L g1142 ( .A(n_1084), .B(n_1047), .C(n_1073), .D(n_1051), .Y(n_1142) );
NOR2xp33_ASAP7_75t_L g1143 ( .A(n_1085), .B(n_1066), .Y(n_1143) );
HB1xp67_ASAP7_75t_L g1144 ( .A(n_1097), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1113), .B(n_1025), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1092), .B(n_1025), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1120), .B(n_1025), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1094), .B(n_1106), .Y(n_1148) );
OR2x2_ASAP7_75t_L g1149 ( .A(n_1114), .B(n_1051), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1091), .Y(n_1150) );
XOR2x2_ASAP7_75t_L g1151 ( .A(n_1083), .B(n_1016), .Y(n_1151) );
INVx3_ASAP7_75t_L g1152 ( .A(n_1123), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1079), .B(n_1102), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1136), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1146), .B(n_1109), .Y(n_1155) );
BUFx3_ASAP7_75t_L g1156 ( .A(n_1138), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1146), .B(n_1098), .Y(n_1157) );
NAND2xp5_ASAP7_75t_SL g1158 ( .A(n_1151), .B(n_1121), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1144), .B(n_1122), .Y(n_1159) );
NOR2x1_ASAP7_75t_L g1160 ( .A(n_1152), .B(n_1105), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1136), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1137), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1137), .Y(n_1163) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1140), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1145), .B(n_1098), .Y(n_1165) );
NOR2xp67_ASAP7_75t_SL g1166 ( .A(n_1152), .B(n_1076), .Y(n_1166) );
AOI211xp5_ASAP7_75t_L g1167 ( .A1(n_1139), .A2(n_1115), .B(n_1082), .C(n_1089), .Y(n_1167) );
AOI221xp5_ASAP7_75t_L g1168 ( .A1(n_1139), .A2(n_1115), .B1(n_1080), .B2(n_1100), .C(n_1125), .Y(n_1168) );
AOI22xp5_ASAP7_75t_L g1169 ( .A1(n_1142), .A2(n_1103), .B1(n_1090), .B2(n_1100), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1126), .Y(n_1170) );
NOR2x1_ASAP7_75t_L g1171 ( .A(n_1152), .B(n_1103), .Y(n_1171) );
OAI21xp33_ASAP7_75t_L g1172 ( .A1(n_1143), .A2(n_1112), .B(n_1103), .Y(n_1172) );
AOI21xp5_ASAP7_75t_L g1173 ( .A1(n_1151), .A2(n_1088), .B(n_1108), .Y(n_1173) );
NAND2xp33_ASAP7_75t_L g1174 ( .A(n_1142), .B(n_1108), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1129), .B(n_1118), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1145), .B(n_1091), .Y(n_1176) );
XOR2x2_ASAP7_75t_L g1177 ( .A(n_1133), .B(n_1090), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1126), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1127), .B(n_1101), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1131), .Y(n_1180) );
O2A1O1Ixp33_ASAP7_75t_L g1181 ( .A1(n_1153), .A2(n_1119), .B(n_1117), .C(n_1110), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1131), .Y(n_1182) );
XOR2x2_ASAP7_75t_L g1183 ( .A(n_1148), .B(n_1095), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1127), .B(n_1101), .Y(n_1184) );
OAI21xp5_ASAP7_75t_L g1185 ( .A1(n_1135), .A2(n_1016), .B(n_1138), .Y(n_1185) );
NOR2xp33_ASAP7_75t_L g1186 ( .A(n_1130), .B(n_1147), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1150), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1150), .Y(n_1188) );
AOI21xp5_ASAP7_75t_L g1189 ( .A1(n_1138), .A2(n_1128), .B(n_1132), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1149), .Y(n_1190) );
AOI21xp5_ASAP7_75t_L g1191 ( .A1(n_1158), .A2(n_1160), .B(n_1173), .Y(n_1191) );
OAI211xp5_ASAP7_75t_L g1192 ( .A1(n_1167), .A2(n_1168), .B(n_1172), .C(n_1181), .Y(n_1192) );
AO21x1_ASAP7_75t_L g1193 ( .A1(n_1189), .A2(n_1174), .B(n_1185), .Y(n_1193) );
NOR2x1_ASAP7_75t_L g1194 ( .A(n_1171), .B(n_1174), .Y(n_1194) );
OAI21xp33_ASAP7_75t_SL g1195 ( .A1(n_1186), .A2(n_1169), .B(n_1183), .Y(n_1195) );
INVx2_ASAP7_75t_SL g1196 ( .A(n_1177), .Y(n_1196) );
OAI21xp5_ASAP7_75t_L g1197 ( .A1(n_1177), .A2(n_1159), .B(n_1186), .Y(n_1197) );
NOR2xp67_ASAP7_75t_L g1198 ( .A(n_1156), .B(n_1157), .Y(n_1198) );
OAI211xp5_ASAP7_75t_SL g1199 ( .A1(n_1191), .A2(n_1159), .B(n_1182), .C(n_1180), .Y(n_1199) );
NOR3xp33_ASAP7_75t_SL g1200 ( .A(n_1192), .B(n_1175), .C(n_1161), .Y(n_1200) );
O2A1O1Ixp33_ASAP7_75t_L g1201 ( .A1(n_1195), .A2(n_1132), .B(n_1162), .C(n_1154), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1196), .Y(n_1202) );
HB1xp67_ASAP7_75t_L g1203 ( .A(n_1198), .Y(n_1203) );
NAND2xp33_ASAP7_75t_SL g1204 ( .A(n_1197), .B(n_1166), .Y(n_1204) );
OAI211xp5_ASAP7_75t_L g1205 ( .A1(n_1194), .A2(n_1155), .B(n_1157), .C(n_1165), .Y(n_1205) );
AND3x4_ASAP7_75t_L g1206 ( .A(n_1200), .B(n_1193), .C(n_1156), .Y(n_1206) );
NOR2xp67_ASAP7_75t_L g1207 ( .A(n_1205), .B(n_1163), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1202), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_1204), .A2(n_1166), .B1(n_1155), .B2(n_1128), .Y(n_1209) );
OAI222xp33_ASAP7_75t_L g1210 ( .A1(n_1201), .A2(n_1165), .B1(n_1190), .B2(n_1188), .C1(n_1187), .C2(n_1132), .Y(n_1210) );
OR4x2_ASAP7_75t_L g1211 ( .A(n_1206), .B(n_1204), .C(n_1199), .D(n_1203), .Y(n_1211) );
NOR3xp33_ASAP7_75t_L g1212 ( .A(n_1208), .B(n_1178), .C(n_1170), .Y(n_1212) );
INVx2_ASAP7_75t_L g1213 ( .A(n_1207), .Y(n_1213) );
OAI21xp5_ASAP7_75t_L g1214 ( .A1(n_1213), .A2(n_1209), .B(n_1210), .Y(n_1214) );
XNOR2xp5_ASAP7_75t_L g1215 ( .A(n_1211), .B(n_1134), .Y(n_1215) );
OAI22xp5_ASAP7_75t_SL g1216 ( .A1(n_1212), .A2(n_1128), .B1(n_1164), .B2(n_1141), .Y(n_1216) );
XNOR2xp5_ASAP7_75t_L g1217 ( .A(n_1215), .B(n_1179), .Y(n_1217) );
OAI22x1_ASAP7_75t_L g1218 ( .A1(n_1214), .A2(n_1179), .B1(n_1184), .B2(n_1176), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1216), .Y(n_1219) );
HB1xp67_ASAP7_75t_L g1220 ( .A(n_1219), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1217), .Y(n_1221) );
INVx4_ASAP7_75t_L g1222 ( .A(n_1218), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1221), .Y(n_1223) );
AOI21xp5_ASAP7_75t_L g1224 ( .A1(n_1223), .A2(n_1220), .B(n_1222), .Y(n_1224) );
endmodule