module fake_jpeg_30521_n_354 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_354);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_354;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_1),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_1),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_16),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_55),
.A2(n_18),
.B1(n_35),
.B2(n_25),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_63),
.A2(n_64),
.B1(n_70),
.B2(n_87),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_18),
.B1(n_35),
.B2(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_77),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_26),
.B1(n_25),
.B2(n_20),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_28),
.B1(n_38),
.B2(n_21),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_71),
.A2(n_40),
.B1(n_3),
.B2(n_4),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_52),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_94),
.Y(n_114)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_102),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_41),
.B(n_38),
.Y(n_94)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_95),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_16),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_100),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_47),
.A2(n_32),
.B1(n_33),
.B2(n_31),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_130)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_23),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_13),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_31),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_104),
.Y(n_174)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_39),
.B(n_17),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_109),
.C(n_129),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_21),
.B(n_23),
.C(n_32),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_107),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_32),
.C(n_39),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_39),
.B1(n_17),
.B2(n_15),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_17),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_122),
.Y(n_144)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_17),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_50),
.B1(n_42),
.B2(n_40),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_127),
.B1(n_74),
.B2(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_1),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_86),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_85),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_2),
.C(n_3),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_112),
.B1(n_121),
.B2(n_107),
.Y(n_153)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_133),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_88),
.A2(n_73),
.B1(n_79),
.B2(n_93),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_89),
.Y(n_145)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_135),
.Y(n_143)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_83),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_137),
.Y(n_146)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_82),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_96),
.B1(n_66),
.B2(n_90),
.Y(n_159)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_5),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_158),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_150),
.A2(n_108),
.B1(n_119),
.B2(n_131),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_153),
.A2(n_156),
.B1(n_160),
.B2(n_150),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_73),
.B1(n_88),
.B2(n_93),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_172),
.B1(n_178),
.B2(n_179),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_110),
.A2(n_109),
.B(n_106),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_155),
.B(n_162),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_82),
.B1(n_67),
.B2(n_96),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_110),
.B(n_67),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_159),
.A2(n_168),
.B1(n_177),
.B2(n_174),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_115),
.A2(n_68),
.B1(n_95),
.B2(n_74),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_90),
.Y(n_162)
);

AO22x2_ASAP7_75t_L g163 ( 
.A1(n_104),
.A2(n_68),
.B1(n_6),
.B2(n_7),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_163),
.B(n_175),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_170),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_114),
.A2(n_118),
.B1(n_126),
.B2(n_139),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_12),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_119),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_135),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_108),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_117),
.C(n_113),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_103),
.A2(n_137),
.B1(n_120),
.B2(n_105),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_118),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_200),
.B1(n_214),
.B2(n_161),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_146),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_197),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_189),
.B(n_199),
.Y(n_228)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_158),
.B(n_144),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_194),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_133),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_151),
.A2(n_125),
.B(n_141),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_171),
.B(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_143),
.B(n_125),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_11),
.B1(n_170),
.B2(n_145),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_198),
.A2(n_205),
.B1(n_212),
.B2(n_180),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_147),
.B(n_11),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_203),
.Y(n_229)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_149),
.B(n_175),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_165),
.B(n_169),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_207),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_145),
.A2(n_156),
.B1(n_159),
.B2(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_210),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_155),
.B(n_160),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_173),
.B(n_157),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_215),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_152),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_152),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_213),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_163),
.B(n_176),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_151),
.A2(n_157),
.B1(n_163),
.B2(n_161),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_216),
.A2(n_235),
.B1(n_219),
.B2(n_227),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_163),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_228),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_207),
.A2(n_142),
.B(n_171),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_238),
.B(n_189),
.C(n_188),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_171),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_236),
.C(n_240),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_213),
.B1(n_214),
.B2(n_185),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_226),
.A2(n_235),
.B1(n_217),
.B2(n_240),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_210),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_239),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_183),
.C(n_206),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_SL g238 ( 
.A(n_204),
.B(n_180),
.C(n_209),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_193),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_185),
.B(n_192),
.C(n_188),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_195),
.A2(n_211),
.B(n_198),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_242),
.A2(n_195),
.B(n_194),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_181),
.B1(n_197),
.B2(n_212),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_219),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_245),
.Y(n_284)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_247),
.A2(n_237),
.B(n_241),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_238),
.A2(n_187),
.B1(n_182),
.B2(n_184),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_248),
.A2(n_250),
.B(n_253),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_244),
.A2(n_186),
.B1(n_181),
.B2(n_205),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_252),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_223),
.B1(n_216),
.B2(n_226),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_191),
.B1(n_196),
.B2(n_201),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_261),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_202),
.C(n_208),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_259),
.C(n_255),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_215),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_232),
.A2(n_239),
.B1(n_230),
.B2(n_218),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_222),
.B(n_234),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_224),
.B1(n_220),
.B2(n_217),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_220),
.Y(n_262)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_263),
.A2(n_264),
.B1(n_259),
.B2(n_249),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_233),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_265),
.B(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_228),
.B(n_229),
.Y(n_267)
);

AOI22x1_ASAP7_75t_L g268 ( 
.A1(n_221),
.A2(n_227),
.B1(n_233),
.B2(n_243),
.Y(n_268)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_225),
.A2(n_231),
.B1(n_234),
.B2(n_237),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_225),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_274),
.A2(n_279),
.B(n_253),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_257),
.B(n_222),
.Y(n_278)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_269),
.Y(n_302)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_241),
.Y(n_283)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_257),
.B(n_243),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_256),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_255),
.C(n_258),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_288),
.B(n_252),
.Y(n_290)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_290),
.B(n_291),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_289),
.A2(n_249),
.B(n_247),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_287),
.C(n_281),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_284),
.B(n_263),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_302),
.Y(n_312)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_286),
.B1(n_275),
.B2(n_250),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_296),
.A2(n_300),
.B1(n_303),
.B2(n_270),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_251),
.B1(n_268),
.B2(n_261),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_275),
.A2(n_279),
.B(n_273),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_270),
.Y(n_319)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_284),
.Y(n_305)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_308),
.C(n_313),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_288),
.C(n_248),
.Y(n_308)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_282),
.C(n_273),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_303),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_268),
.C(n_274),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_278),
.C(n_283),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_298),
.C(n_299),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_276),
.Y(n_329)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_297),
.Y(n_317)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_318),
.A2(n_299),
.B1(n_306),
.B2(n_296),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_304),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_326),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_322),
.B(n_312),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_307),
.B(n_314),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_309),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_313),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_329),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_325),
.A2(n_310),
.B1(n_306),
.B2(n_315),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_332),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g332 ( 
.A(n_326),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_336),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_325),
.A2(n_311),
.B1(n_308),
.B2(n_300),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_321),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_276),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_338),
.A2(n_301),
.B(n_272),
.Y(n_343)
);

AOI31xp33_ASAP7_75t_L g340 ( 
.A1(n_332),
.A2(n_323),
.A3(n_320),
.B(n_321),
.Y(n_340)
);

OAI21x1_ASAP7_75t_L g345 ( 
.A1(n_340),
.A2(n_337),
.B(n_334),
.Y(n_345)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_342),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_343),
.B(n_344),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_295),
.C(n_272),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_345),
.A2(n_347),
.B(n_339),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_341),
.A2(n_335),
.B(n_280),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_349),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_348),
.A2(n_340),
.B1(n_271),
.B2(n_285),
.Y(n_350)
);

FAx1_ASAP7_75t_SL g352 ( 
.A(n_351),
.B(n_350),
.CI(n_346),
.CON(n_352),
.SN(n_352)
);

OAI21x1_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_271),
.B(n_330),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_352),
.Y(n_354)
);


endmodule