module fake_netlist_1_8807_n_14 (n_1, n_2, n_0, n_14);
input n_1;
input n_2;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
NAND2xp33_ASAP7_75t_L g3 ( .A(n_1), .B(n_0), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_4), .Y(n_5) );
AND2x2_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_5), .B(n_3), .Y(n_7) );
AO21x2_ASAP7_75t_L g8 ( .A1(n_6), .A2(n_0), .B(n_1), .Y(n_8) );
NAND3xp33_ASAP7_75t_L g9 ( .A(n_7), .B(n_5), .C(n_6), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
OAI211xp5_ASAP7_75t_SL g11 ( .A1(n_9), .A2(n_7), .B(n_8), .C(n_6), .Y(n_11) );
BUFx2_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
AOI22xp5_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_8), .B1(n_1), .B2(n_2), .Y(n_13) );
AOI22xp5_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_2), .B1(n_12), .B2(n_11), .Y(n_14) );
endmodule