module fake_ariane_1622_n_1967 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1967);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1967;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_181;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g179 ( 
.A(n_23),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_14),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_97),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_41),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_0),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_7),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_76),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_107),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_93),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_136),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_115),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_2),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_82),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_135),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_172),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_118),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_109),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_52),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_62),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_66),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_30),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_103),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_167),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_39),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_119),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_72),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_28),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_158),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_110),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_57),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_47),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_69),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_152),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_2),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_30),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_126),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_68),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_150),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_40),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_79),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_67),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_65),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_85),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_176),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_92),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_98),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_154),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_134),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_59),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_83),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_10),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_14),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_27),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_163),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_18),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_8),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_155),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_20),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_95),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_7),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_21),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_10),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_46),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_61),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_17),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_104),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_111),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_124),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_45),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_122),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_74),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_63),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_168),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_128),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_99),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_18),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_77),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_68),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_87),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_20),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_21),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_78),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_11),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_32),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_39),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_174),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_69),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_116),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_0),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_121),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_15),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_6),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_9),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_170),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_47),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_159),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_42),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_54),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_127),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_59),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_75),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_31),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_35),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_144),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_178),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_52),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_112),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_45),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_153),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_132),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_165),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_113),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_63),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_57),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_41),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_175),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_38),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_56),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_8),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_67),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_12),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_42),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_58),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_86),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_70),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_80),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_62),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_26),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_36),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_148),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_177),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_32),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_129),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_58),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_56),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_55),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_71),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_38),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_34),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_5),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_142),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_31),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_131),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_54),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_17),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_146),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_43),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_65),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_143),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_55),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_88),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_6),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_23),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_9),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_34),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_140),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_29),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_16),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_162),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_114),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_33),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_35),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_145),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_27),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_36),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_100),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_102),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_29),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_61),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_161),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_44),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_191),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_216),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_192),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_226),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_200),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_201),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_226),
.B(n_1),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_226),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_226),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_324),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_216),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_188),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_181),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_181),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_190),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_188),
.Y(n_372)
);

BUFx2_ASAP7_75t_SL g373 ( 
.A(n_188),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_208),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_190),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_195),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_201),
.B(n_1),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_234),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_188),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_324),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_195),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_243),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_243),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_199),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_199),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_350),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_205),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_324),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_342),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_258),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_332),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_332),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_350),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_332),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_335),
.Y(n_397)
);

BUFx6f_ASAP7_75t_SL g398 ( 
.A(n_243),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_186),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_325),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_335),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_322),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_218),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_243),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_179),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_187),
.B(n_3),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_180),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_185),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_194),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_221),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_305),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_179),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_202),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_205),
.B(n_232),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_187),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_244),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_210),
.Y(n_418)
);

NOR2xp67_ASAP7_75t_L g419 ( 
.A(n_214),
.B(n_3),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_204),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_210),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_277),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_338),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_242),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_221),
.Y(n_425)
);

BUFx5_ASAP7_75t_L g426 ( 
.A(n_232),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_305),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_242),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_221),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_213),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_215),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_251),
.B(n_4),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_270),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_217),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_251),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_247),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_220),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_222),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_255),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_255),
.B(n_4),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_247),
.Y(n_441)
);

NOR2xp67_ASAP7_75t_L g442 ( 
.A(n_214),
.B(n_11),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_305),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_224),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_262),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_257),
.B(n_12),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_364),
.B(n_257),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_263),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_427),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_358),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_443),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_427),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_365),
.Y(n_454)
);

OR2x6_ASAP7_75t_L g455 ( 
.A(n_377),
.B(n_262),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_360),
.B(n_263),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_365),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_373),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_411),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_369),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_402),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_369),
.B(n_283),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_370),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_370),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_371),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_371),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_375),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_402),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_402),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_375),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_376),
.B(n_305),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_440),
.A2(n_315),
.B(n_225),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

NOR2x1_ASAP7_75t_L g474 ( 
.A(n_373),
.B(n_270),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_426),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_376),
.B(n_283),
.Y(n_477)
);

NAND2x1_ASAP7_75t_L g478 ( 
.A(n_381),
.B(n_225),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_381),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_384),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_362),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_426),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_426),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_393),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_426),
.Y(n_488)
);

BUFx12f_ASAP7_75t_L g489 ( 
.A(n_372),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_386),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_426),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_426),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_426),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_385),
.B(n_285),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_387),
.B(n_305),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_387),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_435),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_396),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_435),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_399),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_439),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_397),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_401),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_404),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_439),
.B(n_285),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_366),
.B(n_292),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_380),
.B(n_305),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_380),
.B(n_270),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_415),
.B(n_336),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_388),
.B(n_389),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_363),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_446),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_406),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_413),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_421),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_395),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_445),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_424),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_357),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_400),
.B(n_291),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_441),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_390),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_391),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_368),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_458),
.B(n_358),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_485),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_482),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_485),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_496),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_496),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_449),
.Y(n_532)
);

NOR2x1p5_ASAP7_75t_L g533 ( 
.A(n_489),
.B(n_377),
.Y(n_533)
);

INVxp33_ASAP7_75t_SL g534 ( 
.A(n_450),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_458),
.B(n_372),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_455),
.A2(n_432),
.B1(n_416),
.B2(n_398),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_496),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_496),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_496),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_521),
.B(n_490),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_379),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_459),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_459),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_474),
.B(n_379),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_455),
.A2(n_367),
.B1(n_383),
.B2(n_382),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_492),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_449),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_454),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_457),
.Y(n_550)
);

BUFx8_ASAP7_75t_SL g551 ( 
.A(n_500),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_449),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_457),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_455),
.A2(n_416),
.B1(n_398),
.B2(n_425),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_460),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_492),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_452),
.Y(n_557)
);

BUFx4f_ASAP7_75t_L g558 ( 
.A(n_512),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_512),
.B(n_225),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_459),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_460),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_455),
.A2(n_398),
.B1(n_433),
.B2(n_429),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_452),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_485),
.Y(n_564)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_455),
.A2(n_367),
.B1(n_521),
.B2(n_383),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_455),
.A2(n_405),
.B1(n_382),
.B2(n_408),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_500),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_447),
.B(n_405),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_509),
.B(n_408),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_447),
.B(n_409),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_509),
.B(n_409),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_485),
.Y(n_572)
);

INVx5_ASAP7_75t_L g573 ( 
.A(n_482),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_452),
.Y(n_574)
);

OR2x6_ASAP7_75t_L g575 ( 
.A(n_455),
.B(n_407),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_485),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_508),
.A2(n_474),
.B1(n_489),
.B2(n_509),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_509),
.B(n_414),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_509),
.A2(n_442),
.B1(n_419),
.B2(n_306),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_451),
.B(n_414),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_463),
.Y(n_581)
);

BUFx10_ASAP7_75t_L g582 ( 
.A(n_508),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_463),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_451),
.B(n_512),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_508),
.A2(n_306),
.B1(n_291),
.B2(n_271),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_512),
.B(n_420),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_464),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_521),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_464),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_512),
.B(n_420),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_507),
.B(n_428),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_485),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_508),
.A2(n_327),
.B1(n_300),
.B2(n_271),
.Y(n_593)
);

CKINVDCx11_ASAP7_75t_R g594 ( 
.A(n_489),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_512),
.B(n_430),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_490),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_492),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_485),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_465),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_485),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_486),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_520),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_512),
.B(n_430),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_486),
.Y(n_604)
);

AND2x2_ASAP7_75t_SL g605 ( 
.A(n_450),
.B(n_315),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_465),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_513),
.B(n_515),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_486),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_466),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_512),
.B(n_431),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_466),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_467),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_486),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_450),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_492),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_482),
.Y(n_616)
);

AO22x2_ASAP7_75t_L g617 ( 
.A1(n_478),
.A2(n_339),
.B1(n_203),
.B2(n_315),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_507),
.B(n_431),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_482),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_508),
.B(n_434),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_481),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_467),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_506),
.B(n_434),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_507),
.A2(n_524),
.B1(n_506),
.B2(n_515),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_486),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_507),
.A2(n_524),
.B1(n_516),
.B2(n_519),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_507),
.B(n_470),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_523),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_470),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_486),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_479),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_486),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_479),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_480),
.B(n_437),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_480),
.B(n_437),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_484),
.B(n_487),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_484),
.B(n_444),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_487),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_497),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_497),
.B(n_444),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_499),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_499),
.B(n_410),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_448),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_482),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_501),
.B(n_438),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_486),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_501),
.B(n_448),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_502),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_514),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_514),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_481),
.A2(n_436),
.B1(n_260),
.B2(n_308),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_513),
.A2(n_516),
.B1(n_519),
.B2(n_518),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_517),
.B(n_359),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_502),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_502),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_514),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_502),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_518),
.B(n_325),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_517),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_502),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_514),
.B(n_325),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_514),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_523),
.B(n_183),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_483),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_523),
.B(n_310),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_523),
.B(n_292),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_523),
.B(n_483),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_502),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_514),
.Y(n_669)
);

INVx5_ASAP7_75t_L g670 ( 
.A(n_483),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_471),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_514),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_514),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_471),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_483),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_502),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_502),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_605),
.B(n_483),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_544),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_540),
.B(n_614),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_544),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_568),
.B(n_462),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_532),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_532),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_549),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_596),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_596),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_549),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_570),
.B(n_462),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_541),
.B(n_361),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_623),
.B(n_374),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_580),
.B(n_477),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_SL g693 ( 
.A(n_605),
.B(n_378),
.Y(n_693)
);

AO22x2_ASAP7_75t_L g694 ( 
.A1(n_658),
.A2(n_478),
.B1(n_279),
.B2(n_284),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_658),
.B(n_477),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_534),
.B(n_392),
.Y(n_696)
);

NOR3xp33_ASAP7_75t_L g697 ( 
.A(n_565),
.B(n_207),
.C(n_275),
.Y(n_697)
);

O2A1O1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_627),
.A2(n_456),
.B(n_505),
.C(n_494),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_548),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_628),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_617),
.A2(n_478),
.B1(n_518),
.B2(n_522),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_550),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_548),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_552),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_550),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_586),
.B(n_494),
.Y(n_706)
);

AND2x6_ASAP7_75t_SL g707 ( 
.A(n_551),
.B(n_275),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_610),
.B(n_505),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_540),
.B(n_510),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_628),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_635),
.B(n_491),
.Y(n_711)
);

AOI21x1_ASAP7_75t_L g712 ( 
.A1(n_667),
.A2(n_472),
.B(n_475),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_552),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_620),
.A2(n_522),
.B1(n_229),
.B2(n_510),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_553),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_572),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_553),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_617),
.A2(n_522),
.B1(n_471),
.B2(n_495),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_575),
.B(n_471),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_582),
.B(n_491),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_637),
.A2(n_522),
.B1(n_456),
.B2(n_471),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_557),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_557),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_555),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_647),
.B(n_491),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_525),
.B(n_491),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_526),
.B(n_491),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_563),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_582),
.B(n_475),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_534),
.B(n_403),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_563),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_582),
.B(n_475),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_558),
.B(n_616),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_528),
.B(n_476),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_558),
.B(n_616),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_588),
.B(n_417),
.Y(n_736)
);

AND2x2_ASAP7_75t_SL g737 ( 
.A(n_536),
.B(n_344),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_624),
.B(n_522),
.Y(n_738)
);

NOR3xp33_ASAP7_75t_L g739 ( 
.A(n_535),
.B(n_284),
.C(n_279),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_674),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_607),
.B(n_591),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_567),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_574),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_555),
.Y(n_744)
);

AND2x2_ASAP7_75t_SL g745 ( 
.A(n_562),
.B(n_344),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_588),
.B(n_422),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_607),
.B(n_522),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_561),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_659),
.B(n_423),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_L g750 ( 
.A1(n_675),
.A2(n_472),
.B(n_476),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_558),
.B(n_476),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_566),
.B(n_522),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_616),
.B(n_488),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_643),
.B(n_522),
.Y(n_754)
);

INVx5_ASAP7_75t_L g755 ( 
.A(n_559),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_591),
.B(n_634),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_574),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_561),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_575),
.A2(n_495),
.B1(n_294),
.B2(n_295),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_542),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_643),
.B(n_488),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_591),
.B(n_495),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_640),
.B(n_495),
.Y(n_763)
);

BUFx6f_ASAP7_75t_SL g764 ( 
.A(n_575),
.Y(n_764)
);

INVx5_ASAP7_75t_L g765 ( 
.A(n_559),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_619),
.B(n_488),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_542),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_619),
.B(n_493),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_674),
.Y(n_769)
);

BUFx8_ASAP7_75t_L g770 ( 
.A(n_671),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_581),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_584),
.B(n_495),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_643),
.B(n_493),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_602),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_581),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_530),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_626),
.B(n_493),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_618),
.B(n_233),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_590),
.B(n_498),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_530),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_595),
.B(n_498),
.Y(n_781)
);

NAND3xp33_ASAP7_75t_L g782 ( 
.A(n_603),
.B(n_236),
.C(n_235),
.Y(n_782)
);

AND2x4_ASAP7_75t_SL g783 ( 
.A(n_575),
.B(n_325),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_583),
.Y(n_784)
);

INVx8_ASAP7_75t_L g785 ( 
.A(n_559),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_619),
.B(n_472),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_583),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_674),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_L g789 ( 
.A(n_528),
.B(n_237),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_L g790 ( 
.A(n_528),
.B(n_239),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_531),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_671),
.B(n_498),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_531),
.Y(n_793)
);

NOR3xp33_ASAP7_75t_L g794 ( 
.A(n_569),
.B(n_298),
.C(n_290),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_652),
.B(n_503),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_587),
.B(n_503),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_644),
.B(n_294),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_587),
.Y(n_798)
);

NAND2x1_ASAP7_75t_L g799 ( 
.A(n_547),
.B(n_468),
.Y(n_799)
);

AOI221xp5_ASAP7_75t_L g800 ( 
.A1(n_651),
.A2(n_290),
.B1(n_298),
.B2(n_299),
.C(n_300),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_537),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_589),
.B(n_503),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_571),
.B(n_578),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_617),
.A2(n_504),
.B1(n_336),
.B2(n_344),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_547),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_546),
.A2(n_253),
.B1(n_356),
.B2(n_354),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_545),
.B(n_240),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_543),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_644),
.B(n_664),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_537),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_589),
.B(n_504),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_599),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_594),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_599),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_606),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_547),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_538),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_606),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_609),
.B(n_504),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_621),
.B(n_642),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_645),
.B(n_577),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_609),
.B(n_611),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_585),
.B(n_299),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_611),
.B(n_295),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_612),
.B(n_622),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_538),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_593),
.B(n_317),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_612),
.B(n_309),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_602),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_527),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_622),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_629),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_629),
.B(n_631),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_554),
.B(n_245),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_631),
.B(n_309),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_653),
.Y(n_836)
);

OAI21xp33_ASAP7_75t_L g837 ( 
.A1(n_663),
.A2(n_248),
.B(n_246),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_539),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_665),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_543),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_527),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_644),
.B(n_318),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_664),
.B(n_318),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_533),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_617),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_633),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_560),
.B(n_249),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_664),
.B(n_345),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_633),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_742),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_680),
.B(n_533),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_680),
.B(n_579),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_750),
.A2(n_539),
.B(n_649),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_706),
.A2(n_597),
.B(n_556),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_686),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_692),
.A2(n_638),
.B(n_639),
.C(n_641),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_689),
.B(n_638),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_708),
.A2(n_597),
.B(n_556),
.Y(n_858)
);

BUFx4f_ASAP7_75t_L g859 ( 
.A(n_774),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_682),
.A2(n_639),
.B1(n_641),
.B2(n_636),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_821),
.A2(n_666),
.B(n_327),
.C(n_346),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_740),
.B(n_556),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_786),
.A2(n_650),
.B(n_649),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_803),
.A2(n_317),
.B(n_343),
.C(n_353),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_695),
.B(n_560),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_839),
.B(n_528),
.Y(n_866)
);

OAI321xp33_ASAP7_75t_L g867 ( 
.A1(n_691),
.A2(n_834),
.A3(n_800),
.B1(n_806),
.B2(n_804),
.C(n_837),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_756),
.B(n_528),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_786),
.A2(n_656),
.B(n_650),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_741),
.A2(n_346),
.B(n_343),
.C(n_349),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_740),
.B(n_597),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_760),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_760),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_809),
.A2(n_615),
.B(n_573),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_687),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_769),
.B(n_615),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_829),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_809),
.A2(n_615),
.B(n_573),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_683),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_736),
.B(n_347),
.Y(n_880)
);

NAND2x1p5_ASAP7_75t_L g881 ( 
.A(n_788),
.B(n_572),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_769),
.B(n_573),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_725),
.A2(n_670),
.B(n_573),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_753),
.A2(n_670),
.B(n_573),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_679),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_683),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_678),
.B(n_670),
.Y(n_887)
);

AOI21x1_ASAP7_75t_L g888 ( 
.A1(n_751),
.A2(n_662),
.B(n_656),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_822),
.A2(n_670),
.B1(n_600),
.B2(n_601),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_L g890 ( 
.A(n_730),
.B(n_349),
.C(n_347),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_753),
.A2(n_670),
.B(n_669),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_684),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_766),
.A2(n_669),
.B(n_662),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_792),
.B(n_559),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_766),
.A2(n_673),
.B(n_672),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_746),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_770),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_770),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_678),
.B(n_527),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_690),
.A2(n_693),
.B1(n_697),
.B2(n_737),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_684),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_737),
.A2(n_778),
.B1(n_847),
.B2(n_745),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_745),
.A2(n_661),
.B1(n_559),
.B2(n_673),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_768),
.A2(n_672),
.B(n_600),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_699),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_768),
.A2(n_735),
.B(n_733),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_699),
.Y(n_907)
);

INVx1_ASAP7_75t_SL g908 ( 
.A(n_749),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_SL g909 ( 
.A1(n_733),
.A2(n_345),
.B(n_353),
.C(n_668),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_805),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_827),
.A2(n_823),
.B1(n_845),
.B2(n_795),
.Y(n_911)
);

OAI21xp33_ASAP7_75t_L g912 ( 
.A1(n_696),
.A2(n_264),
.B(n_256),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_788),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_681),
.Y(n_914)
);

AND2x6_ASAP7_75t_L g915 ( 
.A(n_719),
.B(n_576),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_792),
.B(n_559),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_761),
.B(n_527),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_735),
.A2(n_600),
.B(n_572),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_825),
.A2(n_833),
.B1(n_688),
.B2(n_702),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_685),
.Y(n_920)
);

O2A1O1Ixp5_ASAP7_75t_L g921 ( 
.A1(n_754),
.A2(n_601),
.B(n_646),
.C(n_657),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_727),
.A2(n_646),
.B(n_601),
.Y(n_922)
);

AOI21x1_ASAP7_75t_L g923 ( 
.A1(n_751),
.A2(n_592),
.B(n_576),
.Y(n_923)
);

AO21x1_ASAP7_75t_L g924 ( 
.A1(n_752),
.A2(n_598),
.B(n_592),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_709),
.B(n_559),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_726),
.A2(n_657),
.B(n_646),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_705),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_820),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_763),
.B(n_657),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_805),
.B(n_527),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_715),
.A2(n_677),
.B1(n_676),
.B2(n_668),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_762),
.B(n_717),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_734),
.A2(n_604),
.B(n_598),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_734),
.A2(n_608),
.B(n_604),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_724),
.B(n_608),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_711),
.A2(n_625),
.B(n_613),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_744),
.B(n_748),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_836),
.B(n_265),
.Y(n_938)
);

INVx4_ASAP7_75t_L g939 ( 
.A(n_785),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_827),
.B(n_267),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_773),
.A2(n_625),
.B(n_613),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_758),
.B(n_677),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_698),
.A2(n_676),
.B(n_655),
.C(n_654),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_779),
.A2(n_632),
.B(n_630),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_771),
.B(n_630),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_823),
.B(n_268),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_703),
.Y(n_947)
);

BUFx12f_ASAP7_75t_L g948 ( 
.A(n_813),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_703),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_770),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_805),
.B(n_529),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_775),
.B(n_632),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_704),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_781),
.A2(n_654),
.B(n_648),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_784),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_720),
.A2(n_655),
.B(n_648),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_783),
.B(n_660),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_719),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_787),
.B(n_529),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_704),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_713),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_720),
.A2(n_564),
.B(n_529),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_798),
.B(n_812),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_814),
.A2(n_564),
.B1(n_529),
.B2(n_660),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_815),
.B(n_529),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_818),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_797),
.A2(n_660),
.B(n_564),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_816),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_831),
.B(n_564),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_832),
.B(n_564),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_783),
.B(n_660),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_846),
.B(n_660),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_795),
.A2(n_336),
.B1(n_273),
.B2(n_276),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_797),
.A2(n_468),
.B(n_453),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_849),
.B(n_269),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_719),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_842),
.A2(n_468),
.B(n_453),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_764),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_842),
.A2(n_468),
.B(n_453),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_764),
.Y(n_980)
);

AOI21x1_ASAP7_75t_L g981 ( 
.A1(n_712),
.A2(n_469),
.B(n_468),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_843),
.A2(n_469),
.B(n_212),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_843),
.A2(n_469),
.B(n_211),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_848),
.A2(n_209),
.B(n_355),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_694),
.B(n_281),
.Y(n_985)
);

AO21x1_ASAP7_75t_L g986 ( 
.A1(n_738),
.A2(n_322),
.B(n_173),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_694),
.B(n_282),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_848),
.A2(n_206),
.B(n_352),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_777),
.A2(n_473),
.B(n_461),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_844),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_SL g991 ( 
.A1(n_813),
.A2(n_286),
.B1(n_287),
.B2(n_293),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_721),
.A2(n_302),
.B(n_303),
.C(n_304),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_816),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_694),
.B(n_794),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_772),
.B(n_307),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_808),
.B(n_312),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_729),
.A2(n_189),
.B(n_351),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_807),
.B(n_313),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_808),
.B(n_314),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_776),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_729),
.A2(n_182),
.B(n_348),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_816),
.B(n_461),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_840),
.B(n_319),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_840),
.B(n_320),
.Y(n_1004)
);

BUFx8_ASAP7_75t_SL g1005 ( 
.A(n_764),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_747),
.B(n_321),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_700),
.B(n_323),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_713),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_722),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_732),
.A2(n_802),
.B(n_796),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_760),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_732),
.A2(n_278),
.B(n_193),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_776),
.B(n_780),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_700),
.B(n_329),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_780),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_700),
.A2(n_330),
.B1(n_333),
.B2(n_337),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_791),
.B(n_340),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_710),
.A2(n_266),
.B1(n_196),
.B2(n_341),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_791),
.B(n_184),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_811),
.A2(n_272),
.B(n_198),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_819),
.A2(n_274),
.B(n_219),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_767),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_710),
.B(n_13),
.Y(n_1023)
);

OAI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_824),
.A2(n_331),
.B(n_223),
.Y(n_1024)
);

BUFx8_ASAP7_75t_L g1025 ( 
.A(n_760),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_828),
.A2(n_322),
.B(n_197),
.C(n_334),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_793),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_793),
.A2(n_838),
.B(n_826),
.C(n_817),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_801),
.A2(n_13),
.B(n_15),
.C(n_16),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_801),
.B(n_227),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_810),
.A2(n_288),
.B(n_230),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_810),
.B(n_228),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_817),
.A2(n_289),
.B(n_238),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_826),
.A2(n_296),
.B(n_241),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_838),
.B(n_231),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_716),
.A2(n_301),
.B(n_252),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_714),
.B(n_250),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_835),
.A2(n_322),
.B(n_254),
.C(n_328),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_767),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_718),
.A2(n_322),
.B1(n_259),
.B2(n_326),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_710),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_759),
.A2(n_311),
.B1(n_280),
.B2(n_297),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_722),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_948),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_879),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_857),
.A2(n_789),
.B(n_790),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_915),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_928),
.B(n_716),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_1025),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_885),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_902),
.A2(n_782),
.B1(n_716),
.B2(n_830),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_908),
.B(n_739),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_896),
.B(n_830),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_919),
.B(n_830),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_867),
.B(n_723),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_940),
.B(n_701),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_850),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_854),
.A2(n_790),
.B(n_789),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_943),
.A2(n_799),
.B(n_723),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_900),
.B(n_728),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_875),
.B(n_841),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_998),
.B(n_728),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_858),
.A2(n_841),
.B(n_830),
.Y(n_1063)
);

NOR2xp67_ASAP7_75t_L g1064 ( 
.A(n_978),
.B(n_765),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_914),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_851),
.B(n_841),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_859),
.B(n_841),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_860),
.A2(n_785),
.B(n_731),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_865),
.A2(n_785),
.B(n_731),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_855),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_946),
.B(n_757),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_920),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_998),
.A2(n_743),
.B(n_757),
.C(n_24),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_911),
.B(n_743),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_852),
.B(n_19),
.Y(n_1075)
);

O2A1O1Ixp5_ASAP7_75t_L g1076 ( 
.A1(n_917),
.A2(n_943),
.B(n_951),
.C(n_930),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_872),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_856),
.A2(n_785),
.B(n_765),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_911),
.B(n_880),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_861),
.A2(n_765),
.B(n_755),
.C(n_316),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_890),
.A2(n_19),
.B(n_22),
.C(n_24),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_932),
.B(n_976),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_856),
.A2(n_765),
.B(n_755),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_937),
.A2(n_765),
.B1(n_755),
.B2(n_261),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_879),
.Y(n_1085)
);

AND2x2_ASAP7_75t_SL g1086 ( 
.A(n_1040),
.B(n_322),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_886),
.Y(n_1087)
);

OAI21xp33_ASAP7_75t_L g1088 ( 
.A1(n_912),
.A2(n_22),
.B(n_25),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_886),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_877),
.Y(n_1090)
);

OA22x2_ASAP7_75t_L g1091 ( 
.A1(n_898),
.A2(n_707),
.B1(n_755),
.B2(n_28),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_958),
.B(n_755),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_995),
.B(n_25),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_906),
.A2(n_473),
.B(n_461),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1010),
.A2(n_473),
.B(n_461),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_915),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_963),
.B(n_26),
.Y(n_1097)
);

NOR2x1_ASAP7_75t_L g1098 ( 
.A(n_897),
.B(n_473),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_990),
.B(n_33),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_892),
.Y(n_1100)
);

O2A1O1Ixp5_ASAP7_75t_L g1101 ( 
.A1(n_917),
.A2(n_37),
.B(n_40),
.C(n_43),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1022),
.B(n_37),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_938),
.A2(n_473),
.B1(n_461),
.B2(n_48),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_883),
.A2(n_473),
.B(n_461),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_927),
.B(n_44),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_859),
.B(n_461),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_955),
.B(n_46),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_872),
.Y(n_1108)
);

NAND3xp33_ASAP7_75t_SL g1109 ( 
.A(n_864),
.B(n_48),
.C(n_49),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_892),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_1025),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_1025),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_922),
.A2(n_473),
.B(n_461),
.Y(n_1113)
);

CKINVDCx16_ASAP7_75t_R g1114 ( 
.A(n_948),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_864),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_966),
.B(n_50),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_853),
.A2(n_473),
.B(n_117),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_1039),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_996),
.B(n_51),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_897),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1041),
.B(n_53),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1005),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_861),
.A2(n_53),
.B(n_60),
.C(n_64),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1028),
.A2(n_1007),
.B(n_1014),
.C(n_1023),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_SL g1125 ( 
.A1(n_930),
.A2(n_60),
.B(n_64),
.C(n_66),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_929),
.A2(n_73),
.B(n_81),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_901),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_901),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_973),
.B(n_84),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_926),
.A2(n_89),
.B(n_90),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_973),
.B(n_91),
.Y(n_1131)
);

NAND2x1_ASAP7_75t_L g1132 ( 
.A(n_939),
.B(n_94),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1000),
.B(n_96),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1007),
.A2(n_101),
.B(n_106),
.C(n_108),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1015),
.B(n_120),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_905),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_991),
.B(n_169),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_905),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_999),
.B(n_123),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_1005),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_872),
.Y(n_1141)
);

AO22x1_ASAP7_75t_L g1142 ( 
.A1(n_950),
.A2(n_125),
.B1(n_130),
.B2(n_133),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_964),
.A2(n_137),
.B(n_139),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_1003),
.B(n_1004),
.Y(n_1144)
);

BUFx2_ASAP7_75t_SL g1145 ( 
.A(n_978),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1041),
.B(n_147),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_992),
.A2(n_151),
.B(n_156),
.C(n_157),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_872),
.Y(n_1148)
);

NAND2xp33_ASAP7_75t_L g1149 ( 
.A(n_910),
.B(n_164),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_980),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_975),
.B(n_166),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_913),
.B(n_939),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1014),
.A2(n_1023),
.B(n_992),
.C(n_929),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_873),
.B(n_910),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1026),
.A2(n_1038),
.B(n_1017),
.C(n_1006),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_SL g1156 ( 
.A(n_913),
.B(n_957),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_941),
.A2(n_936),
.B(n_918),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_873),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1027),
.Y(n_1159)
);

NOR2x1_ASAP7_75t_L g1160 ( 
.A(n_1011),
.B(n_957),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_933),
.A2(n_934),
.B(n_1013),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_873),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1026),
.A2(n_1038),
.B(n_1016),
.C(n_1029),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_915),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_915),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_863),
.A2(n_869),
.B(n_944),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_994),
.B(n_915),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_907),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_887),
.B(n_925),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_870),
.A2(n_1033),
.B(n_887),
.C(n_1035),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1040),
.A2(n_965),
.B1(n_970),
.B2(n_972),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_971),
.B(n_866),
.Y(n_1172)
);

AND2x2_ASAP7_75t_SL g1173 ( 
.A(n_939),
.B(n_971),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_868),
.B(n_899),
.Y(n_1174)
);

INVx8_ASAP7_75t_L g1175 ( 
.A(n_873),
.Y(n_1175)
);

INVxp67_ASAP7_75t_SL g1176 ( 
.A(n_894),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_1011),
.Y(n_1177)
);

AOI21x1_ASAP7_75t_L g1178 ( 
.A1(n_989),
.A2(n_981),
.B(n_923),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_968),
.B(n_993),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_954),
.A2(n_956),
.B(n_874),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_L g1181 ( 
.A(n_1024),
.B(n_1042),
.C(n_1018),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_878),
.A2(n_891),
.B(n_904),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_968),
.B(n_993),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_882),
.B(n_951),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_884),
.A2(n_1002),
.B(n_969),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1043),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_916),
.B(n_959),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_881),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_899),
.B(n_985),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_903),
.B(n_889),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1019),
.A2(n_1032),
.B(n_1030),
.C(n_987),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_881),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_984),
.B(n_988),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_947),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_947),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_921),
.A2(n_967),
.B(n_895),
.C(n_893),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_949),
.Y(n_1197)
);

BUFx2_ASAP7_75t_SL g1198 ( 
.A(n_953),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_953),
.B(n_960),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1002),
.A2(n_962),
.B(n_952),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_960),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_961),
.B(n_1009),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_961),
.B(n_1008),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_935),
.B(n_942),
.Y(n_1204)
);

NOR2xp67_ASAP7_75t_SL g1205 ( 
.A(n_882),
.B(n_862),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_931),
.A2(n_945),
.B(n_977),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1178),
.A2(n_888),
.B(n_924),
.Y(n_1207)
);

AO21x1_ASAP7_75t_L g1208 ( 
.A1(n_1062),
.A2(n_862),
.B(n_871),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1159),
.Y(n_1209)
);

AOI221x1_ASAP7_75t_L g1210 ( 
.A1(n_1088),
.A2(n_1037),
.B1(n_974),
.B2(n_979),
.C(n_1034),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1152),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1161),
.A2(n_986),
.B(n_1009),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1186),
.Y(n_1213)
);

CKINVDCx9p33_ASAP7_75t_R g1214 ( 
.A(n_1052),
.Y(n_1214)
);

AO31x2_ASAP7_75t_L g1215 ( 
.A1(n_1055),
.A2(n_1008),
.A3(n_1031),
.B(n_1021),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_SL g1216 ( 
.A1(n_1170),
.A2(n_1191),
.B(n_1155),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1182),
.A2(n_871),
.B(n_876),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1049),
.Y(n_1218)
);

AOI221x1_ASAP7_75t_L g1219 ( 
.A1(n_1153),
.A2(n_1020),
.B1(n_997),
.B2(n_1012),
.C(n_1001),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_1090),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1055),
.A2(n_982),
.A3(n_983),
.B(n_1036),
.Y(n_1221)
);

CKINVDCx16_ASAP7_75t_R g1222 ( 
.A(n_1114),
.Y(n_1222)
);

AO22x2_ASAP7_75t_L g1223 ( 
.A1(n_1079),
.A2(n_876),
.B1(n_909),
.B2(n_1056),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1062),
.B(n_1060),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1050),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1075),
.B(n_909),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1054),
.A2(n_1124),
.B(n_1046),
.Y(n_1227)
);

NAND2xp33_ASAP7_75t_L g1228 ( 
.A(n_1181),
.B(n_1184),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1070),
.Y(n_1229)
);

INVxp67_ASAP7_75t_SL g1230 ( 
.A(n_1082),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1054),
.A2(n_1068),
.B(n_1058),
.Y(n_1231)
);

OAI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1052),
.A2(n_1091),
.B1(n_1109),
.B2(n_1093),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1086),
.A2(n_1093),
.B1(n_1097),
.B2(n_1060),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1074),
.B(n_1169),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1144),
.B(n_1048),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1065),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1190),
.A2(n_1149),
.B(n_1180),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1122),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1072),
.Y(n_1239)
);

NOR4xp25_ASAP7_75t_L g1240 ( 
.A(n_1123),
.B(n_1115),
.C(n_1081),
.D(n_1163),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1049),
.B(n_1111),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1194),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1190),
.A2(n_1166),
.B(n_1157),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1076),
.A2(n_1174),
.B(n_1169),
.Y(n_1244)
);

INVx3_ASAP7_75t_SL g1245 ( 
.A(n_1044),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1063),
.A2(n_1078),
.B(n_1069),
.Y(n_1246)
);

OAI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1137),
.A2(n_1119),
.B1(n_1097),
.B2(n_1144),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1099),
.B(n_1057),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1195),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1122),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1045),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1077),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1196),
.A2(n_1189),
.A3(n_1174),
.B(n_1200),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1086),
.A2(n_1119),
.B1(n_1099),
.B2(n_1102),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1085),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1048),
.B(n_1071),
.Y(n_1256)
);

BUFx10_ASAP7_75t_L g1257 ( 
.A(n_1102),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1189),
.A2(n_1117),
.A3(n_1185),
.B(n_1051),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_SL g1259 ( 
.A1(n_1121),
.A2(n_1183),
.B(n_1179),
.C(n_1154),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1173),
.B(n_1176),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1139),
.A2(n_1073),
.B(n_1131),
.C(n_1129),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1206),
.A2(n_1204),
.B(n_1083),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1118),
.B(n_1120),
.Y(n_1263)
);

INVx3_ASAP7_75t_SL g1264 ( 
.A(n_1140),
.Y(n_1264)
);

OAI22x1_ASAP7_75t_L g1265 ( 
.A1(n_1103),
.A2(n_1150),
.B1(n_1139),
.B2(n_1066),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1151),
.A2(n_1126),
.B(n_1147),
.C(n_1080),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1095),
.A2(n_1094),
.B(n_1113),
.Y(n_1267)
);

AOI221xp5_ASAP7_75t_L g1268 ( 
.A1(n_1105),
.A2(n_1107),
.B1(n_1116),
.B2(n_1125),
.C(n_1101),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1085),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1167),
.A2(n_1092),
.B(n_1134),
.C(n_1172),
.Y(n_1270)
);

AOI221x1_ASAP7_75t_L g1271 ( 
.A1(n_1143),
.A2(n_1130),
.B1(n_1171),
.B2(n_1059),
.C(n_1104),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1091),
.B(n_1112),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_SL g1273 ( 
.A(n_1156),
.B(n_1121),
.C(n_1067),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1087),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1204),
.A2(n_1193),
.B(n_1187),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1173),
.B(n_1203),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1164),
.A2(n_1184),
.B1(n_1158),
.B2(n_1198),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1089),
.A2(n_1128),
.B1(n_1168),
.B2(n_1127),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1187),
.A2(n_1146),
.B(n_1154),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1199),
.A2(n_1202),
.B(n_1135),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1077),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1089),
.A2(n_1138),
.B1(n_1100),
.B2(n_1110),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1146),
.A2(n_1084),
.B(n_1133),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1061),
.A2(n_1053),
.B(n_1106),
.C(n_1140),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1145),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1175),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1205),
.A2(n_1160),
.B(n_1142),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1047),
.A2(n_1165),
.B1(n_1096),
.B2(n_1192),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1152),
.B(n_1047),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1100),
.A2(n_1136),
.A3(n_1128),
.B(n_1127),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1136),
.B(n_1201),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1132),
.A2(n_1092),
.B(n_1162),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1201),
.B(n_1096),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1165),
.A2(n_1098),
.B(n_1064),
.Y(n_1294)
);

AOI221xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1177),
.A2(n_1188),
.B1(n_1108),
.B2(n_1077),
.C(n_1197),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_SL g1296 ( 
.A1(n_1175),
.A2(n_1077),
.B(n_1108),
.C(n_1141),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1108),
.A2(n_1175),
.B(n_1197),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1141),
.A2(n_1148),
.B(n_1108),
.C(n_1197),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1197),
.A2(n_1148),
.A3(n_924),
.B(n_986),
.Y(n_1299)
);

AOI221xp5_ASAP7_75t_L g1300 ( 
.A1(n_1052),
.A2(n_691),
.B1(n_890),
.B2(n_998),
.C(n_800),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1178),
.A2(n_981),
.B(n_989),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1178),
.A2(n_981),
.B(n_989),
.Y(n_1303)
);

INVxp67_ASAP7_75t_L g1304 ( 
.A(n_1090),
.Y(n_1304)
);

O2A1O1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1153),
.A2(n_998),
.B(n_691),
.C(n_896),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1306)
);

BUFx12f_ASAP7_75t_L g1307 ( 
.A(n_1044),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1157),
.A2(n_1180),
.B(n_1166),
.Y(n_1308)
);

AO21x1_ASAP7_75t_L g1309 ( 
.A1(n_1062),
.A2(n_902),
.B(n_998),
.Y(n_1309)
);

A2O1A1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1093),
.A2(n_902),
.B(n_998),
.C(n_867),
.Y(n_1310)
);

OA21x2_ASAP7_75t_L g1311 ( 
.A1(n_1157),
.A2(n_1180),
.B(n_1166),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1052),
.B(n_908),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1313)
);

AOI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1178),
.A2(n_989),
.B(n_981),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1153),
.A2(n_998),
.B(n_691),
.C(n_896),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1178),
.A2(n_981),
.B(n_989),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1178),
.A2(n_981),
.B(n_989),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1052),
.B(n_534),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1178),
.A2(n_981),
.B(n_989),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1062),
.B(n_908),
.Y(n_1322)
);

OR2x6_ASAP7_75t_L g1323 ( 
.A(n_1049),
.B(n_1198),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1178),
.A2(n_981),
.B(n_989),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1325)
);

BUFx10_ASAP7_75t_L g1326 ( 
.A(n_1044),
.Y(n_1326)
);

BUFx8_ASAP7_75t_L g1327 ( 
.A(n_1122),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1052),
.B(n_534),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_1090),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1090),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1050),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1153),
.A2(n_902),
.B(n_1124),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1086),
.A2(n_902),
.B1(n_1097),
.B2(n_605),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1090),
.B(n_680),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1178),
.A2(n_981),
.B(n_989),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1062),
.B(n_908),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1178),
.A2(n_981),
.B(n_989),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1050),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1153),
.A2(n_902),
.B(n_1124),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1050),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1062),
.B(n_857),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1122),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1153),
.A2(n_902),
.B(n_1124),
.Y(n_1347)
);

NOR2xp67_ASAP7_75t_L g1348 ( 
.A(n_1057),
.B(n_742),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1122),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1062),
.B(n_857),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_SL g1352 ( 
.A1(n_1170),
.A2(n_1191),
.B(n_1155),
.Y(n_1352)
);

AO31x2_ASAP7_75t_L g1353 ( 
.A1(n_1055),
.A2(n_924),
.A3(n_986),
.B(n_1157),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1354)
);

BUFx2_ASAP7_75t_R g1355 ( 
.A(n_1044),
.Y(n_1355)
);

AO32x2_ASAP7_75t_L g1356 ( 
.A1(n_1171),
.A2(n_1051),
.A3(n_919),
.B1(n_860),
.B2(n_931),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1086),
.A2(n_902),
.B1(n_1097),
.B2(n_605),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1052),
.B(n_534),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1360)
);

INVx8_ASAP7_75t_L g1361 ( 
.A(n_1175),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1178),
.A2(n_981),
.B(n_989),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1054),
.A2(n_708),
.B(n_706),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1052),
.B(n_534),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1050),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1050),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1050),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1114),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1050),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1090),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1225),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1337),
.B(n_1224),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1336),
.A2(n_1357),
.B1(n_1359),
.B2(n_1329),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1236),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1239),
.Y(n_1375)
);

CKINVDCx11_ASAP7_75t_R g1376 ( 
.A(n_1307),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1254),
.A2(n_1300),
.B(n_1233),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1361),
.Y(n_1378)
);

INVx4_ASAP7_75t_SL g1379 ( 
.A(n_1323),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1327),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1254),
.A2(n_1233),
.B1(n_1357),
.B2(n_1336),
.Y(n_1381)
);

OAI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1224),
.A2(n_1232),
.B1(n_1235),
.B2(n_1247),
.Y(n_1382)
);

INVx8_ASAP7_75t_L g1383 ( 
.A(n_1361),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1333),
.Y(n_1384)
);

INVx6_ASAP7_75t_L g1385 ( 
.A(n_1361),
.Y(n_1385)
);

INVx3_ASAP7_75t_SL g1386 ( 
.A(n_1368),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1370),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1238),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1320),
.A2(n_1364),
.B1(n_1309),
.B2(n_1342),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1341),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1343),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1209),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1335),
.A2(n_1342),
.B1(n_1347),
.B2(n_1344),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1365),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1312),
.B(n_1230),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1335),
.A2(n_1347),
.B1(n_1351),
.B2(n_1344),
.Y(n_1396)
);

INVx4_ASAP7_75t_L g1397 ( 
.A(n_1285),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1351),
.A2(n_1223),
.B1(n_1257),
.B2(n_1272),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1322),
.B(n_1339),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1245),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1223),
.A2(n_1257),
.B1(n_1248),
.B2(n_1352),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1216),
.A2(n_1265),
.B1(n_1268),
.B2(n_1226),
.Y(n_1402)
);

BUFx4_ASAP7_75t_SL g1403 ( 
.A(n_1250),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1366),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1222),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1228),
.A2(n_1310),
.B1(n_1214),
.B2(n_1244),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1327),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1213),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1229),
.B(n_1331),
.Y(n_1409)
);

BUFx10_ASAP7_75t_L g1410 ( 
.A(n_1241),
.Y(n_1410)
);

INVx6_ASAP7_75t_L g1411 ( 
.A(n_1218),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1218),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1331),
.B(n_1332),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1264),
.Y(n_1414)
);

INVx6_ASAP7_75t_L g1415 ( 
.A(n_1218),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1244),
.A2(n_1260),
.B1(n_1277),
.B2(n_1256),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1249),
.A2(n_1332),
.B1(n_1367),
.B2(n_1369),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1234),
.A2(n_1276),
.B1(n_1260),
.B2(n_1242),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1234),
.A2(n_1276),
.B1(n_1304),
.B2(n_1220),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1263),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1251),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1345),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1286),
.Y(n_1423)
);

INVx3_ASAP7_75t_SL g1424 ( 
.A(n_1326),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1350),
.Y(n_1425)
);

BUFx4_ASAP7_75t_R g1426 ( 
.A(n_1326),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1252),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1273),
.A2(n_1348),
.B1(n_1360),
.B2(n_1358),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1277),
.A2(n_1305),
.B1(n_1315),
.B2(n_1237),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1255),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1323),
.A2(n_1240),
.B1(n_1283),
.B2(n_1211),
.Y(n_1431)
);

BUFx12f_ASAP7_75t_L g1432 ( 
.A(n_1323),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1301),
.A2(n_1363),
.B1(n_1306),
.B2(n_1313),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1269),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1252),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1281),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_1355),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1261),
.A2(n_1266),
.B1(n_1270),
.B2(n_1243),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1274),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1316),
.A2(n_1334),
.B1(n_1325),
.B2(n_1317),
.Y(n_1440)
);

OAI21xp33_ASAP7_75t_L g1441 ( 
.A1(n_1240),
.A2(n_1227),
.B(n_1328),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1330),
.A2(n_1354),
.B1(n_1349),
.B2(n_1346),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1281),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_1289),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1281),
.Y(n_1445)
);

INVx6_ASAP7_75t_L g1446 ( 
.A(n_1296),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1291),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1291),
.A2(n_1280),
.B1(n_1208),
.B2(n_1288),
.Y(n_1448)
);

INVx6_ASAP7_75t_L g1449 ( 
.A(n_1295),
.Y(n_1449)
);

CKINVDCx11_ASAP7_75t_R g1450 ( 
.A(n_1295),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1280),
.A2(n_1278),
.B1(n_1282),
.B2(n_1293),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1253),
.B(n_1293),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1284),
.A2(n_1271),
.B(n_1287),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1262),
.A2(n_1356),
.B1(n_1279),
.B2(n_1275),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1294),
.Y(n_1455)
);

INVx6_ASAP7_75t_L g1456 ( 
.A(n_1298),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1356),
.A2(n_1311),
.B1(n_1308),
.B2(n_1292),
.Y(n_1457)
);

OAI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1356),
.A2(n_1219),
.B1(n_1210),
.B2(n_1231),
.Y(n_1458)
);

BUFx4f_ASAP7_75t_SL g1459 ( 
.A(n_1259),
.Y(n_1459)
);

INVx6_ASAP7_75t_L g1460 ( 
.A(n_1297),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1308),
.A2(n_1311),
.B1(n_1246),
.B2(n_1253),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1253),
.A2(n_1314),
.B1(n_1258),
.B2(n_1353),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1299),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1258),
.A2(n_1353),
.B1(n_1215),
.B2(n_1217),
.Y(n_1464)
);

INVx8_ASAP7_75t_L g1465 ( 
.A(n_1299),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1207),
.A2(n_1212),
.B1(n_1353),
.B2(n_1267),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1290),
.B(n_1258),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1215),
.A2(n_1221),
.B1(n_1302),
.B2(n_1303),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1318),
.A2(n_1362),
.B1(n_1319),
.B2(n_1321),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1324),
.B(n_1338),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1221),
.B(n_1340),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1221),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1307),
.Y(n_1473)
);

BUFx12f_ASAP7_75t_L g1474 ( 
.A(n_1327),
.Y(n_1474)
);

CKINVDCx11_ASAP7_75t_R g1475 ( 
.A(n_1307),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1224),
.B(n_1235),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1307),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_1222),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1225),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1218),
.Y(n_1480)
);

INVx3_ASAP7_75t_SL g1481 ( 
.A(n_1368),
.Y(n_1481)
);

INVx6_ASAP7_75t_L g1482 ( 
.A(n_1361),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1209),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1336),
.A2(n_1357),
.B1(n_1300),
.B2(n_745),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1254),
.A2(n_1320),
.B1(n_1359),
.B2(n_1329),
.Y(n_1485)
);

AO22x1_ASAP7_75t_L g1486 ( 
.A1(n_1320),
.A2(n_691),
.B1(n_1359),
.B2(n_1329),
.Y(n_1486)
);

BUFx8_ASAP7_75t_SL g1487 ( 
.A(n_1307),
.Y(n_1487)
);

OAI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1254),
.A2(n_1233),
.B1(n_1357),
.B2(n_1336),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_1222),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1307),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1225),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1225),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1209),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1337),
.Y(n_1494)
);

INVx6_ASAP7_75t_L g1495 ( 
.A(n_1361),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1225),
.Y(n_1496)
);

OAI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1254),
.A2(n_1233),
.B1(n_1357),
.B2(n_1336),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1336),
.A2(n_1357),
.B1(n_1300),
.B2(n_745),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1254),
.A2(n_1320),
.B1(n_1359),
.B2(n_1329),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1238),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1336),
.A2(n_693),
.B1(n_1357),
.B2(n_691),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1361),
.Y(n_1502)
);

BUFx10_ASAP7_75t_L g1503 ( 
.A(n_1368),
.Y(n_1503)
);

INVx6_ASAP7_75t_L g1504 ( 
.A(n_1361),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_1222),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1336),
.A2(n_1357),
.B1(n_1300),
.B2(n_745),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1225),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1336),
.A2(n_693),
.B1(n_1357),
.B2(n_691),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1336),
.A2(n_1357),
.B1(n_1300),
.B2(n_745),
.Y(n_1509)
);

BUFx8_ASAP7_75t_L g1510 ( 
.A(n_1307),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1238),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1225),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1225),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1336),
.A2(n_1357),
.B1(n_1300),
.B2(n_745),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1300),
.A2(n_691),
.B1(n_1329),
.B2(n_1320),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1225),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1336),
.A2(n_1357),
.B1(n_1300),
.B2(n_745),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1430),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1439),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1395),
.B(n_1476),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1515),
.A2(n_1377),
.B(n_1485),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1461),
.A2(n_1471),
.B(n_1442),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1372),
.B(n_1396),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1420),
.Y(n_1524)
);

CKINVDCx16_ASAP7_75t_R g1525 ( 
.A(n_1405),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1387),
.Y(n_1526)
);

INVx4_ASAP7_75t_SL g1527 ( 
.A(n_1449),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1452),
.Y(n_1528)
);

INVx4_ASAP7_75t_L g1529 ( 
.A(n_1449),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1393),
.B(n_1371),
.Y(n_1530)
);

OAI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1499),
.A2(n_1389),
.B(n_1438),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1472),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1449),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1470),
.A2(n_1466),
.B(n_1464),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1466),
.A2(n_1469),
.B(n_1440),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1409),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1373),
.A2(n_1389),
.B1(n_1514),
.B2(n_1484),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1413),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1469),
.A2(n_1440),
.B(n_1433),
.Y(n_1539)
);

AO31x2_ASAP7_75t_L g1540 ( 
.A1(n_1462),
.A2(n_1463),
.A3(n_1467),
.B(n_1434),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1421),
.Y(n_1541)
);

OA21x2_ASAP7_75t_L g1542 ( 
.A1(n_1457),
.A2(n_1441),
.B(n_1454),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1393),
.B(n_1374),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1375),
.Y(n_1544)
);

CKINVDCx20_ASAP7_75t_R g1545 ( 
.A(n_1437),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1384),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1455),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1390),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1391),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1446),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1501),
.A2(n_1508),
.B1(n_1484),
.B2(n_1506),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1394),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1381),
.B(n_1488),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1465),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1404),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1479),
.B(n_1491),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1381),
.B(n_1488),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1400),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1433),
.A2(n_1457),
.B(n_1454),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1447),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1486),
.B(n_1397),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1460),
.Y(n_1562)
);

NOR2xp67_ASAP7_75t_L g1563 ( 
.A(n_1453),
.B(n_1427),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1492),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1496),
.B(n_1507),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1396),
.B(n_1494),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1498),
.A2(n_1517),
.B1(n_1506),
.B2(n_1509),
.Y(n_1567)
);

NOR2x1_ASAP7_75t_R g1568 ( 
.A(n_1474),
.B(n_1376),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1512),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1513),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1516),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1398),
.B(n_1418),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1446),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1459),
.Y(n_1574)
);

OAI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1448),
.A2(n_1428),
.B(n_1451),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1459),
.Y(n_1576)
);

AO21x2_ASAP7_75t_L g1577 ( 
.A1(n_1458),
.A2(n_1468),
.B(n_1497),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1379),
.B(n_1398),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1392),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1399),
.Y(n_1580)
);

INVxp33_ASAP7_75t_SL g1581 ( 
.A(n_1403),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1408),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1448),
.A2(n_1451),
.B(n_1517),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1446),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1410),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1483),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1493),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1487),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1468),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1419),
.B(n_1418),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1458),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1397),
.B(n_1386),
.Y(n_1592)
);

OAI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1428),
.A2(n_1402),
.B(n_1401),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1416),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1402),
.A2(n_1401),
.B(n_1436),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1456),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1497),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1498),
.A2(n_1514),
.B(n_1509),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1410),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1419),
.B(n_1382),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1417),
.B(n_1406),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1417),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1456),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1429),
.A2(n_1382),
.B(n_1431),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1456),
.Y(n_1605)
);

AO21x2_ASAP7_75t_L g1606 ( 
.A1(n_1450),
.A2(n_1445),
.B(n_1444),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1443),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1412),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1412),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1480),
.Y(n_1610)
);

OA21x2_ASAP7_75t_L g1611 ( 
.A1(n_1388),
.A2(n_1511),
.B(n_1425),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1502),
.B(n_1422),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1500),
.B(n_1481),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1502),
.B(n_1423),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1478),
.A2(n_1489),
.B1(n_1505),
.B2(n_1482),
.Y(n_1615)
);

AOI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1423),
.A2(n_1490),
.B1(n_1477),
.B2(n_1473),
.C(n_1424),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1411),
.B(n_1415),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1432),
.A2(n_1415),
.B1(n_1475),
.B2(n_1435),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1386),
.B(n_1481),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1378),
.A2(n_1504),
.B(n_1495),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1385),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1385),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1403),
.Y(n_1623)
);

OR2x6_ASAP7_75t_L g1624 ( 
.A(n_1383),
.B(n_1482),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1536),
.B(n_1503),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1521),
.B(n_1426),
.Y(n_1626)
);

A2O1A1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1604),
.A2(n_1598),
.B(n_1521),
.C(n_1531),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1531),
.A2(n_1383),
.B(n_1414),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1562),
.Y(n_1629)
);

O2A1O1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1537),
.A2(n_1503),
.B(n_1510),
.C(n_1383),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1548),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1560),
.B(n_1524),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1569),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_SL g1634 ( 
.A1(n_1594),
.A2(n_1380),
.B(n_1407),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1567),
.A2(n_1495),
.B(n_1504),
.C(n_1510),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1600),
.A2(n_1591),
.B1(n_1590),
.B2(n_1572),
.C(n_1601),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1570),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1570),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1556),
.B(n_1565),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1556),
.B(n_1565),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1611),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1553),
.A2(n_1557),
.B(n_1593),
.Y(n_1642)
);

AO32x2_ASAP7_75t_L g1643 ( 
.A1(n_1529),
.A2(n_1573),
.A3(n_1550),
.B1(n_1585),
.B2(n_1599),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1528),
.B(n_1577),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1557),
.A2(n_1567),
.B1(n_1551),
.B2(n_1597),
.Y(n_1645)
);

AND2x2_ASAP7_75t_SL g1646 ( 
.A(n_1572),
.B(n_1583),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1538),
.B(n_1570),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1601),
.A2(n_1603),
.B1(n_1533),
.B2(n_1597),
.Y(n_1648)
);

OA21x2_ASAP7_75t_L g1649 ( 
.A1(n_1522),
.A2(n_1539),
.B(n_1559),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1544),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1574),
.B(n_1576),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1580),
.B(n_1566),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1530),
.B(n_1543),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1574),
.A2(n_1576),
.B1(n_1533),
.B2(n_1529),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1530),
.B(n_1543),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1520),
.B(n_1526),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1589),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1611),
.B(n_1608),
.Y(n_1658)
);

NAND2xp33_ASAP7_75t_R g1659 ( 
.A(n_1584),
.B(n_1611),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1523),
.B(n_1546),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1611),
.B(n_1533),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1546),
.B(n_1549),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1617),
.B(n_1609),
.Y(n_1663)
);

A2O1A1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1593),
.A2(n_1575),
.B(n_1595),
.C(n_1561),
.Y(n_1664)
);

OA21x2_ASAP7_75t_L g1665 ( 
.A1(n_1535),
.A2(n_1534),
.B(n_1595),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1578),
.B(n_1527),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1602),
.A2(n_1577),
.B1(n_1571),
.B2(n_1564),
.C(n_1555),
.Y(n_1667)
);

INVx4_ASAP7_75t_L g1668 ( 
.A(n_1527),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1552),
.B(n_1555),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1603),
.A2(n_1583),
.B1(n_1596),
.B2(n_1605),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_SL g1671 ( 
.A1(n_1615),
.A2(n_1602),
.B1(n_1616),
.B2(n_1621),
.C(n_1610),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1578),
.B(n_1527),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1583),
.A2(n_1605),
.B1(n_1596),
.B2(n_1577),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1518),
.B(n_1519),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1519),
.B(n_1541),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1563),
.A2(n_1605),
.B(n_1535),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1583),
.A2(n_1578),
.B1(n_1542),
.B2(n_1606),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1579),
.B(n_1607),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1525),
.A2(n_1623),
.B1(n_1624),
.B2(n_1581),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1584),
.A2(n_1620),
.B(n_1542),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_L g1681 ( 
.A(n_1542),
.B(n_1607),
.C(n_1584),
.Y(n_1681)
);

AOI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1532),
.A2(n_1618),
.B1(n_1587),
.B2(n_1582),
.C(n_1586),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1525),
.A2(n_1624),
.B1(n_1613),
.B2(n_1622),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_SL g1684 ( 
.A1(n_1545),
.A2(n_1588),
.B1(n_1558),
.B2(n_1619),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1637),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1638),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1639),
.B(n_1542),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1650),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1643),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1641),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1640),
.B(n_1534),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1658),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1644),
.B(n_1547),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1649),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1660),
.B(n_1540),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1641),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1649),
.B(n_1547),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1653),
.B(n_1655),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1657),
.B(n_1656),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1657),
.B(n_1540),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1667),
.B(n_1540),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1675),
.Y(n_1702)
);

AND2x4_ASAP7_75t_SL g1703 ( 
.A(n_1668),
.B(n_1666),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1661),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1631),
.B(n_1540),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1633),
.B(n_1540),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1662),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1627),
.B(n_1540),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1669),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1629),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1659),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1665),
.B(n_1532),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1674),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1699),
.Y(n_1714)
);

INVx4_ASAP7_75t_L g1715 ( 
.A(n_1710),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1685),
.Y(n_1716)
);

OAI33xp33_ASAP7_75t_L g1717 ( 
.A1(n_1708),
.A2(n_1645),
.A3(n_1652),
.B1(n_1679),
.B2(n_1647),
.B3(n_1683),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1708),
.A2(n_1626),
.B(n_1627),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1685),
.Y(n_1719)
);

AOI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1708),
.A2(n_1636),
.B1(n_1671),
.B2(n_1664),
.C(n_1642),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1712),
.Y(n_1721)
);

AOI221xp5_ASAP7_75t_L g1722 ( 
.A1(n_1701),
.A2(n_1711),
.B1(n_1689),
.B2(n_1695),
.C(n_1700),
.Y(n_1722)
);

OAI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1711),
.A2(n_1664),
.B1(n_1659),
.B2(n_1626),
.C(n_1677),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1698),
.B(n_1632),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1698),
.B(n_1663),
.Y(n_1725)
);

OAI21x1_ASAP7_75t_L g1726 ( 
.A1(n_1694),
.A2(n_1680),
.B(n_1676),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1707),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1698),
.B(n_1673),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1701),
.A2(n_1646),
.B1(n_1677),
.B2(n_1606),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1699),
.B(n_1646),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1712),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1707),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1689),
.B(n_1625),
.Y(n_1733)
);

OAI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1700),
.A2(n_1648),
.B1(n_1670),
.B2(n_1634),
.C(n_1682),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1694),
.Y(n_1735)
);

NOR3xp33_ASAP7_75t_L g1736 ( 
.A(n_1705),
.B(n_1630),
.C(n_1654),
.Y(n_1736)
);

BUFx5_ASAP7_75t_L g1737 ( 
.A(n_1712),
.Y(n_1737)
);

NOR2xp67_ASAP7_75t_L g1738 ( 
.A(n_1700),
.B(n_1681),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1687),
.B(n_1678),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1709),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1687),
.A2(n_1606),
.B1(n_1672),
.B2(n_1554),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1703),
.B(n_1672),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1685),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1691),
.B(n_1651),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1686),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1691),
.B(n_1643),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1704),
.B(n_1643),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1747),
.B(n_1692),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1715),
.B(n_1721),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1747),
.B(n_1692),
.Y(n_1750)
);

OAI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1718),
.A2(n_1634),
.B1(n_1635),
.B2(n_1695),
.C(n_1705),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1716),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1746),
.B(n_1704),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1746),
.B(n_1704),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1714),
.B(n_1706),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1737),
.B(n_1704),
.Y(n_1756)
);

INVxp67_ASAP7_75t_SL g1757 ( 
.A(n_1738),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1737),
.B(n_1744),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1742),
.B(n_1703),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1737),
.B(n_1687),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1716),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1737),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1737),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1737),
.B(n_1687),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1719),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1714),
.B(n_1706),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1719),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1737),
.B(n_1693),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1718),
.B(n_1713),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1737),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1728),
.B(n_1713),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1721),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1721),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1744),
.B(n_1693),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1727),
.B(n_1688),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1743),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1728),
.B(n_1702),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1743),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_L g1779 ( 
.A(n_1720),
.B(n_1694),
.C(n_1697),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1745),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1739),
.B(n_1702),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1715),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1731),
.B(n_1697),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1739),
.B(n_1702),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1731),
.B(n_1697),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1769),
.B(n_1732),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1753),
.B(n_1733),
.Y(n_1787)
);

NAND2x1_ASAP7_75t_L g1788 ( 
.A(n_1756),
.B(n_1782),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1757),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1752),
.Y(n_1790)
);

AOI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1779),
.A2(n_1723),
.B1(n_1717),
.B2(n_1729),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1752),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1769),
.B(n_1722),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1752),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1772),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_R g1796 ( 
.A(n_1756),
.B(n_1592),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_1759),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1771),
.B(n_1740),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1753),
.B(n_1754),
.Y(n_1799)
);

INVxp67_ASAP7_75t_SL g1800 ( 
.A(n_1757),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1761),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1761),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1771),
.B(n_1725),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1771),
.B(n_1725),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1761),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1753),
.B(n_1733),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1772),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1765),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1765),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1779),
.B(n_1738),
.Y(n_1810)
);

NOR2xp67_ASAP7_75t_L g1811 ( 
.A(n_1759),
.B(n_1715),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1775),
.B(n_1730),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1751),
.B(n_1568),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1772),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1777),
.Y(n_1815)
);

OAI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1751),
.A2(n_1734),
.B1(n_1741),
.B2(n_1736),
.C(n_1696),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1765),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1767),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1767),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1777),
.B(n_1568),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1754),
.B(n_1742),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1775),
.B(n_1724),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1767),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1754),
.B(n_1742),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1776),
.Y(n_1825)
);

OR2x2_ASAP7_75t_SL g1826 ( 
.A(n_1762),
.B(n_1613),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1776),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1774),
.B(n_1756),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1815),
.B(n_1776),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1800),
.B(n_1774),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1803),
.B(n_1804),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1789),
.B(n_1774),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1799),
.B(n_1758),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1794),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1789),
.B(n_1748),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1794),
.Y(n_1836)
);

NAND4xp25_ASAP7_75t_L g1837 ( 
.A(n_1810),
.B(n_1684),
.C(n_1782),
.D(n_1628),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1793),
.B(n_1778),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1791),
.B(n_1778),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1795),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1801),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1801),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1786),
.B(n_1748),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1802),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1795),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1803),
.B(n_1781),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1802),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1786),
.B(n_1748),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1799),
.B(n_1821),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1821),
.B(n_1824),
.Y(n_1850)
);

BUFx2_ASAP7_75t_SL g1851 ( 
.A(n_1811),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1805),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1804),
.B(n_1781),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1805),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1798),
.B(n_1750),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1824),
.B(n_1758),
.Y(n_1856)
);

INVx2_ASAP7_75t_SL g1857 ( 
.A(n_1788),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1787),
.B(n_1758),
.Y(n_1858)
);

BUFx2_ASAP7_75t_L g1859 ( 
.A(n_1797),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1787),
.B(n_1750),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1825),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1806),
.B(n_1750),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1806),
.B(n_1768),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1820),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1864),
.B(n_1813),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1850),
.B(n_1849),
.Y(n_1866)
);

AOI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1839),
.A2(n_1816),
.B1(n_1812),
.B2(n_1814),
.C(n_1807),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1839),
.A2(n_1797),
.B1(n_1826),
.B2(n_1798),
.Y(n_1868)
);

NAND2xp33_ASAP7_75t_SL g1869 ( 
.A(n_1859),
.B(n_1788),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1859),
.Y(n_1870)
);

O2A1O1Ixp5_ASAP7_75t_SL g1871 ( 
.A1(n_1834),
.A2(n_1825),
.B(n_1827),
.C(n_1790),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_SL g1872 ( 
.A1(n_1837),
.A2(n_1828),
.B(n_1782),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1850),
.B(n_1828),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1838),
.A2(n_1826),
.B1(n_1822),
.B2(n_1777),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1838),
.B(n_1792),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1831),
.B(n_1781),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1849),
.Y(n_1877)
);

AOI22xp5_ASAP7_75t_SL g1878 ( 
.A1(n_1864),
.A2(n_1796),
.B1(n_1764),
.B2(n_1760),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1834),
.Y(n_1879)
);

AOI31xp33_ASAP7_75t_L g1880 ( 
.A1(n_1835),
.A2(n_1796),
.A3(n_1760),
.B(n_1764),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1843),
.A2(n_1848),
.B1(n_1830),
.B2(n_1832),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1837),
.A2(n_1696),
.B1(n_1690),
.B2(n_1807),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_SL g1883 ( 
.A1(n_1851),
.A2(n_1770),
.B1(n_1762),
.B2(n_1763),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1856),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1856),
.Y(n_1885)
);

OAI21xp33_ASAP7_75t_L g1886 ( 
.A1(n_1855),
.A2(n_1809),
.B(n_1808),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1836),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1840),
.A2(n_1696),
.B1(n_1690),
.B2(n_1814),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1840),
.A2(n_1845),
.B1(n_1831),
.B2(n_1862),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1829),
.A2(n_1766),
.B(n_1755),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1876),
.B(n_1846),
.Y(n_1891)
);

INVxp67_ASAP7_75t_L g1892 ( 
.A(n_1870),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1879),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1877),
.B(n_1860),
.Y(n_1894)
);

A2O1A1Ixp33_ASAP7_75t_SL g1895 ( 
.A1(n_1889),
.A2(n_1847),
.B(n_1841),
.C(n_1861),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1866),
.B(n_1860),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1887),
.Y(n_1897)
);

NOR3xp33_ASAP7_75t_L g1898 ( 
.A(n_1868),
.B(n_1829),
.C(n_1836),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1873),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1875),
.Y(n_1900)
);

AOI221x1_ASAP7_75t_L g1901 ( 
.A1(n_1865),
.A2(n_1851),
.B1(n_1854),
.B2(n_1861),
.C(n_1841),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1884),
.B(n_1862),
.Y(n_1902)
);

INVxp67_ASAP7_75t_SL g1903 ( 
.A(n_1868),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1867),
.A2(n_1840),
.B1(n_1845),
.B2(n_1846),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1885),
.B(n_1833),
.Y(n_1905)
);

OAI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1882),
.A2(n_1853),
.B1(n_1845),
.B2(n_1766),
.Y(n_1906)
);

AOI222xp33_ASAP7_75t_L g1907 ( 
.A1(n_1874),
.A2(n_1842),
.B1(n_1844),
.B2(n_1854),
.C1(n_1847),
.C2(n_1852),
.Y(n_1907)
);

OAI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1880),
.A2(n_1853),
.B1(n_1755),
.B2(n_1766),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1881),
.B(n_1857),
.Y(n_1909)
);

NAND2xp33_ASAP7_75t_SL g1910 ( 
.A(n_1881),
.B(n_1857),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1891),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1892),
.Y(n_1912)
);

OAI22xp33_ASAP7_75t_L g1913 ( 
.A1(n_1903),
.A2(n_1872),
.B1(n_1874),
.B2(n_1875),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1905),
.B(n_1886),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1899),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1892),
.Y(n_1916)
);

O2A1O1Ixp33_ASAP7_75t_L g1917 ( 
.A1(n_1895),
.A2(n_1890),
.B(n_1871),
.C(n_1852),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1894),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1909),
.B(n_1878),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1902),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1896),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1900),
.Y(n_1922)
);

NAND4xp25_ASAP7_75t_L g1923 ( 
.A(n_1917),
.B(n_1901),
.C(n_1910),
.D(n_1898),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1911),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1921),
.B(n_1898),
.Y(n_1925)
);

OAI21xp33_ASAP7_75t_L g1926 ( 
.A1(n_1919),
.A2(n_1914),
.B(n_1918),
.Y(n_1926)
);

OAI21xp33_ASAP7_75t_SL g1927 ( 
.A1(n_1919),
.A2(n_1907),
.B(n_1897),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1912),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1913),
.B(n_1869),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1915),
.B(n_1833),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1913),
.A2(n_1904),
.B(n_1908),
.Y(n_1931)
);

NAND3xp33_ASAP7_75t_L g1932 ( 
.A(n_1915),
.B(n_1893),
.C(n_1906),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1916),
.Y(n_1933)
);

AOI211x1_ASAP7_75t_L g1934 ( 
.A1(n_1920),
.A2(n_1844),
.B(n_1842),
.C(n_1858),
.Y(n_1934)
);

OAI221xp5_ASAP7_75t_SL g1935 ( 
.A1(n_1927),
.A2(n_1922),
.B1(n_1888),
.B2(n_1858),
.C(n_1883),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1923),
.B(n_1922),
.Y(n_1936)
);

O2A1O1Ixp33_ASAP7_75t_L g1937 ( 
.A1(n_1931),
.A2(n_1823),
.B(n_1819),
.C(n_1818),
.Y(n_1937)
);

O2A1O1Ixp33_ASAP7_75t_L g1938 ( 
.A1(n_1929),
.A2(n_1817),
.B(n_1863),
.C(n_1755),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1930),
.Y(n_1939)
);

NAND4xp25_ASAP7_75t_L g1940 ( 
.A(n_1926),
.B(n_1863),
.C(n_1782),
.D(n_1760),
.Y(n_1940)
);

OAI221xp5_ASAP7_75t_L g1941 ( 
.A1(n_1935),
.A2(n_1932),
.B1(n_1925),
.B2(n_1928),
.C(n_1933),
.Y(n_1941)
);

AOI211xp5_ASAP7_75t_SL g1942 ( 
.A1(n_1936),
.A2(n_1928),
.B(n_1924),
.C(n_1934),
.Y(n_1942)
);

AOI221xp5_ASAP7_75t_L g1943 ( 
.A1(n_1937),
.A2(n_1694),
.B1(n_1772),
.B2(n_1773),
.C(n_1785),
.Y(n_1943)
);

AOI221xp5_ASAP7_75t_L g1944 ( 
.A1(n_1938),
.A2(n_1694),
.B1(n_1773),
.B2(n_1785),
.C(n_1783),
.Y(n_1944)
);

OAI211xp5_ASAP7_75t_L g1945 ( 
.A1(n_1939),
.A2(n_1940),
.B(n_1782),
.C(n_1763),
.Y(n_1945)
);

NOR3xp33_ASAP7_75t_L g1946 ( 
.A(n_1936),
.B(n_1635),
.C(n_1726),
.Y(n_1946)
);

XNOR2xp5_ASAP7_75t_L g1947 ( 
.A(n_1941),
.B(n_1612),
.Y(n_1947)
);

NAND4xp75_ASAP7_75t_L g1948 ( 
.A(n_1944),
.B(n_1764),
.C(n_1763),
.D(n_1770),
.Y(n_1948)
);

XNOR2x1_ASAP7_75t_L g1949 ( 
.A(n_1942),
.B(n_1726),
.Y(n_1949)
);

XOR2xp5_ASAP7_75t_L g1950 ( 
.A(n_1946),
.B(n_1784),
.Y(n_1950)
);

OAI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1943),
.A2(n_1770),
.B1(n_1762),
.B2(n_1763),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1947),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1949),
.B(n_1945),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1950),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1953),
.A2(n_1951),
.B1(n_1782),
.B2(n_1948),
.Y(n_1955)
);

INVxp67_ASAP7_75t_SL g1956 ( 
.A(n_1955),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_SL g1957 ( 
.A1(n_1956),
.A2(n_1954),
.B1(n_1952),
.B2(n_1953),
.Y(n_1957)
);

AOI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1956),
.A2(n_1952),
.B1(n_1773),
.B2(n_1770),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1957),
.Y(n_1959)
);

NOR2x1_ASAP7_75t_L g1960 ( 
.A(n_1958),
.B(n_1749),
.Y(n_1960)
);

AO21x2_ASAP7_75t_L g1961 ( 
.A1(n_1959),
.A2(n_1780),
.B(n_1778),
.Y(n_1961)
);

AOI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1960),
.A2(n_1773),
.B(n_1785),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1961),
.Y(n_1963)
);

OAI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1963),
.A2(n_1962),
.B1(n_1762),
.B2(n_1784),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1964),
.Y(n_1965)
);

OAI221xp5_ASAP7_75t_R g1966 ( 
.A1(n_1965),
.A2(n_1749),
.B1(n_1735),
.B2(n_1780),
.C(n_1783),
.Y(n_1966)
);

AOI211xp5_ASAP7_75t_L g1967 ( 
.A1(n_1966),
.A2(n_1612),
.B(n_1614),
.C(n_1749),
.Y(n_1967)
);


endmodule