module fake_jpeg_29339_n_102 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_20),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_51),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_38),
.B1(n_43),
.B2(n_4),
.Y(n_61)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_53),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_13),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_40),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_3),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_41),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_7),
.B(n_8),
.Y(n_80)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_42),
.B1(n_34),
.B2(n_14),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_74),
.B1(n_75),
.B2(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_68),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_1),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_73),
.B(n_6),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_72),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_5),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_61),
.B1(n_73),
.B2(n_74),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_79),
.Y(n_91)
);

AND2x6_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_18),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

AOI22x1_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_21),
.B1(n_28),
.B2(n_10),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_22),
.B(n_27),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_87),
.A2(n_15),
.B(n_26),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_93),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_8),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_85),
.C(n_82),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_92),
.C(n_91),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_79),
.A3(n_89),
.B1(n_81),
.B2(n_84),
.C1(n_86),
.C2(n_90),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_94),
.B(n_11),
.Y(n_101)
);

A2O1A1O1Ixp25_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_12),
.B(n_24),
.C(n_32),
.D(n_9),
.Y(n_102)
);


endmodule