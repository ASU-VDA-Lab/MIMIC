module real_aes_7936_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_704, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_704;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_404;
wire n_147;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
wire n_237;
A2O1A1Ixp33_ASAP7_75t_SL g157 ( .A1(n_0), .A2(n_158), .B(n_159), .C(n_163), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_1), .B(n_152), .Y(n_165) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_3), .B(n_137), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_4), .A2(n_126), .B(n_143), .C(n_434), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_5), .A2(n_146), .B(n_455), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_6), .A2(n_146), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_7), .B(n_152), .Y(n_461) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_8), .A2(n_118), .B(n_205), .Y(n_204) );
AND2x6_ASAP7_75t_L g143 ( .A(n_9), .B(n_144), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_10), .A2(n_126), .B(n_143), .C(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g426 ( .A(n_11), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_12), .B(n_40), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_13), .B(n_162), .Y(n_436) );
INVx1_ASAP7_75t_L g123 ( .A(n_14), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_15), .B(n_137), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g444 ( .A1(n_16), .A2(n_138), .B(n_445), .C(n_447), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_17), .B(n_152), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g689 ( .A1(n_18), .A2(n_65), .B1(n_690), .B2(n_691), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_18), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_19), .B(n_195), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_20), .A2(n_126), .B(n_189), .C(n_194), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g415 ( .A1(n_21), .A2(n_161), .B(n_213), .C(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_22), .B(n_162), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_23), .B(n_162), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_24), .Y(n_464) );
INVx1_ASAP7_75t_L g476 ( .A(n_25), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_26), .A2(n_126), .B(n_194), .C(n_208), .Y(n_207) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_27), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_28), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_29), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g493 ( .A(n_30), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_31), .A2(n_146), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g128 ( .A(n_32), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_33), .A2(n_141), .B(n_173), .C(n_174), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_34), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_35), .A2(n_161), .B(n_458), .C(n_460), .Y(n_457) );
INVxp67_ASAP7_75t_L g494 ( .A(n_36), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_37), .B(n_210), .Y(n_209) );
CKINVDCx14_ASAP7_75t_R g456 ( .A(n_38), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_39), .A2(n_126), .B(n_194), .C(n_475), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g423 ( .A1(n_41), .A2(n_163), .B(n_424), .C(n_425), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_42), .B(n_187), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_43), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_44), .B(n_137), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_45), .B(n_146), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_46), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_47), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_48), .A2(n_141), .B(n_173), .C(n_234), .Y(n_233) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_49), .A2(n_103), .B1(n_666), .B2(n_667), .C1(n_670), .C2(n_674), .Y(n_102) );
INVx1_ASAP7_75t_L g160 ( .A(n_50), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_51), .A2(n_81), .B1(n_668), .B2(n_669), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_51), .Y(n_669) );
INVx1_ASAP7_75t_L g235 ( .A(n_52), .Y(n_235) );
INVx1_ASAP7_75t_L g414 ( .A(n_53), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_54), .B(n_146), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_55), .Y(n_198) );
CKINVDCx14_ASAP7_75t_R g422 ( .A(n_56), .Y(n_422) );
INVx1_ASAP7_75t_L g144 ( .A(n_57), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_58), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_59), .B(n_152), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_60), .A2(n_133), .B(n_193), .C(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g122 ( .A(n_61), .Y(n_122) );
INVx1_ASAP7_75t_SL g459 ( .A(n_62), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_63), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_64), .B(n_137), .Y(n_178) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_65), .A2(n_101), .B1(n_678), .B2(n_687), .C1(n_696), .C2(n_700), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_65), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_66), .B(n_152), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_67), .B(n_138), .Y(n_224) );
INVx1_ASAP7_75t_L g467 ( .A(n_68), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g155 ( .A(n_69), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_70), .B(n_177), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g125 ( .A1(n_71), .A2(n_126), .B(n_131), .C(n_141), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g249 ( .A(n_72), .Y(n_249) );
INVx1_ASAP7_75t_L g682 ( .A(n_73), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_74), .A2(n_146), .B(n_421), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_75), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_76), .A2(n_146), .B(n_442), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_77), .A2(n_187), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g443 ( .A(n_78), .Y(n_443) );
CKINVDCx16_ASAP7_75t_R g473 ( .A(n_79), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_80), .B(n_176), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_81), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_82), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_83), .A2(n_146), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g446 ( .A(n_84), .Y(n_446) );
INVx2_ASAP7_75t_L g120 ( .A(n_85), .Y(n_120) );
INVx1_ASAP7_75t_L g435 ( .A(n_86), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_87), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_88), .B(n_162), .Y(n_225) );
OR2x2_ASAP7_75t_L g106 ( .A(n_89), .B(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g404 ( .A(n_89), .Y(n_404) );
OR2x2_ASAP7_75t_L g686 ( .A(n_89), .B(n_673), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_90), .A2(n_126), .B(n_141), .C(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_91), .B(n_146), .Y(n_171) );
INVx1_ASAP7_75t_L g175 ( .A(n_92), .Y(n_175) );
INVxp67_ASAP7_75t_L g252 ( .A(n_93), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_94), .B(n_118), .Y(n_427) );
INVx1_ASAP7_75t_L g132 ( .A(n_95), .Y(n_132) );
INVx1_ASAP7_75t_L g220 ( .A(n_96), .Y(n_220) );
INVx2_ASAP7_75t_L g417 ( .A(n_97), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_98), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g237 ( .A(n_99), .B(n_180), .Y(n_237) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_110), .B1(n_402), .B2(n_405), .Y(n_104) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_105), .A2(n_111), .B1(n_676), .B2(n_677), .Y(n_675) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g403 ( .A(n_107), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g673 ( .A(n_107), .Y(n_673) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
XNOR2xp5_ASAP7_75t_L g688 ( .A(n_111), .B(n_689), .Y(n_688) );
NAND2x1p5_ASAP7_75t_L g111 ( .A(n_112), .B(n_345), .Y(n_111) );
AND4x1_ASAP7_75t_L g112 ( .A(n_113), .B(n_285), .C(n_300), .D(n_325), .Y(n_112) );
NOR2xp33_ASAP7_75t_SL g113 ( .A(n_114), .B(n_258), .Y(n_113) );
OAI21xp33_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_166), .B(n_238), .Y(n_114) );
AND2x2_ASAP7_75t_L g288 ( .A(n_115), .B(n_184), .Y(n_288) );
AND2x2_ASAP7_75t_L g301 ( .A(n_115), .B(n_183), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_115), .B(n_167), .Y(n_351) );
INVx1_ASAP7_75t_L g355 ( .A(n_115), .Y(n_355) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_151), .Y(n_115) );
INVx2_ASAP7_75t_L g272 ( .A(n_116), .Y(n_272) );
BUFx2_ASAP7_75t_L g299 ( .A(n_116), .Y(n_299) );
AO21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_124), .B(n_149), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_117), .B(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g152 ( .A(n_117), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_117), .B(n_182), .Y(n_181) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_117), .A2(n_219), .B(n_226), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_117), .B(n_439), .Y(n_438) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_117), .A2(n_463), .B(n_469), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_117), .B(n_479), .Y(n_478) );
INVx4_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_118), .A2(n_206), .B(n_207), .Y(n_205) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_118), .Y(n_246) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g228 ( .A(n_119), .Y(n_228) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_120), .B(n_121), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_145), .Y(n_124) );
INVx5_ASAP7_75t_L g156 ( .A(n_126), .Y(n_156) );
AND2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_127), .Y(n_140) );
BUFx3_ASAP7_75t_L g164 ( .A(n_127), .Y(n_164) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g148 ( .A(n_128), .Y(n_148) );
INVx1_ASAP7_75t_L g214 ( .A(n_128), .Y(n_214) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_130), .Y(n_135) );
INVx3_ASAP7_75t_L g138 ( .A(n_130), .Y(n_138) );
AND2x2_ASAP7_75t_L g147 ( .A(n_130), .B(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_130), .Y(n_162) );
INVx1_ASAP7_75t_L g210 ( .A(n_130), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_136), .C(n_139), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_134), .B(n_417), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_134), .B(n_446), .Y(n_445) );
OAI22xp33_ASAP7_75t_L g492 ( .A1(n_134), .A2(n_137), .B1(n_493), .B2(n_494), .Y(n_492) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g177 ( .A(n_135), .Y(n_177) );
INVx2_ASAP7_75t_L g158 ( .A(n_137), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_137), .B(n_252), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_137), .A2(n_192), .B(n_476), .C(n_477), .Y(n_475) );
INVx5_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_138), .B(n_426), .Y(n_425) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g460 ( .A(n_140), .Y(n_460) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_SL g154 ( .A1(n_142), .A2(n_155), .B(n_156), .C(n_157), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_142), .A2(n_156), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g413 ( .A1(n_142), .A2(n_156), .B(n_414), .C(n_415), .Y(n_413) );
O2A1O1Ixp33_ASAP7_75t_SL g421 ( .A1(n_142), .A2(n_156), .B(n_422), .C(n_423), .Y(n_421) );
O2A1O1Ixp33_ASAP7_75t_SL g442 ( .A1(n_142), .A2(n_156), .B(n_443), .C(n_444), .Y(n_442) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_142), .A2(n_156), .B(n_456), .C(n_457), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_SL g489 ( .A1(n_142), .A2(n_156), .B(n_490), .C(n_491), .Y(n_489) );
INVx4_ASAP7_75t_SL g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g146 ( .A(n_143), .B(n_147), .Y(n_146) );
BUFx3_ASAP7_75t_L g194 ( .A(n_143), .Y(n_194) );
NAND2x1p5_ASAP7_75t_L g221 ( .A(n_143), .B(n_147), .Y(n_221) );
BUFx2_ASAP7_75t_L g187 ( .A(n_146), .Y(n_187) );
INVx1_ASAP7_75t_L g193 ( .A(n_148), .Y(n_193) );
AND2x2_ASAP7_75t_L g239 ( .A(n_151), .B(n_184), .Y(n_239) );
INVx2_ASAP7_75t_L g255 ( .A(n_151), .Y(n_255) );
AND2x2_ASAP7_75t_L g264 ( .A(n_151), .B(n_183), .Y(n_264) );
AND2x2_ASAP7_75t_L g343 ( .A(n_151), .B(n_272), .Y(n_343) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_165), .Y(n_151) );
INVx2_ASAP7_75t_L g173 ( .A(n_156), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_161), .B(n_459), .Y(n_458) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g424 ( .A(n_162), .Y(n_424) );
INVx2_ASAP7_75t_L g437 ( .A(n_163), .Y(n_437) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
INVx1_ASAP7_75t_L g447 ( .A(n_164), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_200), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_167), .B(n_270), .Y(n_308) );
INVx1_ASAP7_75t_L g396 ( .A(n_167), .Y(n_396) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_183), .Y(n_167) );
AND2x2_ASAP7_75t_L g254 ( .A(n_168), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g268 ( .A(n_168), .B(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_168), .Y(n_297) );
OR2x2_ASAP7_75t_L g329 ( .A(n_168), .B(n_271), .Y(n_329) );
AND2x2_ASAP7_75t_L g337 ( .A(n_168), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g370 ( .A(n_168), .B(n_339), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_168), .B(n_239), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_168), .B(n_299), .Y(n_395) );
AND2x2_ASAP7_75t_L g401 ( .A(n_168), .B(n_288), .Y(n_401) );
INVx5_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx2_ASAP7_75t_L g261 ( .A(n_169), .Y(n_261) );
AND2x2_ASAP7_75t_L g291 ( .A(n_169), .B(n_271), .Y(n_291) );
AND2x2_ASAP7_75t_L g324 ( .A(n_169), .B(n_284), .Y(n_324) );
AND2x2_ASAP7_75t_L g344 ( .A(n_169), .B(n_184), .Y(n_344) );
AND2x2_ASAP7_75t_L g378 ( .A(n_169), .B(n_244), .Y(n_378) );
OR2x6_ASAP7_75t_L g169 ( .A(n_170), .B(n_181), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_180), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_178), .C(n_179), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_176), .A2(n_179), .B(n_235), .C(n_236), .Y(n_234) );
O2A1O1Ixp5_ASAP7_75t_L g434 ( .A1(n_176), .A2(n_435), .B(n_436), .C(n_437), .Y(n_434) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_176), .A2(n_437), .B(n_467), .C(n_468), .Y(n_466) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g196 ( .A(n_180), .Y(n_196) );
INVx1_ASAP7_75t_L g199 ( .A(n_180), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_180), .A2(n_232), .B(n_233), .Y(n_231) );
OA21x2_ASAP7_75t_L g419 ( .A1(n_180), .A2(n_420), .B(n_427), .Y(n_419) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_180), .A2(n_221), .B(n_473), .C(n_474), .Y(n_472) );
AND2x4_ASAP7_75t_L g284 ( .A(n_183), .B(n_255), .Y(n_284) );
AND2x2_ASAP7_75t_L g295 ( .A(n_183), .B(n_291), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_183), .B(n_271), .Y(n_334) );
INVx2_ASAP7_75t_L g349 ( .A(n_183), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_183), .B(n_283), .Y(n_372) );
AND2x2_ASAP7_75t_L g391 ( .A(n_183), .B(n_343), .Y(n_391) );
INVx5_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_184), .Y(n_290) );
AND2x2_ASAP7_75t_L g298 ( .A(n_184), .B(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_L g339 ( .A(n_184), .B(n_255), .Y(n_339) );
OR2x6_ASAP7_75t_L g184 ( .A(n_185), .B(n_197), .Y(n_184) );
AOI21xp5_ASAP7_75t_SL g185 ( .A1(n_186), .A2(n_188), .B(n_195), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_192), .Y(n_189) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_193), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_196), .B(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
AO21x2_ASAP7_75t_L g430 ( .A1(n_199), .A2(n_431), .B(n_438), .Y(n_430) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_215), .Y(n_201) );
AND2x2_ASAP7_75t_L g262 ( .A(n_202), .B(n_245), .Y(n_262) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_203), .B(n_218), .Y(n_242) );
OR2x2_ASAP7_75t_L g275 ( .A(n_203), .B(n_245), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_203), .B(n_245), .Y(n_280) );
AND2x2_ASAP7_75t_L g307 ( .A(n_203), .B(n_244), .Y(n_307) );
AND2x2_ASAP7_75t_L g359 ( .A(n_203), .B(n_217), .Y(n_359) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_204), .B(n_229), .Y(n_267) );
AND2x2_ASAP7_75t_L g303 ( .A(n_204), .B(n_218), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_211), .B(n_212), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_212), .A2(n_224), .B(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_215), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_L g293 ( .A(n_216), .B(n_275), .Y(n_293) );
OR2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_229), .Y(n_216) );
OAI322xp33_ASAP7_75t_L g258 ( .A1(n_217), .A2(n_259), .A3(n_263), .B1(n_265), .B2(n_268), .C1(n_273), .C2(n_281), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_217), .B(n_244), .Y(n_266) );
OR2x2_ASAP7_75t_L g276 ( .A(n_217), .B(n_230), .Y(n_276) );
AND2x2_ASAP7_75t_L g278 ( .A(n_217), .B(n_230), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_217), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_217), .B(n_245), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_217), .B(n_374), .Y(n_373) );
INVx5_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_218), .B(n_262), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_222), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_221), .A2(n_432), .B(n_433), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_221), .A2(n_464), .B(n_465), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g487 ( .A(n_228), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_229), .B(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g256 ( .A(n_229), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_229), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g318 ( .A(n_229), .B(n_245), .Y(n_318) );
AOI211xp5_ASAP7_75t_SL g346 ( .A1(n_229), .A2(n_347), .B(n_350), .C(n_362), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_229), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g384 ( .A(n_229), .B(n_359), .Y(n_384) );
INVx5_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g312 ( .A(n_230), .B(n_245), .Y(n_312) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_230), .Y(n_321) );
AND2x2_ASAP7_75t_L g361 ( .A(n_230), .B(n_359), .Y(n_361) );
AND2x2_ASAP7_75t_SL g392 ( .A(n_230), .B(n_262), .Y(n_392) );
AND2x2_ASAP7_75t_L g399 ( .A(n_230), .B(n_358), .Y(n_399) );
OR2x6_ASAP7_75t_L g230 ( .A(n_231), .B(n_237), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B1(n_254), .B2(n_256), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_239), .B(n_261), .Y(n_309) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g257 ( .A(n_242), .Y(n_257) );
OR2x2_ASAP7_75t_L g317 ( .A(n_242), .B(n_318), .Y(n_317) );
OAI221xp5_ASAP7_75t_SL g365 ( .A1(n_242), .A2(n_366), .B1(n_368), .B2(n_369), .C(n_371), .Y(n_365) );
INVx2_ASAP7_75t_L g304 ( .A(n_243), .Y(n_304) );
AND2x2_ASAP7_75t_L g277 ( .A(n_244), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g367 ( .A(n_244), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_244), .B(n_359), .Y(n_380) );
INVx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVxp67_ASAP7_75t_L g322 ( .A(n_245), .Y(n_322) );
AND2x2_ASAP7_75t_L g358 ( .A(n_245), .B(n_359), .Y(n_358) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_253), .Y(n_245) );
OA21x2_ASAP7_75t_L g411 ( .A1(n_246), .A2(n_412), .B(n_418), .Y(n_411) );
OA21x2_ASAP7_75t_L g440 ( .A1(n_246), .A2(n_441), .B(n_448), .Y(n_440) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_246), .A2(n_454), .B(n_461), .Y(n_453) );
AND2x2_ASAP7_75t_L g360 ( .A(n_254), .B(n_299), .Y(n_360) );
AND2x2_ASAP7_75t_L g270 ( .A(n_255), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_255), .B(n_328), .Y(n_327) );
NOR2xp33_ASAP7_75t_SL g341 ( .A(n_257), .B(n_304), .Y(n_341) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g347 ( .A(n_260), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
OR2x2_ASAP7_75t_L g333 ( .A(n_261), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g398 ( .A(n_261), .B(n_343), .Y(n_398) );
INVx2_ASAP7_75t_L g331 ( .A(n_262), .Y(n_331) );
NAND4xp25_ASAP7_75t_SL g394 ( .A(n_263), .B(n_395), .C(n_396), .D(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_264), .B(n_328), .Y(n_363) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_SL g400 ( .A(n_267), .Y(n_400) );
O2A1O1Ixp33_ASAP7_75t_SL g362 ( .A1(n_268), .A2(n_331), .B(n_335), .C(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g357 ( .A(n_270), .B(n_349), .Y(n_357) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_271), .Y(n_283) );
INVx1_ASAP7_75t_L g338 ( .A(n_271), .Y(n_338) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_272), .Y(n_315) );
AOI211xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_276), .B(n_277), .C(n_279), .Y(n_273) );
AND2x2_ASAP7_75t_L g294 ( .A(n_274), .B(n_278), .Y(n_294) );
OAI322xp33_ASAP7_75t_SL g332 ( .A1(n_274), .A2(n_333), .A3(n_335), .B1(n_336), .B2(n_340), .C1(n_341), .C2(n_342), .Y(n_332) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g354 ( .A(n_276), .B(n_280), .Y(n_354) );
INVx1_ASAP7_75t_L g335 ( .A(n_278), .Y(n_335) );
INVx1_ASAP7_75t_SL g353 ( .A(n_280), .Y(n_353) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
AOI222xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_292), .B1(n_294), .B2(n_295), .C1(n_296), .C2(n_704), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_287), .B(n_289), .Y(n_286) );
OAI322xp33_ASAP7_75t_L g375 ( .A1(n_287), .A2(n_349), .A3(n_354), .B1(n_376), .B2(n_377), .C1(n_379), .C2(n_380), .Y(n_375) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_288), .A2(n_302), .B1(n_326), .B2(n_330), .C(n_332), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OAI222xp33_ASAP7_75t_L g305 ( .A1(n_293), .A2(n_306), .B1(n_308), .B2(n_309), .C1(n_310), .C2(n_313), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_295), .A2(n_302), .B1(n_372), .B2(n_373), .Y(n_371) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AOI211xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B(n_305), .C(n_316), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_L g381 ( .A1(n_302), .A2(n_339), .B(n_382), .C(n_385), .Y(n_381) );
AND2x4_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x2_ASAP7_75t_L g311 ( .A(n_303), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_SL g374 ( .A(n_307), .Y(n_374) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_314), .B(n_339), .Y(n_368) );
BUFx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI21xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_319), .B(n_323), .Y(n_316) );
OAI221xp5_ASAP7_75t_SL g385 ( .A1(n_317), .A2(n_386), .B1(n_387), .B2(n_388), .C(n_389), .Y(n_385) );
INVxp33_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_321), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_328), .B(n_339), .Y(n_379) );
INVx2_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AND2x2_ASAP7_75t_L g390 ( .A(n_343), .B(n_349), .Y(n_390) );
AND4x1_ASAP7_75t_L g345 ( .A(n_346), .B(n_364), .C(n_381), .D(n_393), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI221xp5_ASAP7_75t_SL g350 ( .A1(n_351), .A2(n_352), .B1(n_354), .B2(n_355), .C(n_356), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .B1(n_360), .B2(n_361), .Y(n_356) );
INVx1_ASAP7_75t_L g386 ( .A(n_357), .Y(n_386) );
INVx1_ASAP7_75t_SL g376 ( .A(n_361), .Y(n_376) );
NOR2xp33_ASAP7_75t_SL g364 ( .A(n_365), .B(n_375), .Y(n_364) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_377), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_384), .A2(n_390), .B1(n_391), .B2(n_392), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_399), .B1(n_400), .B2(n_401), .Y(n_393) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx6_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g676 ( .A(n_403), .Y(n_676) );
NOR2x2_ASAP7_75t_L g672 ( .A(n_404), .B(n_673), .Y(n_672) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g677 ( .A(n_406), .Y(n_677) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_592), .Y(n_406) );
NOR4xp25_ASAP7_75t_L g407 ( .A(n_408), .B(n_534), .C(n_564), .D(n_574), .Y(n_407) );
OAI211xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_449), .B(n_497), .C(n_524), .Y(n_408) );
OAI222xp33_ASAP7_75t_L g619 ( .A1(n_409), .A2(n_539), .B1(n_620), .B2(n_621), .C1(n_622), .C2(n_623), .Y(n_619) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_428), .Y(n_409) );
AOI33xp33_ASAP7_75t_L g545 ( .A1(n_410), .A2(n_532), .A3(n_533), .B1(n_546), .B2(n_551), .B3(n_553), .Y(n_545) );
OAI211xp5_ASAP7_75t_SL g602 ( .A1(n_410), .A2(n_603), .B(n_605), .C(n_607), .Y(n_602) );
OR2x2_ASAP7_75t_L g618 ( .A(n_410), .B(n_604), .Y(n_618) );
INVx1_ASAP7_75t_L g651 ( .A(n_410), .Y(n_651) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_419), .Y(n_410) );
INVx2_ASAP7_75t_L g528 ( .A(n_411), .Y(n_528) );
AND2x2_ASAP7_75t_L g544 ( .A(n_411), .B(n_440), .Y(n_544) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_411), .Y(n_579) );
AND2x2_ASAP7_75t_L g608 ( .A(n_411), .B(n_419), .Y(n_608) );
INVx2_ASAP7_75t_L g508 ( .A(n_419), .Y(n_508) );
BUFx3_ASAP7_75t_L g516 ( .A(n_419), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_419), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g527 ( .A(n_419), .B(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_419), .B(n_429), .Y(n_556) );
AND2x2_ASAP7_75t_L g625 ( .A(n_419), .B(n_559), .Y(n_625) );
INVx2_ASAP7_75t_SL g519 ( .A(n_428), .Y(n_519) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_440), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_429), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g561 ( .A(n_429), .Y(n_561) );
AND2x2_ASAP7_75t_L g572 ( .A(n_429), .B(n_528), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_429), .B(n_557), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_429), .B(n_559), .Y(n_604) );
AND2x2_ASAP7_75t_L g663 ( .A(n_429), .B(n_608), .Y(n_663) );
INVx4_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g533 ( .A(n_430), .B(n_440), .Y(n_533) );
AND2x2_ASAP7_75t_L g543 ( .A(n_430), .B(n_544), .Y(n_543) );
BUFx3_ASAP7_75t_L g565 ( .A(n_430), .Y(n_565) );
AND3x2_ASAP7_75t_L g624 ( .A(n_430), .B(n_625), .C(n_626), .Y(n_624) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_440), .Y(n_515) );
INVx1_ASAP7_75t_SL g559 ( .A(n_440), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_440), .B(n_508), .C(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_480), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g594 ( .A1(n_450), .A2(n_543), .B(n_595), .C(n_597), .Y(n_594) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_452), .B(n_471), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_452), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_SL g611 ( .A(n_452), .Y(n_611) );
AND2x2_ASAP7_75t_L g632 ( .A(n_452), .B(n_482), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_452), .B(n_541), .Y(n_660) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_462), .Y(n_452) );
AND2x2_ASAP7_75t_L g505 ( .A(n_453), .B(n_496), .Y(n_505) );
INVx2_ASAP7_75t_L g512 ( .A(n_453), .Y(n_512) );
AND2x2_ASAP7_75t_L g532 ( .A(n_453), .B(n_482), .Y(n_532) );
AND2x2_ASAP7_75t_L g582 ( .A(n_453), .B(n_471), .Y(n_582) );
INVx1_ASAP7_75t_L g586 ( .A(n_453), .Y(n_586) );
INVx2_ASAP7_75t_SL g496 ( .A(n_462), .Y(n_496) );
BUFx2_ASAP7_75t_L g522 ( .A(n_462), .Y(n_522) );
AND2x2_ASAP7_75t_L g649 ( .A(n_462), .B(n_471), .Y(n_649) );
INVx3_ASAP7_75t_SL g482 ( .A(n_471), .Y(n_482) );
AND2x2_ASAP7_75t_L g504 ( .A(n_471), .B(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_L g511 ( .A(n_471), .B(n_512), .Y(n_511) );
OR2x2_ASAP7_75t_L g541 ( .A(n_471), .B(n_501), .Y(n_541) );
OR2x2_ASAP7_75t_L g550 ( .A(n_471), .B(n_496), .Y(n_550) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_471), .Y(n_568) );
AND2x2_ASAP7_75t_L g573 ( .A(n_471), .B(n_526), .Y(n_573) );
AND2x2_ASAP7_75t_L g601 ( .A(n_471), .B(n_484), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_471), .B(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g639 ( .A(n_471), .B(n_483), .Y(n_639) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_478), .Y(n_471) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
AND2x2_ASAP7_75t_L g563 ( .A(n_482), .B(n_512), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_482), .B(n_505), .Y(n_591) );
AND2x2_ASAP7_75t_L g609 ( .A(n_482), .B(n_526), .Y(n_609) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_496), .Y(n_483) );
AND2x2_ASAP7_75t_L g510 ( .A(n_484), .B(n_496), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_484), .B(n_539), .Y(n_538) );
BUFx3_ASAP7_75t_L g548 ( .A(n_484), .Y(n_548) );
OR2x2_ASAP7_75t_L g596 ( .A(n_484), .B(n_516), .Y(n_596) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_488), .B(n_495), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_486), .A2(n_502), .B(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g502 ( .A(n_488), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_495), .Y(n_503) );
AND2x2_ASAP7_75t_L g531 ( .A(n_496), .B(n_501), .Y(n_531) );
INVx1_ASAP7_75t_L g539 ( .A(n_496), .Y(n_539) );
AND2x2_ASAP7_75t_L g634 ( .A(n_496), .B(n_512), .Y(n_634) );
AOI222xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_506), .B1(n_509), .B2(n_513), .C1(n_517), .C2(n_520), .Y(n_497) );
INVx1_ASAP7_75t_L g629 ( .A(n_498), .Y(n_629) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_504), .Y(n_498) );
AND2x2_ASAP7_75t_L g525 ( .A(n_499), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g536 ( .A(n_499), .B(n_505), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_499), .B(n_527), .Y(n_552) );
OAI222xp33_ASAP7_75t_L g574 ( .A1(n_499), .A2(n_575), .B1(n_580), .B2(n_581), .C1(n_589), .C2(n_591), .Y(n_574) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g562 ( .A(n_501), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_501), .B(n_582), .Y(n_622) );
AND2x2_ASAP7_75t_L g633 ( .A(n_501), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g641 ( .A(n_504), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_506), .B(n_557), .Y(n_620) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_508), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g578 ( .A(n_508), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx3_ASAP7_75t_L g523 ( .A(n_511), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_511), .A2(n_614), .B(n_617), .C(n_619), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_511), .B(n_548), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_511), .B(n_531), .Y(n_653) );
AND2x2_ASAP7_75t_L g526 ( .A(n_512), .B(n_522), .Y(n_526) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g553 ( .A(n_515), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_516), .B(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g605 ( .A(n_516), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g644 ( .A(n_516), .B(n_544), .Y(n_644) );
INVx1_ASAP7_75t_L g656 ( .A(n_516), .Y(n_656) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_519), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g637 ( .A(n_522), .Y(n_637) );
A2O1A1Ixp33_ASAP7_75t_SL g524 ( .A1(n_525), .A2(n_527), .B(n_529), .C(n_533), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_525), .A2(n_555), .B1(n_570), .B2(n_573), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_526), .B(n_540), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_526), .B(n_548), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_527), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_SL g590 ( .A(n_527), .Y(n_590) );
AND2x2_ASAP7_75t_L g597 ( .A(n_527), .B(n_577), .Y(n_597) );
INVx2_ASAP7_75t_L g558 ( .A(n_528), .Y(n_558) );
INVxp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
NOR4xp25_ASAP7_75t_L g535 ( .A(n_532), .B(n_536), .C(n_537), .D(n_540), .Y(n_535) );
INVx1_ASAP7_75t_SL g606 ( .A(n_533), .Y(n_606) );
AND2x2_ASAP7_75t_L g650 ( .A(n_533), .B(n_651), .Y(n_650) );
OAI211xp5_ASAP7_75t_SL g534 ( .A1(n_535), .A2(n_542), .B(n_545), .C(n_554), .Y(n_534) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_541), .B(n_611), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_543), .A2(n_662), .B1(n_663), .B2(n_664), .Y(n_661) );
INVx1_ASAP7_75t_SL g616 ( .A(n_544), .Y(n_616) );
AND2x2_ASAP7_75t_L g655 ( .A(n_544), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_548), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_552), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_553), .B(n_578), .Y(n_638) );
OAI21xp5_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_560), .B(n_562), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx1_ASAP7_75t_L g630 ( .A(n_557), .Y(n_630) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx2_ASAP7_75t_L g658 ( .A(n_558), .Y(n_658) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_559), .Y(n_585) );
OAI21xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B(n_569), .Y(n_564) );
CKINVDCx16_ASAP7_75t_R g577 ( .A(n_565), .Y(n_577) );
OR2x2_ASAP7_75t_L g615 ( .A(n_565), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AOI21xp33_ASAP7_75t_SL g610 ( .A1(n_568), .A2(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g598 ( .A1(n_572), .A2(n_599), .B1(n_602), .B2(n_609), .C(n_610), .Y(n_598) );
INVx1_ASAP7_75t_SL g642 ( .A(n_573), .Y(n_642) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
OR2x2_ASAP7_75t_L g589 ( .A(n_577), .B(n_590), .Y(n_589) );
INVxp67_ASAP7_75t_L g626 ( .A(n_579), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B1(n_586), .B2(n_587), .Y(n_581) );
INVx1_ASAP7_75t_L g621 ( .A(n_582), .Y(n_621) );
INVxp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_585), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NOR4xp25_ASAP7_75t_L g592 ( .A(n_593), .B(n_627), .C(n_640), .D(n_652), .Y(n_592) );
NAND3xp33_ASAP7_75t_SL g593 ( .A(n_594), .B(n_598), .C(n_613), .Y(n_593) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_596), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_603), .B(n_608), .Y(n_612) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI221xp5_ASAP7_75t_SL g640 ( .A1(n_615), .A2(n_641), .B1(n_642), .B2(n_643), .C(n_645), .Y(n_640) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_617), .A2(n_632), .B(n_633), .C(n_635), .Y(n_631) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_618), .A2(n_636), .B1(n_638), .B2(n_639), .Y(n_635) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B(n_630), .C(n_631), .Y(n_627) );
INVx1_ASAP7_75t_L g646 ( .A(n_639), .Y(n_646) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI21xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_647), .B(n_650), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI221xp5_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B1(n_657), .B2(n_659), .C(n_661), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
INVx3_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_684), .Y(n_679) );
NOR2xp33_ASAP7_75t_SL g680 ( .A(n_681), .B(n_683), .Y(n_680) );
INVx1_ASAP7_75t_SL g699 ( .A(n_681), .Y(n_699) );
INVx1_ASAP7_75t_L g698 ( .A(n_683), .Y(n_698) );
OA21x2_ASAP7_75t_L g701 ( .A1(n_683), .A2(n_699), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_686), .Y(n_693) );
INVx2_ASAP7_75t_L g695 ( .A(n_686), .Y(n_695) );
BUFx2_ASAP7_75t_L g702 ( .A(n_686), .Y(n_702) );
OAI21xp5_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_692), .B(n_694), .Y(n_687) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_701), .Y(n_700) );
endmodule