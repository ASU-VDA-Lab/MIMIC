module fake_jpeg_19352_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_2),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_21),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_74),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_62),
.Y(n_73)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_1),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_51),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_78),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_68),
.Y(n_92)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_68),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_66),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_59),
.B1(n_63),
.B2(n_53),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_77),
.B1(n_45),
.B2(n_67),
.Y(n_96)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_57),
.B1(n_71),
.B2(n_52),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_96),
.B1(n_102),
.B2(n_86),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_85),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_45),
.B(n_67),
.C(n_47),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_103),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_47),
.B1(n_56),
.B2(n_64),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_54),
.B1(n_69),
.B2(n_70),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_60),
.B1(n_66),
.B2(n_50),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_1),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_55),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_117),
.B1(n_7),
.B2(n_8),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_114),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_3),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_5),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_6),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_7),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_116),
.B(n_11),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_111),
.B1(n_117),
.B2(n_112),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_113),
.B1(n_14),
.B2(n_15),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_127),
.B1(n_119),
.B2(n_122),
.Y(n_131)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_108),
.A3(n_115),
.B1(n_104),
.B2(n_48),
.C1(n_20),
.C2(n_22),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.C(n_121),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_131),
.C(n_124),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_132),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_120),
.C(n_19),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_13),
.B(n_25),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_28),
.C(n_29),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_30),
.B(n_31),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_34),
.B(n_35),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_37),
.C(n_39),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_41),
.Y(n_141)
);


endmodule