module real_aes_15640_n_4 (n_0, n_3, n_2, n_1, n_4);
input n_0;
input n_3;
input n_2;
input n_1;
output n_4;
wire n_16;
wire n_17;
wire n_13;
wire n_18;
wire n_5;
wire n_15;
wire n_7;
wire n_8;
wire n_6;
wire n_12;
wire n_9;
wire n_14;
wire n_10;
wire n_11;
INVx1_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
BUFx3_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
INVx1_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
AND2x4_ASAP7_75t_L g14 ( .A(n_2), .B(n_7), .Y(n_14) );
INVx1_ASAP7_75t_L g7 ( .A(n_3), .Y(n_7) );
AOI21xp5_ASAP7_75t_L g12 ( .A1(n_3), .A2(n_13), .B(n_14), .Y(n_12) );
AOI21xp33_ASAP7_75t_SL g4 ( .A1(n_5), .A2(n_15), .B(n_16), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_6), .Y(n_5) );
AOI21xp33_ASAP7_75t_SL g6 ( .A1(n_7), .A2(n_8), .B(n_12), .Y(n_6) );
INVx3_ASAP7_75t_L g8 ( .A(n_9), .Y(n_8) );
BUFx8_ASAP7_75t_SL g9 ( .A(n_10), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
BUFx2_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
INVx2_ASAP7_75t_SL g17 ( .A(n_14), .Y(n_17) );
NOR3x1_ASAP7_75t_L g16 ( .A(n_15), .B(n_17), .C(n_18), .Y(n_16) );
endmodule