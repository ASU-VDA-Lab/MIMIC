module fake_jpeg_6190_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_27),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_10),
.B1(n_13),
.B2(n_17),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_34),
.B1(n_12),
.B2(n_19),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_13),
.B1(n_10),
.B2(n_17),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_10),
.B(n_13),
.C(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_33),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_32),
.B1(n_36),
.B2(n_38),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_19),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_20),
.B(n_18),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_26),
.B(n_22),
.C(n_28),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_45),
.B1(n_32),
.B2(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_48),
.Y(n_58)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_44),
.B1(n_48),
.B2(n_36),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_43),
.C(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_16),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

OAI32xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_39),
.A3(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_29),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_15),
.B1(n_14),
.B2(n_2),
.Y(n_72)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_68),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_64),
.Y(n_78)
);

AOI322xp5_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_54),
.A3(n_15),
.B1(n_14),
.B2(n_9),
.C1(n_4),
.C2(n_5),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_29),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_29),
.C(n_27),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_58),
.C(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_0),
.Y(n_75)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_66),
.C(n_60),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_1),
.B(n_3),
.C(n_6),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_75),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_14),
.B1(n_15),
.B2(n_9),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_1),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_76),
.C(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_78),
.C(n_69),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_75),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_83),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_92),
.B1(n_93),
.B2(n_83),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_82),
.C(n_14),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_61),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_97),
.Y(n_101)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_87),
.Y(n_102)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_99),
.A2(n_82),
.B1(n_14),
.B2(n_15),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_98),
.B1(n_91),
.B2(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_105),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_102),
.B1(n_99),
.B2(n_100),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_104),
.A2(n_101),
.B(n_100),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_105),
.C(n_6),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_15),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_107),
.Y(n_110)
);


endmodule