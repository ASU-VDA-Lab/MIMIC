module fake_jpeg_26726_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx8_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

CKINVDCx6p67_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_27),
.B1(n_19),
.B2(n_20),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_43),
.B1(n_50),
.B2(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_47),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_27),
.B1(n_19),
.B2(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_14),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_35),
.B1(n_30),
.B2(n_36),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_44),
.B1(n_41),
.B2(n_45),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_58),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_15),
.B1(n_41),
.B2(n_44),
.Y(n_74)
);

AOI32xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_33),
.A3(n_36),
.B1(n_17),
.B2(n_24),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_24),
.Y(n_68)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_61),
.Y(n_71)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_63),
.Y(n_76)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_65),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_57),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_28),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_74),
.B(n_75),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_37),
.A3(n_16),
.B1(n_23),
.B2(n_21),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_42),
.B(n_49),
.C(n_15),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_21),
.B(n_16),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_65),
.C(n_58),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_42),
.B1(n_49),
.B2(n_24),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_60),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_91),
.Y(n_99)
);

OA21x2_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_12),
.B(n_11),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_90),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_61),
.C(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_69),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_97),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_84),
.B1(n_74),
.B2(n_72),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_81),
.B1(n_82),
.B2(n_66),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_79),
.C(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_70),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_0),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_106),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_103),
.A2(n_72),
.B1(n_75),
.B2(n_80),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

XNOR2x2_ASAP7_75t_SL g109 ( 
.A(n_99),
.B(n_80),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_98),
.A3(n_95),
.B1(n_80),
.B2(n_0),
.C1(n_3),
.C2(n_1),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_5),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_107),
.A2(n_101),
.B1(n_99),
.B2(n_97),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_118),
.B1(n_119),
.B2(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_124),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_109),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_117),
.C(n_115),
.Y(n_127)
);

AOI31xp67_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_1),
.A3(n_6),
.B(n_9),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_115),
.B(n_6),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_125),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_130),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_126),
.Y(n_132)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_132),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);


endmodule