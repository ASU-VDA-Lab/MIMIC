module real_jpeg_465_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_2),
.A2(n_21),
.B1(n_35),
.B2(n_43),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_2),
.A2(n_26),
.B1(n_35),
.B2(n_47),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_2),
.A2(n_35),
.B1(n_58),
.B2(n_59),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_25),
.C(n_26),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_21),
.B1(n_37),
.B2(n_43),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_3),
.A2(n_26),
.B1(n_37),
.B2(n_47),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_3),
.A2(n_37),
.B1(n_58),
.B2(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_3),
.B(n_46),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_3),
.B(n_55),
.C(n_59),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_3),
.B(n_33),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_3),
.B(n_70),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_3),
.B(n_32),
.C(n_71),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_3),
.B(n_61),
.Y(n_162)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_108),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_10),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_112),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_111),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_91),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_15),
.B(n_91),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_65),
.C(n_82),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_16),
.A2(n_17),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_38),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_18),
.B(n_40),
.C(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_28),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_19),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_43),
.Y(n_45)
);

AO22x1_ASAP7_75t_SL g46 ( 
.A1(n_25),
.A2(n_26),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_26),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_26),
.A2(n_47),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_26),
.B(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_28),
.A2(n_29),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_29),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_29),
.B(n_150),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_29),
.B(n_110),
.C(n_162),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_30),
.B(n_36),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

AO22x1_ASAP7_75t_L g70 ( 
.A1(n_31),
.A2(n_32),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_32),
.B(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_34),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_36),
.B(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_50),
.B2(n_64),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_46),
.B2(n_49),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OA21x2_ASAP7_75t_L g88 ( 
.A1(n_42),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_50),
.B(n_124),
.C(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_50),
.A2(n_64),
.B1(n_130),
.B2(n_133),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_61),
.B2(n_62),
.Y(n_50)
);

AO21x1_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_61),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_63),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_57),
.B(n_63),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

AOI22x1_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_59),
.B1(n_71),
.B2(n_72),
.Y(n_73)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_59),
.B(n_155),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_65),
.A2(n_82),
.B1(n_83),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_65),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_76),
.B2(n_77),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_77),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_66),
.A2(n_67),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_66),
.B(n_156),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_66),
.A2(n_67),
.B1(n_84),
.B2(n_120),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_66),
.B(n_84),
.C(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_69),
.B(n_74),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_68),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_80),
.B(n_81),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_80),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_80),
.A2(n_81),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_80),
.B(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.C(n_87),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_86),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_88),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_88),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_102),
.B2(n_103),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_109),
.A2(n_110),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_109),
.A2(n_110),
.B1(n_134),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_129),
.C(n_134),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_179),
.B(n_186),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_141),
.B(n_178),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_128),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_128),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_117),
.B(n_123),
.C(n_127),
.Y(n_181)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_125),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_153),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_172),
.B(n_177),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_166),
.B(n_171),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_158),
.B(n_165),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_152),
.B(n_157),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_149),
.B(n_151),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_154),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_164),
.Y(n_165)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_168),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_176),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_182),
.Y(n_186)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);


endmodule