module fake_jpeg_22511_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_7),
.B(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_41),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_26),
.C(n_27),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_28),
.C(n_24),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_46),
.Y(n_65)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_55),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_21),
.B1(n_16),
.B2(n_23),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_57),
.B1(n_64),
.B2(n_31),
.Y(n_73)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_25),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_18),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_29),
.B1(n_25),
.B2(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_63),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_70),
.C(n_3),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_69),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_40),
.A2(n_24),
.B(n_32),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_86),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_83),
.B1(n_49),
.B2(n_58),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_19),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_85),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_30),
.B1(n_34),
.B2(n_32),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_2),
.Y(n_84)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_9),
.B(n_14),
.C(n_13),
.D(n_11),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_3),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_65),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_9),
.B(n_14),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_34),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_3),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_99),
.B1(n_79),
.B2(n_77),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_49),
.B(n_57),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_104),
.C(n_106),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_49),
.B1(n_52),
.B2(n_56),
.Y(n_99)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_56),
.B(n_5),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_69),
.C(n_63),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_75),
.C(n_92),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_62),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_118),
.Y(n_119)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_116),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_127),
.B1(n_132),
.B2(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_88),
.B1(n_84),
.B2(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_83),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_136),
.C(n_138),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_86),
.B1(n_80),
.B2(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_135),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_78),
.B1(n_90),
.B2(n_80),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_103),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_75),
.C(n_71),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_104),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_144),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_101),
.Y(n_143)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_137),
.A2(n_71),
.B1(n_116),
.B2(n_113),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_139),
.B(n_141),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_148),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_117),
.B(n_102),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_136),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_101),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_110),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_151),
.B(n_156),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

AO221x1_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_125),
.B1(n_140),
.B2(n_141),
.C(n_144),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_115),
.B1(n_111),
.B2(n_108),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_154),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_124),
.C(n_138),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_163),
.C(n_165),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_151),
.Y(n_159)
);

BUFx24_ASAP7_75t_SL g176 ( 
.A(n_159),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_161),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_134),
.C(n_128),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_142),
.B(n_133),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_120),
.C(n_111),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_148),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g175 ( 
.A(n_170),
.B(n_149),
.CI(n_142),
.CON(n_175),
.SN(n_175)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_172),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_174),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_155),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_SL g181 ( 
.A(n_175),
.B(n_178),
.C(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_139),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_177),
.A2(n_164),
.B(n_158),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_184),
.C(n_176),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_149),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_188),
.Y(n_191)
);

OAI21x1_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_156),
.B(n_162),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_11),
.B(n_13),
.C(n_7),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_163),
.C(n_120),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_87),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_87),
.B1(n_93),
.B2(n_62),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_183),
.B(n_185),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_192),
.B(n_194),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_180),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_193),
.C(n_6),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_4),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_6),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_78),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_78),
.B(n_8),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_200),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_195),
.B(n_8),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);


endmodule