module fake_jpeg_14902_n_293 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2x1_ASAP7_75t_SL g38 ( 
.A(n_20),
.B(n_1),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_20),
.CON(n_58),
.SN(n_58)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_14),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_17),
.Y(n_57)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_16),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_38),
.B1(n_15),
.B2(n_30),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_38),
.B(n_26),
.Y(n_77)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_48),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_16),
.B1(n_37),
.B2(n_21),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_37),
.B1(n_25),
.B2(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_29),
.B1(n_19),
.B2(n_46),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_32),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_64),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_79),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_38),
.B1(n_23),
.B2(n_26),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_81),
.B1(n_67),
.B2(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_33),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_77),
.B(n_18),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_83),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_42),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_50),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_44),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_100),
.B(n_73),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_44),
.B(n_28),
.Y(n_90)
);

OR2x4_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_28),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_29),
.B(n_25),
.C(n_15),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_95),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_107),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_101),
.B1(n_109),
.B2(n_113),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_65),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_70),
.B(n_32),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_74),
.A2(n_54),
.B1(n_53),
.B2(n_43),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_61),
.B1(n_55),
.B2(n_59),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_110),
.B1(n_83),
.B2(n_114),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_87),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_43),
.B1(n_55),
.B2(n_50),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_50),
.B1(n_19),
.B2(n_26),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_85),
.B1(n_76),
.B2(n_82),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_130),
.B(n_134),
.Y(n_159)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_85),
.B1(n_62),
.B2(n_71),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_66),
.B(n_84),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_93),
.C(n_88),
.Y(n_155)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_76),
.B1(n_78),
.B2(n_82),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_127),
.B1(n_92),
.B2(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_131),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_86),
.B(n_42),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_133),
.B(n_136),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_75),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_99),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_111),
.B(n_114),
.C(n_99),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_89),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_1),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_80),
.C(n_41),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_153),
.C(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_148),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_98),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_152),
.B(n_155),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_98),
.B1(n_105),
.B2(n_90),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_147),
.A2(n_157),
.B1(n_116),
.B2(n_127),
.Y(n_169)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_97),
.Y(n_151)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_93),
.B(n_104),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_89),
.Y(n_153)
);

OAI22x1_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_132),
.B1(n_111),
.B2(n_116),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_88),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_125),
.B1(n_132),
.B2(n_133),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_91),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_120),
.A3(n_136),
.B1(n_123),
.B2(n_138),
.C1(n_132),
.C2(n_119),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_118),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_164),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_91),
.B1(n_111),
.B2(n_94),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_35),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_111),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_118),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_184),
.B(n_166),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_168),
.A2(n_185),
.B1(n_150),
.B2(n_160),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_189),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_141),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_170),
.B(n_178),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_139),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_174),
.C(n_175),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_131),
.B1(n_134),
.B2(n_130),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_180),
.B1(n_183),
.B2(n_149),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_134),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_130),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_103),
.B1(n_99),
.B2(n_117),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_41),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_150),
.C(n_163),
.Y(n_202)
);

NOR2x1_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_126),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_146),
.A2(n_126),
.B1(n_117),
.B2(n_87),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_145),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_146),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_159),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_193),
.B(n_194),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_179),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_203),
.B(n_211),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_182),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_197),
.B(n_195),
.Y(n_220)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_206),
.B1(n_208),
.B2(n_210),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_212),
.C(n_181),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_188),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_209),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_149),
.B1(n_152),
.B2(n_165),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_207),
.A2(n_189),
.B1(n_154),
.B2(n_169),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_168),
.A2(n_143),
.B1(n_158),
.B2(n_154),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_154),
.B1(n_156),
.B2(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_162),
.C(n_126),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_204),
.B(n_87),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_177),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_223),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_226),
.C(n_228),
.Y(n_234)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_176),
.B1(n_172),
.B2(n_154),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_224),
.B1(n_200),
.B2(n_193),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_171),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_174),
.B1(n_175),
.B2(n_14),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_126),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_229),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_198),
.C(n_210),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_80),
.C(n_18),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_48),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_48),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_208),
.C(n_196),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_203),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_235),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_201),
.Y(n_233)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_236),
.Y(n_257)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_228),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_191),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_240),
.B(n_242),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_229),
.A2(n_211),
.B(n_207),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_217),
.C(n_225),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_204),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_1),
.B(n_2),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_22),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_245),
.B(n_22),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_255),
.C(n_28),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_253),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_213),
.B1(n_223),
.B2(n_216),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_241),
.B1(n_234),
.B2(n_243),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_213),
.B(n_11),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_251),
.A2(n_13),
.B(n_12),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_232),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_13),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_234),
.C(n_243),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_2),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_242),
.B(n_240),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_252),
.B(n_247),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_263),
.Y(n_273)
);

AOI21x1_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_238),
.B(n_12),
.Y(n_261)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_267),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_270)
);

AO21x1_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_264),
.B(n_265),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_13),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_268),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_2),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_22),
.Y(n_268)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_277),
.B1(n_5),
.B2(n_7),
.Y(n_280)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_275),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_250),
.A3(n_255),
.B1(n_26),
.B2(n_23),
.C1(n_17),
.C2(n_9),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_5),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_265),
.A3(n_17),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_277)
);

AOI31xp33_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_5),
.A3(n_7),
.B(n_8),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_279),
.B1(n_282),
.B2(n_277),
.Y(n_285)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_273),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_18),
.C(n_22),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_18),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_285),
.Y(n_289)
);

AO21x1_ASAP7_75t_L g290 ( 
.A1(n_286),
.A2(n_287),
.B(n_288),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_284),
.A2(n_8),
.B(n_9),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_18),
.C(n_22),
.Y(n_288)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_9),
.A3(n_10),
.B1(n_22),
.B2(n_285),
.C1(n_280),
.C2(n_283),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_291),
.B(n_290),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_292),
.Y(n_293)
);


endmodule