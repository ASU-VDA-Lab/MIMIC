module real_aes_3109_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_564;
wire n_519;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_601;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g288 ( .A(n_0), .B(n_268), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_1), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_2), .A2(n_64), .B1(n_159), .B2(n_160), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_SL g340 ( .A1(n_3), .A2(n_213), .B(n_341), .C(n_342), .Y(n_340) );
OAI22xp33_ASAP7_75t_L g293 ( .A1(n_4), .A2(n_63), .B1(n_211), .B2(n_240), .Y(n_293) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_5), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_6), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_7), .A2(n_51), .B1(n_238), .B2(n_240), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_8), .Y(n_259) );
INVx1_ASAP7_75t_L g106 ( .A(n_9), .Y(n_106) );
INVxp67_ASAP7_75t_L g116 ( .A(n_9), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_9), .B(n_54), .Y(n_137) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_10), .A2(n_38), .B1(n_145), .B2(n_149), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_11), .A2(n_43), .B1(n_211), .B2(n_236), .Y(n_235) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_12), .A2(n_50), .B(n_226), .Y(n_225) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_12), .A2(n_50), .B(n_226), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g102 ( .A(n_13), .B(n_91), .Y(n_102) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_14), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_15), .Y(n_314) );
BUFx3_ASAP7_75t_L g183 ( .A(n_16), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g346 ( .A1(n_17), .A2(n_294), .B(n_347), .C(n_348), .Y(n_346) );
OAI22xp33_ASAP7_75t_SL g291 ( .A1(n_18), .A2(n_32), .B1(n_211), .B2(n_258), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_19), .A2(n_24), .B1(n_258), .B2(n_263), .Y(n_278) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_20), .Y(n_91) );
O2A1O1Ixp5_ASAP7_75t_L g206 ( .A1(n_21), .A2(n_207), .B(n_210), .C(n_213), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_22), .A2(n_56), .B1(n_162), .B2(n_163), .Y(n_161) );
INVx1_ASAP7_75t_L g95 ( .A(n_23), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_23), .B(n_53), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_25), .A2(n_29), .B1(n_119), .B2(n_121), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_26), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_27), .A2(n_52), .B1(n_151), .B2(n_156), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_28), .B(n_284), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_30), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g86 ( .A1(n_31), .A2(n_41), .B1(n_87), .B2(n_109), .Y(n_86) );
INVx1_ASAP7_75t_L g226 ( .A(n_33), .Y(n_226) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_34), .Y(n_194) );
AND2x4_ASAP7_75t_L g222 ( .A(n_34), .B(n_192), .Y(n_222) );
AND2x4_ASAP7_75t_L g243 ( .A(n_34), .B(n_192), .Y(n_243) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_35), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_36), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_37), .Y(n_81) );
INVx2_ASAP7_75t_L g264 ( .A(n_39), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g316 ( .A1(n_40), .A2(n_213), .B(n_317), .C(n_318), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_42), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_44), .A2(n_60), .B1(n_280), .B2(n_281), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_45), .B(n_244), .Y(n_306) );
OA22x2_ASAP7_75t_L g89 ( .A1(n_46), .A2(n_54), .B1(n_90), .B2(n_91), .Y(n_89) );
INVx1_ASAP7_75t_L g126 ( .A(n_46), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_47), .A2(n_71), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_48), .Y(n_305) );
NAND2xp33_ASAP7_75t_R g245 ( .A(n_49), .B(n_230), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_49), .A2(n_76), .B1(n_284), .B2(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g108 ( .A(n_53), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_53), .B(n_124), .Y(n_140) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_53), .Y(n_186) );
OAI21xp33_ASAP7_75t_L g127 ( .A1(n_54), .A2(n_61), .B(n_117), .Y(n_127) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_55), .Y(n_172) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_57), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_58), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_59), .Y(n_260) );
INVx1_ASAP7_75t_L g97 ( .A(n_61), .Y(n_97) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_61), .B(n_73), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_62), .B(n_142), .Y(n_141) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_65), .Y(n_209) );
BUFx5_ASAP7_75t_L g211 ( .A(n_65), .Y(n_211) );
INVx1_ASAP7_75t_L g239 ( .A(n_65), .Y(n_239) );
INVx2_ASAP7_75t_L g352 ( .A(n_66), .Y(n_352) );
INVx2_ASAP7_75t_L g321 ( .A(n_67), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_68), .A2(n_82), .B1(n_83), .B2(n_606), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_68), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_69), .Y(n_349) );
INVx2_ASAP7_75t_SL g192 ( .A(n_70), .Y(n_192) );
INVx1_ASAP7_75t_L g218 ( .A(n_72), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g100 ( .A(n_73), .B(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g228 ( .A(n_74), .Y(n_228) );
OAI21xp33_ASAP7_75t_SL g312 ( .A1(n_75), .A2(n_211), .B(n_313), .Y(n_312) );
INVxp67_ASAP7_75t_SL g266 ( .A(n_76), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_76), .B(n_284), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_178), .B1(n_195), .B2(n_591), .C(n_598), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_165), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_82), .B1(n_83), .B2(n_164), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_80), .Y(n_164) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_81), .B(n_211), .Y(n_219) );
AOI22xp5_ASAP7_75t_SL g599 ( .A1(n_82), .A2(n_83), .B1(n_600), .B2(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
OR2x2_ASAP7_75t_L g84 ( .A(n_85), .B(n_143), .Y(n_84) );
NAND4xp25_ASAP7_75t_L g85 ( .A(n_86), .B(n_118), .C(n_130), .D(n_141), .Y(n_85) );
AND2x4_ASAP7_75t_L g87 ( .A(n_88), .B(n_98), .Y(n_87) );
AND2x2_ASAP7_75t_L g131 ( .A(n_88), .B(n_128), .Y(n_131) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_92), .Y(n_88) );
AND2x2_ASAP7_75t_L g114 ( .A(n_89), .B(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g120 ( .A(n_89), .B(n_93), .Y(n_120) );
INVx1_ASAP7_75t_L g153 ( .A(n_89), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g96 ( .A(n_90), .B(n_97), .Y(n_96) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
NAND2xp33_ASAP7_75t_L g94 ( .A(n_91), .B(n_95), .Y(n_94) );
INVx3_ASAP7_75t_L g101 ( .A(n_91), .Y(n_101) );
NAND2xp33_ASAP7_75t_L g107 ( .A(n_91), .B(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_91), .Y(n_112) );
INVx1_ASAP7_75t_L g117 ( .A(n_91), .Y(n_117) );
AND2x4_ASAP7_75t_L g152 ( .A(n_92), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g93 ( .A(n_94), .B(n_96), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_95), .B(n_126), .Y(n_125) );
INVxp67_ASAP7_75t_L g187 ( .A(n_95), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g115 ( .A1(n_97), .A2(n_116), .B(n_117), .Y(n_115) );
AND2x4_ASAP7_75t_L g119 ( .A(n_98), .B(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g162 ( .A(n_98), .B(n_152), .Y(n_162) );
AND2x4_ASAP7_75t_L g98 ( .A(n_99), .B(n_103), .Y(n_98) );
AND2x2_ASAP7_75t_L g110 ( .A(n_99), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g129 ( .A(n_99), .Y(n_129) );
OR2x2_ASAP7_75t_L g147 ( .A(n_99), .B(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g154 ( .A(n_99), .B(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_102), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_101), .B(n_106), .Y(n_105) );
INVxp67_ASAP7_75t_L g124 ( .A(n_101), .Y(n_124) );
NAND3xp33_ASAP7_75t_L g139 ( .A(n_102), .B(n_123), .C(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g128 ( .A(n_103), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g148 ( .A(n_104), .Y(n_148) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_114), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g135 ( .A(n_112), .Y(n_135) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_113), .Y(n_184) );
AND2x2_ASAP7_75t_L g142 ( .A(n_120), .B(n_128), .Y(n_142) );
AND2x4_ASAP7_75t_L g145 ( .A(n_120), .B(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g159 ( .A(n_120), .B(n_154), .Y(n_159) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_128), .Y(n_121) );
AND2x4_ASAP7_75t_L g149 ( .A(n_122), .B(n_146), .Y(n_149) );
AND2x4_ASAP7_75t_L g160 ( .A(n_122), .B(n_154), .Y(n_160) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_127), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_126), .Y(n_188) );
AND2x4_ASAP7_75t_L g163 ( .A(n_128), .B(n_152), .Y(n_163) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_139), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
NAND4xp25_ASAP7_75t_L g143 ( .A(n_144), .B(n_150), .C(n_158), .D(n_161), .Y(n_143) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g157 ( .A(n_147), .Y(n_157) );
INVx1_ASAP7_75t_L g155 ( .A(n_148), .Y(n_155) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_154), .Y(n_151) );
AND2x4_ASAP7_75t_L g156 ( .A(n_152), .B(n_157), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B1(n_176), .B2(n_177), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_166), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_167), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B1(n_170), .B2(n_171), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B1(n_174), .B2(n_175), .Y(n_171) );
INVx1_ASAP7_75t_L g174 ( .A(n_172), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_173), .Y(n_175) );
BUFx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_189), .Y(n_180) );
INVxp67_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g603 ( .A(n_182), .B(n_189), .Y(n_603) );
AOI211xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_185), .C(n_188), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_193), .Y(n_189) );
OR2x2_ASAP7_75t_L g608 ( .A(n_190), .B(n_194), .Y(n_608) );
INVx1_ASAP7_75t_L g611 ( .A(n_190), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_190), .B(n_193), .Y(n_612) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND4x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_449), .C(n_489), .D(n_558), .Y(n_198) );
NOR2x1_ASAP7_75t_L g199 ( .A(n_200), .B(n_387), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_201), .B(n_367), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_246), .B(n_270), .C(n_322), .Y(n_201) );
AND2x2_ASAP7_75t_L g381 ( .A(n_202), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_202), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g435 ( .A(n_202), .Y(n_435) );
AND2x2_ASAP7_75t_L g455 ( .A(n_202), .B(n_324), .Y(n_455) );
AND2x2_ASAP7_75t_L g557 ( .A(n_202), .B(n_538), .Y(n_557) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_231), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_203), .B(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g583 ( .A(n_203), .B(n_522), .Y(n_583) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g354 ( .A(n_204), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g361 ( .A(n_204), .Y(n_361) );
BUFx2_ASAP7_75t_R g421 ( .A(n_204), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_204), .B(n_338), .Y(n_530) );
AND2x2_ASAP7_75t_L g534 ( .A(n_204), .B(n_337), .Y(n_534) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_223), .B(n_227), .Y(n_204) );
NOR3xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_215), .C(n_221), .Y(n_205) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g216 ( .A(n_208), .Y(n_216) );
INVx1_ASAP7_75t_L g317 ( .A(n_208), .Y(n_317) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g236 ( .A(n_209), .Y(n_236) );
INVx2_ASAP7_75t_L g240 ( .A(n_209), .Y(n_240) );
INVx6_ASAP7_75t_L g258 ( .A(n_209), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_211), .A2(n_258), .B1(n_259), .B2(n_260), .Y(n_257) );
AOI22xp33_ASAP7_75t_SL g300 ( .A1(n_211), .A2(n_258), .B1(n_301), .B2(n_302), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_211), .A2(n_236), .B1(n_304), .B2(n_305), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_211), .B(n_314), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_213), .A2(n_220), .B1(n_235), .B2(n_237), .Y(n_234) );
OAI22xp33_ASAP7_75t_L g256 ( .A1(n_213), .A2(n_220), .B1(n_257), .B2(n_261), .Y(n_256) );
OAI221xp5_ASAP7_75t_L g299 ( .A1(n_213), .A2(n_243), .B1(n_294), .B2(n_300), .C(n_303), .Y(n_299) );
INVx1_ASAP7_75t_L g380 ( .A(n_213), .Y(n_380) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_214), .B(n_218), .Y(n_217) );
INVx4_ASAP7_75t_L g220 ( .A(n_214), .Y(n_220) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_214), .Y(n_277) );
INVx1_ASAP7_75t_L g282 ( .A(n_214), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_214), .B(n_291), .Y(n_290) );
INVx3_ASAP7_75t_L g294 ( .A(n_214), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B1(n_219), .B2(n_220), .Y(n_215) );
INVx2_ASAP7_75t_L g315 ( .A(n_220), .Y(n_315) );
NOR2xp33_ASAP7_75t_SL g350 ( .A(n_221), .B(n_268), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_221), .A2(n_315), .B1(n_378), .B2(n_379), .C(n_380), .Y(n_377) );
INVx4_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_222), .B(n_254), .Y(n_275) );
AND2x2_ASAP7_75t_L g309 ( .A(n_222), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_223), .B(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx3_ASAP7_75t_L g244 ( .A(n_224), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_224), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx4_ASAP7_75t_L g269 ( .A(n_225), .Y(n_269) );
BUFx3_ASAP7_75t_L g331 ( .A(n_225), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
BUFx3_ASAP7_75t_L g255 ( .A(n_230), .Y(n_255) );
INVx1_ASAP7_75t_L g310 ( .A(n_230), .Y(n_310) );
INVx2_ASAP7_75t_L g508 ( .A(n_230), .Y(n_508) );
INVx1_ASAP7_75t_SL g248 ( .A(n_231), .Y(n_248) );
INVx1_ASAP7_75t_L g362 ( .A(n_231), .Y(n_362) );
AND2x2_ASAP7_75t_L g444 ( .A(n_231), .B(n_337), .Y(n_444) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g355 ( .A(n_232), .Y(n_355) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_232), .Y(n_371) );
AND2x2_ASAP7_75t_L g459 ( .A(n_232), .B(n_361), .Y(n_459) );
AND2x2_ASAP7_75t_L g531 ( .A(n_232), .B(n_251), .Y(n_531) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_245), .Y(n_232) );
AND2x2_ASAP7_75t_L g505 ( .A(n_233), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_241), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_236), .A2(n_262), .B1(n_263), .B2(n_264), .Y(n_261) );
INVx1_ASAP7_75t_L g347 ( .A(n_236), .Y(n_347) );
INVx2_ASAP7_75t_L g280 ( .A(n_238), .Y(n_280) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g263 ( .A(n_239), .Y(n_263) );
NOR2xp67_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_243), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_243), .B(n_269), .Y(n_295) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_249), .B(n_353), .Y(n_580) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x4_ASAP7_75t_L g446 ( .A(n_251), .B(n_338), .Y(n_446) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_256), .B(n_265), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x2_ASAP7_75t_SL g592 ( .A(n_253), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g378 ( .A(n_257), .Y(n_378) );
INVx2_ASAP7_75t_SL g281 ( .A(n_258), .Y(n_281) );
INVx2_ASAP7_75t_L g343 ( .A(n_258), .Y(n_343) );
INVx1_ASAP7_75t_L g600 ( .A(n_260), .Y(n_600) );
INVx1_ASAP7_75t_L g379 ( .A(n_261), .Y(n_379) );
INVx1_ASAP7_75t_L g614 ( .A(n_262), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_263), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_263), .B(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g298 ( .A(n_267), .Y(n_298) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g284 ( .A(n_269), .Y(n_284) );
NOR2xp33_ASAP7_75t_SL g351 ( .A(n_269), .B(n_352), .Y(n_351) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_285), .Y(n_271) );
AND2x4_ASAP7_75t_L g364 ( .A(n_272), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g448 ( .A(n_273), .B(n_417), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_273), .B(n_442), .Y(n_461) );
OR2x2_ASAP7_75t_L g565 ( .A(n_273), .B(n_521), .Y(n_565) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g401 ( .A(n_274), .Y(n_401) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B(n_283), .Y(n_274) );
INVx1_ASAP7_75t_L g329 ( .A(n_276), .Y(n_329) );
OA22x2_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B1(n_279), .B2(n_282), .Y(n_276) );
INVx4_ASAP7_75t_L g597 ( .A(n_277), .Y(n_597) );
INVx1_ASAP7_75t_L g341 ( .A(n_280), .Y(n_341) );
INVx1_ASAP7_75t_L g332 ( .A(n_283), .Y(n_332) );
BUFx2_ASAP7_75t_SL g429 ( .A(n_285), .Y(n_429) );
NOR2xp67_ASAP7_75t_L g285 ( .A(n_286), .B(n_296), .Y(n_285) );
INVx1_ASAP7_75t_L g384 ( .A(n_286), .Y(n_384) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g366 ( .A(n_287), .Y(n_366) );
INVx3_ASAP7_75t_L g403 ( .A(n_287), .Y(n_403) );
AND2x2_ASAP7_75t_L g438 ( .A(n_287), .B(n_404), .Y(n_438) );
AND2x2_ASAP7_75t_L g468 ( .A(n_287), .B(n_307), .Y(n_468) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B(n_295), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_307), .Y(n_296) );
INVx2_ASAP7_75t_L g333 ( .A(n_297), .Y(n_333) );
INVx2_ASAP7_75t_L g386 ( .A(n_297), .Y(n_386) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_306), .Y(n_297) );
OA21x2_ASAP7_75t_L g404 ( .A1(n_298), .A2(n_299), .B(n_306), .Y(n_404) );
INVx1_ASAP7_75t_L g325 ( .A(n_307), .Y(n_325) );
AND2x2_ASAP7_75t_L g385 ( .A(n_307), .B(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g411 ( .A(n_307), .B(n_366), .Y(n_411) );
INVx2_ASAP7_75t_L g417 ( .A(n_307), .Y(n_417) );
AND2x2_ASAP7_75t_L g442 ( .A(n_307), .B(n_403), .Y(n_442) );
BUFx2_ASAP7_75t_L g511 ( .A(n_307), .Y(n_511) );
INVx2_ASAP7_75t_L g522 ( .A(n_307), .Y(n_522) );
INVx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI21x1_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_311), .B(n_320), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .B(n_316), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_334), .B1(n_356), .B2(n_363), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g423 ( .A(n_327), .B(n_416), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_327), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_SL g517 ( .A(n_327), .Y(n_517) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_333), .Y(n_327) );
OR2x2_ASAP7_75t_L g409 ( .A(n_328), .B(n_404), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B(n_332), .Y(n_328) );
INVx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g365 ( .A(n_333), .B(n_366), .Y(n_365) );
NAND3xp33_ASAP7_75t_L g389 ( .A(n_334), .B(n_390), .C(n_394), .Y(n_389) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_353), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g372 ( .A(n_336), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g382 ( .A(n_338), .B(n_374), .Y(n_382) );
INVx1_ASAP7_75t_L g393 ( .A(n_338), .Y(n_393) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_338), .Y(n_397) );
OR2x2_ASAP7_75t_L g426 ( .A(n_338), .B(n_374), .Y(n_426) );
INVx1_ASAP7_75t_L g463 ( .A(n_338), .Y(n_463) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_338), .Y(n_585) );
AO31x2_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_345), .A3(n_350), .B(n_351), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_347), .Y(n_594) );
OR2x2_ASAP7_75t_L g412 ( .A(n_353), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g424 ( .A(n_354), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g433 ( .A(n_354), .B(n_382), .Y(n_433) );
AND2x4_ASAP7_75t_L g469 ( .A(n_354), .B(n_446), .Y(n_469) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g514 ( .A(n_359), .B(n_397), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_360), .B(n_374), .Y(n_554) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_361), .Y(n_488) );
AND2x2_ASAP7_75t_L g539 ( .A(n_361), .B(n_504), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_363), .B(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g546 ( .A(n_364), .B(n_499), .Y(n_546) );
NAND2x1p5_ASAP7_75t_L g510 ( .A(n_365), .B(n_511), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g556 ( .A(n_365), .B(n_551), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_365), .B(n_448), .Y(n_569) );
AND2x2_ASAP7_75t_L g431 ( .A(n_366), .B(n_401), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_381), .B(n_383), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
AND2x2_ASAP7_75t_L g391 ( .A(n_370), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_370), .B(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g472 ( .A(n_370), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_370), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g518 ( .A(n_372), .Y(n_518) );
INVx1_ASAP7_75t_L g589 ( .A(n_373), .Y(n_589) );
AND2x2_ASAP7_75t_L g392 ( .A(n_374), .B(n_393), .Y(n_392) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_374), .Y(n_478) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
AND2x2_ASAP7_75t_L g504 ( .A(n_376), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_382), .B(n_421), .Y(n_420) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_382), .Y(n_525) );
AOI22xp5_ASAP7_75t_SL g464 ( .A1(n_383), .A2(n_465), .B1(n_466), .B2(n_469), .Y(n_464) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_422), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_398), .B(n_405), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g436 ( .A(n_392), .Y(n_436) );
OR2x2_ASAP7_75t_L g502 ( .A(n_393), .B(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g574 ( .A(n_393), .B(n_531), .Y(n_574) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_394), .Y(n_465) );
BUFx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVxp67_ASAP7_75t_L g413 ( .A(n_396), .Y(n_413) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_399), .A2(n_468), .B(n_471), .C(n_474), .Y(n_470) );
OR2x2_ASAP7_75t_L g543 ( .A(n_399), .B(n_411), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_399), .B(n_402), .Y(n_577) );
AND2x2_ASAP7_75t_L g590 ( .A(n_399), .B(n_438), .Y(n_590) );
INVx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g498 ( .A(n_400), .B(n_402), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_400), .B(n_438), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_400), .B(n_442), .Y(n_561) );
AND2x2_ASAP7_75t_L g566 ( .A(n_400), .B(n_468), .Y(n_566) );
INVx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g454 ( .A(n_401), .Y(n_454) );
AND2x2_ASAP7_75t_L g572 ( .A(n_401), .B(n_404), .Y(n_572) );
AND2x2_ASAP7_75t_L g479 ( .A(n_402), .B(n_448), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_402), .B(n_511), .Y(n_542) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_403), .B(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g453 ( .A(n_404), .B(n_454), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_412), .B1(n_414), .B2(n_418), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
AND2x2_ASAP7_75t_L g415 ( .A(n_408), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_408), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g440 ( .A(n_409), .Y(n_440) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g499 ( .A(n_416), .Y(n_499) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g482 ( .A(n_417), .B(n_431), .Y(n_482) );
AND2x2_ASAP7_75t_L g484 ( .A(n_417), .B(n_438), .Y(n_484) );
INVx1_ASAP7_75t_L g552 ( .A(n_417), .Y(n_552) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_419), .A2(n_557), .B1(n_564), .B2(n_566), .Y(n_563) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g494 ( .A(n_421), .Y(n_494) );
AOI211xp5_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_424), .B(n_427), .C(n_434), .Y(n_422) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_424), .B(n_528), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_425), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B(n_432), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI332xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .A3(n_437), .B1(n_439), .B2(n_441), .B3(n_443), .C1(n_445), .C2(n_447), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_438), .A2(n_528), .B1(n_532), .B2(n_533), .Y(n_527) );
INVxp67_ASAP7_75t_SL g532 ( .A(n_439), .Y(n_532) );
INVx2_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g587 ( .A(n_441), .Y(n_587) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g553 ( .A(n_444), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g588 ( .A(n_444), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_SL g473 ( .A(n_446), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_446), .B(n_459), .Y(n_474) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND4x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_464), .C(n_470), .D(n_475), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_455), .B(n_456), .C(n_462), .Y(n_450) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
OAI321xp33_ASAP7_75t_L g578 ( .A1(n_452), .A2(n_519), .A3(n_532), .B1(n_579), .B2(n_581), .C(n_586), .Y(n_578) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVxp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_SL g538 ( .A(n_463), .Y(n_538) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_473), .A2(n_481), .B(n_483), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_479), .B(n_480), .C(n_485), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVxp67_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_484), .A2(n_501), .B1(n_509), .B2(n_512), .Y(n_500) );
INVxp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_490), .B(n_526), .Y(n_489) );
OAI211xp5_ASAP7_75t_SL g490 ( .A1(n_491), .A2(n_495), .B(n_500), .C(n_515), .Y(n_490) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
OR2x2_ASAP7_75t_L g570 ( .A(n_499), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_502), .B(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g584 ( .A(n_503), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g545 ( .A(n_504), .Y(n_545) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AOI32xp33_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_518), .A3(n_519), .B1(n_520), .B2(n_523), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND3xp33_ASAP7_75t_SL g526 ( .A(n_527), .B(n_535), .C(n_547), .Y(n_526) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g533 ( .A(n_531), .B(n_534), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_531), .A2(n_587), .B1(n_588), .B2(n_590), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_540), .B1(n_544), .B2(n_546), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2x1p5_ASAP7_75t_SL g537 ( .A(n_538), .B(n_539), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .C(n_543), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_543), .A2(n_560), .B(n_562), .C(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_553), .B1(n_555), .B2(n_557), .Y(n_547) );
BUFx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NOR3xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_567), .C(n_578), .Y(n_558) );
BUFx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_570), .B(n_573), .C(n_575), .Y(n_567) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVxp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NOR2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
BUFx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OA21x2_ASAP7_75t_L g610 ( .A1(n_593), .A2(n_611), .B(n_612), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_596), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI222xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_602), .B1(n_604), .B2(n_607), .C1(n_609), .C2(n_613), .Y(n_598) );
INVx1_ASAP7_75t_L g601 ( .A(n_600), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
BUFx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
endmodule