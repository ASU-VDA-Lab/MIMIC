module fake_jpeg_6038_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx9p33_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_26),
.B1(n_23),
.B2(n_15),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_52),
.B1(n_56),
.B2(n_62),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_18),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_60),
.B(n_45),
.C(n_31),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_15),
.B1(n_23),
.B2(n_26),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_26),
.B1(n_15),
.B2(n_23),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_20),
.B1(n_18),
.B2(n_30),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_20),
.B1(n_28),
.B2(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_32),
.B(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_17),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_25),
.B1(n_18),
.B2(n_24),
.Y(n_62)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_31),
.B1(n_40),
.B2(n_37),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_65),
.A2(n_20),
.B1(n_54),
.B2(n_53),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_70),
.Y(n_92)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_42),
.C(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_80),
.B(n_82),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVxp67_ASAP7_75t_SL g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_89),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_99),
.B1(n_81),
.B2(n_72),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_47),
.B1(n_54),
.B2(n_62),
.Y(n_99)
);

AO22x2_ASAP7_75t_L g100 ( 
.A1(n_65),
.A2(n_61),
.B1(n_58),
.B2(n_39),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_66),
.B1(n_75),
.B2(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_119),
.B1(n_92),
.B2(n_87),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_81),
.C(n_72),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_120),
.C(n_92),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_101),
.B1(n_100),
.B2(n_67),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_106),
.A2(n_123),
.B1(n_34),
.B2(n_53),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_114),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_66),
.B1(n_89),
.B2(n_101),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_117),
.Y(n_131)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_67),
.B1(n_54),
.B2(n_46),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_77),
.C(n_43),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_85),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_39),
.B1(n_34),
.B2(n_43),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_84),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_134),
.C(n_135),
.Y(n_151)
);

XOR2x1_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_106),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_145),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_118),
.B1(n_95),
.B2(n_94),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_145),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_136),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_91),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_77),
.C(n_90),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_137),
.B(n_144),
.Y(n_162)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_143),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_61),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_86),
.C(n_53),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_98),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_141),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_88),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_120),
.C(n_112),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_51),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

XOR2x2_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_140),
.Y(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_112),
.B(n_118),
.C(n_121),
.D(n_115),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_156),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_139),
.B1(n_142),
.B2(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_103),
.Y(n_154)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_122),
.B(n_17),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_161),
.B(n_136),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_163),
.C(n_141),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_22),
.B1(n_16),
.B2(n_19),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_22),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_128),
.A2(n_51),
.B(n_71),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_51),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_166),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_179),
.B1(n_163),
.B2(n_148),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_162),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_172),
.B(n_165),
.Y(n_189)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_174),
.B(n_176),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_171),
.C(n_151),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_144),
.C(n_51),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_69),
.B(n_73),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_149),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_173),
.B(n_174),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_73),
.B1(n_19),
.B2(n_16),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_172),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_167),
.B1(n_177),
.B2(n_178),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_187),
.B1(n_21),
.B2(n_22),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_148),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_185),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_168),
.B(n_158),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_191),
.B(n_175),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_147),
.B1(n_159),
.B2(n_157),
.Y(n_187)
);

NAND2x1_ASAP7_75t_SL g199 ( 
.A(n_189),
.B(n_22),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_171),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_176),
.A2(n_0),
.B(n_1),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_164),
.B(n_1),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_179),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_200),
.B1(n_202),
.B2(n_187),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_197),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_29),
.B(n_19),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_181),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_198),
.A2(n_201),
.B1(n_4),
.B2(n_5),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_199),
.A2(n_29),
.B1(n_8),
.B2(n_9),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_3),
.B(n_4),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_189),
.A2(n_22),
.B1(n_19),
.B2(n_16),
.Y(n_201)
);

OAI21x1_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_188),
.B(n_183),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_207),
.C(n_202),
.Y(n_212)
);

OAI221xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_180),
.B1(n_191),
.B2(n_184),
.C(n_29),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_208),
.Y(n_214)
);

AOI31xp33_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_16),
.A3(n_29),
.B(n_6),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_5),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_213),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_5),
.B1(n_10),
.B2(n_12),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_194),
.C(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_10),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_216),
.A2(n_210),
.B1(n_8),
.B2(n_10),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_219),
.C(n_12),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_218),
.A2(n_214),
.B(n_215),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_14),
.C(n_12),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_223),
.B(n_217),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_225),
.C(n_13),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_13),
.B(n_215),
.Y(n_227)
);


endmodule