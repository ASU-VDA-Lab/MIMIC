module fake_jpeg_16955_n_141 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_13),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_21),
.A2(n_0),
.B1(n_2),
.B2(n_6),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_7),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_13),
.B(n_2),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_28),
.B(n_24),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AO21x1_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_48),
.B(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_15),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_31),
.A2(n_30),
.B1(n_34),
.B2(n_33),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_27),
.B(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_15),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_29),
.B(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_21),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_8),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_78),
.B1(n_79),
.B2(n_10),
.Y(n_82)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_53),
.B1(n_59),
.B2(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_75),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_27),
.B1(n_19),
.B2(n_24),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_26),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_10),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_16),
.B1(n_22),
.B2(n_12),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_16),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_59),
.Y(n_94)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_91),
.Y(n_101)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_51),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_72),
.B1(n_79),
.B2(n_63),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_66),
.Y(n_96)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_73),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_64),
.B(n_70),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_107),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_87),
.B(n_85),
.C(n_82),
.D(n_78),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_111),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_88),
.C(n_77),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_94),
.C(n_65),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_114),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_103),
.B1(n_99),
.B2(n_97),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_83),
.C(n_62),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_83),
.C(n_62),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_116),
.B(n_97),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_121),
.C(n_84),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_124),
.B(n_106),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_113),
.B(n_84),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_129),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_127),
.B(n_128),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_128),
.A2(n_122),
.B(n_120),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_130),
.A2(n_131),
.B(n_104),
.Y(n_136)
);

NOR2xp67_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_121),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_104),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_86),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_136),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_81),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_138),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_140),
.Y(n_141)
);


endmodule