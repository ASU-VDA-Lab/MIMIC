module fake_jpeg_16761_n_359 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_359);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_359;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g19 ( 
.A(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_47),
.Y(n_57)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_0),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_32),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_26),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_37),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_22),
.B1(n_37),
.B2(n_26),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_71),
.B1(n_78),
.B2(n_20),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_33),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_64),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_22),
.B1(n_35),
.B2(n_36),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_67),
.B1(n_80),
.B2(n_29),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_28),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_35),
.B1(n_33),
.B2(n_21),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_35),
.B1(n_26),
.B2(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_72),
.B(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_41),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_32),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_79),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_75),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_27),
.C(n_30),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_39),
.B1(n_38),
.B2(n_34),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_32),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_20),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_86),
.B(n_95),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_91),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_90),
.A2(n_114),
.B1(n_25),
.B2(n_63),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_38),
.B1(n_34),
.B2(n_21),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_74),
.Y(n_116)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_21),
.B1(n_25),
.B2(n_29),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_104),
.B1(n_105),
.B2(n_85),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_112),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_51),
.B1(n_48),
.B2(n_46),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_51),
.B1(n_48),
.B2(n_44),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_64),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_29),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_57),
.Y(n_130)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_77),
.A2(n_25),
.B1(n_27),
.B2(n_10),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_122),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_141),
.B1(n_145),
.B2(n_95),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_59),
.Y(n_122)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_126),
.B1(n_143),
.B2(n_92),
.Y(n_156)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_130),
.B(n_12),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_79),
.C(n_73),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_134),
.C(n_86),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_57),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_81),
.C(n_69),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_70),
.Y(n_137)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_70),
.Y(n_139)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_109),
.B(n_69),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_144),
.B(n_121),
.Y(n_150)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_101),
.A2(n_77),
.B1(n_63),
.B2(n_85),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_88),
.A2(n_66),
.B1(n_63),
.B2(n_58),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_153),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_88),
.B1(n_66),
.B2(n_104),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_149),
.B1(n_155),
.B2(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_95),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_157),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_87),
.B(n_27),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_162),
.B(n_166),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_87),
.C(n_55),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_99),
.B1(n_94),
.B2(n_96),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_87),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_110),
.B1(n_103),
.B2(n_105),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_116),
.A2(n_108),
.B1(n_102),
.B2(n_13),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_159),
.A2(n_160),
.B1(n_125),
.B2(n_143),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_12),
.B1(n_18),
.B2(n_17),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_128),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_141),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_163),
.B(n_17),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_119),
.B(n_126),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_27),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_169),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_115),
.B(n_0),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_75),
.B(n_1),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_169),
.B(n_167),
.Y(n_184)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_149),
.A2(n_117),
.B1(n_124),
.B2(n_136),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_179),
.A2(n_190),
.B1(n_159),
.B2(n_150),
.Y(n_211)
);

OAI22x1_ASAP7_75t_SL g180 ( 
.A1(n_158),
.A2(n_135),
.B1(n_138),
.B2(n_123),
.Y(n_180)
);

OAI22x1_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_194),
.B1(n_135),
.B2(n_123),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_184),
.A2(n_192),
.B(n_166),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_185),
.B(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_170),
.B(n_136),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_124),
.B1(n_118),
.B2(n_140),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_161),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_173),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_123),
.B(n_1),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_152),
.A2(n_127),
.B1(n_135),
.B2(n_138),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_162),
.B1(n_147),
.B2(n_146),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_197),
.A2(n_200),
.B1(n_213),
.B2(n_195),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_162),
.B1(n_146),
.B2(n_152),
.Y(n_200)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_174),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_206),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_153),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_207),
.C(n_172),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_153),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_217),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_214),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_189),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_151),
.B(n_157),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_209),
.B(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_154),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_219),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_220),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_180),
.B(n_160),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_197),
.B(n_175),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_232),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_217),
.A2(n_183),
.B1(n_180),
.B2(n_186),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_225),
.A2(n_240),
.B1(n_204),
.B2(n_208),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_175),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_229),
.C(n_230),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_184),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_231),
.B(n_238),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_172),
.C(n_178),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_183),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_235),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_179),
.C(n_148),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_198),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_212),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_212),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_243),
.A2(n_246),
.B(n_208),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_203),
.C(n_211),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_226),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_176),
.Y(n_245)
);

XOR2x2_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_249),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_191),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_248),
.Y(n_251)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_227),
.B(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_210),
.Y(n_256)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_256),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_261),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_222),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_260),
.A2(n_272),
.B1(n_262),
.B2(n_264),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_222),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_265),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_263),
.B(n_128),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_236),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_264),
.A2(n_267),
.B(n_270),
.Y(n_278)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_204),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_244),
.B(n_185),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_271),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_232),
.C(n_230),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_239),
.B(n_223),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_247),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_235),
.B1(n_241),
.B2(n_224),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_274),
.A2(n_270),
.B1(n_254),
.B2(n_261),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_281),
.C(n_282),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_229),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_286),
.Y(n_304)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_228),
.C(n_246),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_240),
.C(n_225),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_128),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_123),
.C(n_127),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_292),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_257),
.B(n_265),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_257),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_251),
.B(n_11),
.Y(n_291)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_30),
.C(n_54),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_300),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_284),
.Y(n_296)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_254),
.B1(n_267),
.B2(n_259),
.Y(n_297)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_308),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_257),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_302),
.A2(n_303),
.B(n_307),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_289),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_278),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_283),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_2),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_288),
.C(n_276),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_317),
.C(n_319),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_300),
.B(n_263),
.CI(n_274),
.CON(n_312),
.SN(n_312)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_295),
.A2(n_290),
.B1(n_282),
.B2(n_272),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_6),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_277),
.C(n_292),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_296),
.C(n_281),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_302),
.A2(n_278),
.B(n_250),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_321),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_256),
.C(n_287),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_280),
.C(n_260),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_311),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_306),
.B1(n_303),
.B2(n_3),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_329),
.C(n_333),
.Y(n_341)
);

FAx1_ASAP7_75t_SL g326 ( 
.A(n_310),
.B(n_10),
.CI(n_16),
.CON(n_326),
.SN(n_326)
);

FAx1_ASAP7_75t_SL g343 ( 
.A(n_326),
.B(n_10),
.CI(n_14),
.CON(n_343),
.SN(n_343)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_0),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_9),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_316),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_332),
.Y(n_338)
);

O2A1O1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_331),
.A2(n_334),
.B(n_317),
.C(n_312),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_321),
.A2(n_2),
.B1(n_6),
.B2(n_9),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_335),
.B(n_336),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_318),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_339),
.Y(n_346)
);

AOI21x1_ASAP7_75t_L g339 ( 
.A1(n_326),
.A2(n_309),
.B(n_14),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_324),
.A2(n_309),
.B(n_14),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_340),
.B(n_342),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_30),
.C(n_54),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_343),
.B(n_326),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_336),
.A2(n_323),
.B(n_328),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_344),
.A2(n_338),
.B(n_332),
.Y(n_352)
);

BUFx24_ASAP7_75t_SL g347 ( 
.A(n_343),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_347),
.B(n_349),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_345),
.B(n_333),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_351),
.B(n_352),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_350),
.C(n_348),
.Y(n_354)
);

AOI21x1_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_346),
.B(n_341),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_335),
.B(n_330),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_356),
.A2(n_15),
.B(n_16),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_15),
.C(n_16),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_15),
.B(n_75),
.Y(n_359)
);


endmodule