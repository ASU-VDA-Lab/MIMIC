module fake_jpeg_29671_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx8_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

AOI21xp33_ASAP7_75t_L g12 ( 
.A1(n_7),
.A2(n_0),
.B(n_2),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_1),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_24),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_2),
.B(n_3),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_20),
.A2(n_14),
.B1(n_8),
.B2(n_11),
.Y(n_36)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx4_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_20),
.B(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_17),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_21),
.B(n_13),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_39),
.C(n_41),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_10),
.B(n_23),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_15),
.C(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_46),
.B1(n_23),
.B2(n_39),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_47),
.B1(n_41),
.B2(n_17),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_51),
.C(n_47),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_50),
.A2(n_30),
.B(n_13),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_32),
.C(n_34),
.Y(n_51)
);

NOR2xp67_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_51),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_30),
.B1(n_27),
.B2(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_55),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_18),
.B1(n_22),
.B2(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_13),
.Y(n_59)
);


endmodule