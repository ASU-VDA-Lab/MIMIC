module fake_jpeg_1870_n_199 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_199);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_3),
.B(n_24),
.C(n_15),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_67),
.Y(n_73)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_62),
.Y(n_81)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_1),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_72),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_3),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_52),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_59),
.B1(n_61),
.B2(n_56),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_45),
.B1(n_61),
.B2(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_53),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_83),
.B(n_84),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_45),
.B1(n_46),
.B2(n_62),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_51),
.B1(n_68),
.B2(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_81),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_63),
.B(n_53),
.C(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_100),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_50),
.B1(n_51),
.B2(n_46),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_80),
.B1(n_82),
.B2(n_75),
.Y(n_103)
);

NAND2x1_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_56),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_75),
.B(n_64),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_55),
.B(n_57),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_64),
.B(n_58),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_95),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_57),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_42),
.B1(n_39),
.B2(n_38),
.Y(n_118)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_47),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_83),
.C(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_109),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_109),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_82),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_108),
.A2(n_112),
.B(n_8),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_89),
.B1(n_88),
.B2(n_90),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_118),
.B1(n_5),
.B2(n_6),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_47),
.C(n_64),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_115),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_4),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_100),
.C(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_117),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_4),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_37),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_36),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_131),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_128),
.A2(n_139),
.B(n_9),
.Y(n_149)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_35),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_118),
.B1(n_114),
.B2(n_12),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_104),
.B(n_7),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_136),
.Y(n_159)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_8),
.Y(n_136)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_9),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_108),
.C(n_114),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_146),
.C(n_126),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_33),
.C(n_30),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_123),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_147),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_149),
.A2(n_131),
.B(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_155),
.B1(n_16),
.B2(n_17),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_121),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_14),
.B(n_15),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_132),
.B(n_137),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_164),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_127),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_171),
.C(n_146),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_169),
.B1(n_173),
.B2(n_157),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_138),
.B(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_153),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_28),
.C(n_27),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_158),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_172),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_179),
.Y(n_188)
);

AOI221xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_150),
.B1(n_145),
.B2(n_141),
.C(n_159),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_182),
.B(n_160),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_162),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_148),
.B1(n_144),
.B2(n_18),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_180),
.B(n_178),
.Y(n_184)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_16),
.A3(n_17),
.B1(n_18),
.B2(n_19),
.C1(n_20),
.C2(n_21),
.Y(n_182)
);

AOI31xp33_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_185),
.A3(n_161),
.B(n_177),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_179),
.B1(n_181),
.B2(n_167),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_163),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_176),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_191),
.Y(n_192)
);

NOR2xp67_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_171),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_191),
.C(n_192),
.Y(n_194)
);

O2A1O1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_194),
.A2(n_188),
.B(n_184),
.C(n_167),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_187),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_166),
.B(n_20),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_19),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_26),
.Y(n_199)
);


endmodule