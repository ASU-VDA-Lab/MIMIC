module fake_netlist_6_316_n_6181 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_625, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_644, n_621, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_648, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_612, n_633, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_110, n_151, n_412, n_640, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_364, n_637, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_171, n_192, n_57, n_169, n_51, n_649, n_283, n_6181);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_625;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_648;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_612;
input n_633;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_364;
input n_637;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_6181;

wire n_5643;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_741;
wire n_1351;
wire n_5254;
wire n_1212;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_6141;
wire n_3849;
wire n_5138;
wire n_4395;
wire n_4388;
wire n_1061;
wire n_3089;
wire n_783;
wire n_5653;
wire n_4978;
wire n_5409;
wire n_5301;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_1387;
wire n_3222;
wire n_677;
wire n_6126;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_5524;
wire n_5345;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_5818;
wire n_2179;
wire n_5963;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_5950;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5548;
wire n_5057;
wire n_3030;
wire n_830;
wire n_5838;
wire n_5725;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_5900;
wire n_4273;
wire n_5545;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_5598;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_5819;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_5279;
wire n_2786;
wire n_5894;
wire n_5930;
wire n_5239;
wire n_1781;
wire n_1971;
wire n_5354;
wire n_5332;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_5908;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_5420;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_6015;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_5638;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_6110;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_5684;
wire n_5729;
wire n_5680;
wire n_6148;
wire n_686;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_5522;
wire n_5828;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_5902;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_6107;
wire n_2832;
wire n_4226;
wire n_5493;
wire n_1762;
wire n_1910;
wire n_3980;
wire n_1075;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_5452;
wire n_3888;
wire n_6151;
wire n_764;
wire n_5476;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_5536;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_6055;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_5532;
wire n_5897;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_5609;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_5922;
wire n_2641;
wire n_5658;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_5667;
wire n_780;
wire n_2624;
wire n_5865;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_5281;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_5314;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_3968;
wire n_2096;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_5795;
wire n_4473;
wire n_6043;
wire n_5552;
wire n_5226;
wire n_687;
wire n_890;
wire n_5457;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_6010;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4289;
wire n_4288;
wire n_3763;
wire n_2712;
wire n_5529;
wire n_3733;
wire n_6042;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_5957;
wire n_4228;
wire n_3423;
wire n_1932;
wire n_925;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_2767;
wire n_4576;
wire n_5929;
wire n_4615;
wire n_5787;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_5445;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_5501;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_6033;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_5748;
wire n_3782;
wire n_6097;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_5870;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_5636;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_989;
wire n_2689;
wire n_1473;
wire n_5286;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_5811;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_705;
wire n_1004;
wire n_1529;
wire n_5530;
wire n_2473;
wire n_5397;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_5595;
wire n_3119;
wire n_5427;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_5388;
wire n_4718;
wire n_1448;
wire n_5901;
wire n_5962;
wire n_3631;
wire n_5599;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_5326;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_6149;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_1398;
wire n_1201;
wire n_884;
wire n_5394;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_5359;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_5741;
wire n_2773;
wire n_5405;
wire n_5288;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_5952;
wire n_3964;
wire n_2416;
wire n_5947;
wire n_1877;
wire n_3944;
wire n_6124;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_5985;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_5761;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_5760;
wire n_2146;
wire n_2131;
wire n_5472;
wire n_3547;
wire n_5679;
wire n_2575;
wire n_5100;
wire n_5973;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_5688;
wire n_5740;
wire n_1731;
wire n_5820;
wire n_5648;
wire n_2135;
wire n_5745;
wire n_4707;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_5180;
wire n_2049;
wire n_858;
wire n_5182;
wire n_956;
wire n_5534;
wire n_663;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_664;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_5949;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_6100;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_5906;
wire n_1934;
wire n_5660;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_5334;
wire n_6024;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_5783;
wire n_3120;
wire n_5821;
wire n_6079;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_5556;
wire n_4932;
wire n_5456;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_5500;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_6059;
wire n_3042;
wire n_6065;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_5433;
wire n_6075;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_6117;
wire n_5618;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_6133;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_5978;
wire n_4996;
wire n_4990;
wire n_5247;
wire n_6127;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_6006;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_5689;
wire n_1043;
wire n_4090;
wire n_6115;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_6048;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_5931;
wire n_2371;
wire n_6139;
wire n_1361;
wire n_662;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_5641;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_6085;
wire n_5731;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_5883;
wire n_5754;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_5629;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_6147;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_5434;
wire n_5934;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_6157;
wire n_4859;
wire n_2626;
wire n_5880;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_5852;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_5960;
wire n_4571;
wire n_3698;
wire n_5358;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_6073;
wire n_1484;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_5571;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_5512;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_6025;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_5607;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_5999;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_6150;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_695;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_5562;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_5911;
wire n_2122;
wire n_5622;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_5577;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_698;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_5413;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_5915;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_5779;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_3617;
wire n_2076;
wire n_6019;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_6036;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_5591;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_6013;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_5518;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_5847;
wire n_6049;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2444;
wire n_2437;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_668;
wire n_4166;
wire n_1821;
wire n_6136;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_6091;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_5541;
wire n_5568;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_5381;
wire n_2408;
wire n_5723;
wire n_5918;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_5696;
wire n_4486;
wire n_1816;
wire n_6131;
wire n_5848;
wire n_3024;
wire n_4612;
wire n_5673;
wire n_5443;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_5485;
wire n_5823;
wire n_2800;
wire n_3496;
wire n_5473;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_5537;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_3288;
wire n_2918;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_6137;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_5630;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_5379;
wire n_5335;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_6113;
wire n_2634;
wire n_1761;
wire n_5424;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_5505;
wire n_5868;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_5018;
wire n_6129;
wire n_3815;
wire n_3896;
wire n_5274;
wire n_3274;
wire n_5401;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_5989;
wire n_4928;
wire n_5769;
wire n_4794;
wire n_722;
wire n_5613;
wire n_5612;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_5581;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_5375;
wire n_2451;
wire n_5370;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_5601;
wire n_5784;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_5248;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_5635;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_5528;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_873;
wire n_3946;
wire n_2989;
wire n_5778;
wire n_3395;
wire n_4474;
wire n_5665;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_6135;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_5788;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_6168;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_666;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_5317;
wire n_1094;
wire n_5430;
wire n_5942;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_5540;
wire n_3532;
wire n_5716;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_5762;
wire n_6132;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_6179;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_659;
wire n_3351;
wire n_6171;
wire n_808;
wire n_5519;
wire n_4047;
wire n_5753;
wire n_3413;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_6083;
wire n_3164;
wire n_4575;
wire n_699;
wire n_4320;
wire n_3884;
wire n_5808;
wire n_5436;
wire n_5139;
wire n_757;
wire n_5231;
wire n_2190;
wire n_6120;
wire n_6068;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_5789;
wire n_2104;
wire n_3883;
wire n_5961;
wire n_5866;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5822;
wire n_5195;
wire n_6121;
wire n_3949;
wire n_5726;
wire n_2792;
wire n_5364;
wire n_3315;
wire n_5533;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_4107;
wire n_1876;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_5953;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_5718;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_6001;
wire n_3686;
wire n_4502;
wire n_5958;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_5792;
wire n_3581;
wire n_3069;
wire n_6023;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_5554;
wire n_1175;
wire n_2311;
wire n_3691;
wire n_1012;
wire n_5553;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_5711;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_5790;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_4004;
wire n_2206;
wire n_2967;
wire n_5404;
wire n_2916;
wire n_5739;
wire n_4292;
wire n_6163;
wire n_5972;
wire n_2467;
wire n_5549;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_3280;
wire n_5757;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_701;
wire n_950;
wire n_3009;
wire n_5824;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_5488;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_5637;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_5728;
wire n_5471;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_5843;
wire n_2078;
wire n_2932;
wire n_3431;
wire n_1767;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_5484;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_5523;
wire n_1067;
wire n_3405;
wire n_5423;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_3442;
wire n_1880;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_5204;
wire n_5333;
wire n_847;
wire n_682;
wire n_851;
wire n_4991;
wire n_5594;
wire n_2554;
wire n_5422;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_5526;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_5551;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_3133;
wire n_1959;
wire n_5257;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4753;
wire n_4688;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_5887;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_5631;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_6008;
wire n_1022;
wire n_5854;
wire n_2667;
wire n_5460;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_5686;
wire n_5899;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_5981;
wire n_3788;
wire n_4891;
wire n_5937;
wire n_777;
wire n_1299;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_6040;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5465;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_6160;
wire n_796;
wire n_1195;
wire n_1811;
wire n_3987;
wire n_1857;
wire n_1519;
wire n_6039;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_5721;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_5719;
wire n_1502;
wire n_5773;
wire n_1659;
wire n_5482;
wire n_3393;
wire n_6012;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_6064;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_5793;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_5578;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_3718;
wire n_5893;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5742;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_5676;
wire n_1220;
wire n_6051;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_5674;
wire n_3270;
wire n_5539;
wire n_2846;
wire n_5282;
wire n_970;
wire n_2488;
wire n_1980;
wire n_5464;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_6026;
wire n_6070;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_5589;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1614;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_5475;
wire n_5807;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_688;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_4386;
wire n_2995;
wire n_5273;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_5439;
wire n_4955;
wire n_4149;
wire n_5936;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_856;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_6069;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_5706;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_5431;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_6153;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_5627;
wire n_5774;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_5798;
wire n_2984;
wire n_5187;
wire n_5875;
wire n_4024;
wire n_1508;
wire n_5621;
wire n_5608;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_5844;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_6164;
wire n_768;
wire n_6173;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_2598;
wire n_1916;
wire n_1683;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_5867;
wire n_750;
wire n_5508;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_6158;
wire n_5597;
wire n_4915;
wire n_4328;
wire n_6090;
wire n_1057;
wire n_2785;
wire n_5515;
wire n_1997;
wire n_5662;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_5862;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_5697;
wire n_3416;
wire n_3498;
wire n_5767;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_5462;
wire n_1497;
wire n_5980;
wire n_3672;
wire n_5318;
wire n_3533;
wire n_1622;
wire n_6105;
wire n_4725;
wire n_6022;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5987;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_5988;
wire n_5585;
wire n_6058;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_5348;
wire n_1332;
wire n_5480;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_936;
wire n_3821;
wire n_3045;
wire n_885;
wire n_6161;
wire n_2970;
wire n_2167;
wire n_2342;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_5904;
wire n_4739;
wire n_6062;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_5461;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_5503;
wire n_5845;
wire n_5945;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_5600;
wire n_5755;
wire n_707;
wire n_1900;
wire n_5048;
wire n_6053;
wire n_3246;
wire n_3381;
wire n_1548;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_6123;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_5448;
wire n_2939;
wire n_5749;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_3517;
wire n_4045;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_5993;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_6020;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_6162;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_1650;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_5418;
wire n_6178;
wire n_4088;
wire n_3398;
wire n_5685;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_5459;
wire n_1019;
wire n_4170;
wire n_4143;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_5839;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_6175;
wire n_3806;
wire n_5514;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_5351;
wire n_5909;
wire n_671;
wire n_6093;
wire n_4543;
wire n_740;
wire n_703;
wire n_4157;
wire n_4229;
wire n_5293;
wire n_6099;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_5400;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_6140;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_5890;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_676;
wire n_832;
wire n_3049;
wire n_5389;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_5891;
wire n_3541;
wire n_6101;
wire n_3117;
wire n_5935;
wire n_4930;
wire n_5623;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_5693;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_5663;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_5990;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_5647;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_5203;
wire n_930;
wire n_2620;
wire n_5162;
wire n_6134;
wire n_1945;
wire n_5426;
wire n_1656;
wire n_5803;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_653;
wire n_1414;
wire n_5285;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_5365;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_5715;
wire n_4920;
wire n_870;
wire n_5395;
wire n_1253;
wire n_5709;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_5634;
wire n_5672;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_5799;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_5617;
wire n_1829;
wire n_5266;
wire n_5580;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_5390;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_5593;
wire n_4769;
wire n_5764;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_5385;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_6177;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_5853;
wire n_5982;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_5917;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5376;
wire n_5106;
wire n_6116;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_5561;
wire n_5410;
wire n_2215;
wire n_6167;
wire n_1884;
wire n_6170;
wire n_665;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_6094;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_6155;
wire n_1833;
wire n_3903;
wire n_5998;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_5378;
wire n_6028;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_5916;
wire n_681;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_5691;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_5615;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_5468;
wire n_4730;
wire n_5399;
wire n_1234;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_700;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_6077;
wire n_1003;
wire n_5713;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_5550;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_5573;
wire n_1553;
wire n_5939;
wire n_5509;
wire n_5382;
wire n_5659;
wire n_3619;
wire n_1415;
wire n_5881;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_5863;
wire n_2645;
wire n_3904;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_5466;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_5955;
wire n_658;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_6076;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_693;
wire n_1056;
wire n_758;
wire n_5851;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_5796;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_6096;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_5492;
wire n_5995;
wire n_2378;
wire n_887;
wire n_5905;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_5829;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_5734;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_5770;
wire n_1333;
wire n_2496;
wire n_5705;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_5525;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_6052;
wire n_2907;
wire n_5374;
wire n_5575;
wire n_1843;
wire n_5675;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_5297;
wire n_1123;
wire n_1309;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_5959;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_5642;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_6109;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_689;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_5302;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_692;
wire n_5639;
wire n_5781;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_5543;
wire n_1251;
wire n_5361;
wire n_2711;
wire n_4199;
wire n_5885;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_1312;
wire n_5668;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_5463;
wire n_3022;
wire n_5489;
wire n_1165;
wire n_5892;
wire n_4773;
wire n_5654;
wire n_2008;
wire n_6009;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5923;
wire n_5113;
wire n_5479;
wire n_3549;
wire n_5714;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_5510;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_690;
wire n_850;
wire n_5692;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_5555;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_825;
wire n_6066;
wire n_3785;
wire n_2963;
wire n_5366;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_696;
wire n_4886;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_3289;
wire n_2733;
wire n_4055;
wire n_2178;
wire n_5968;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_3519;
wire n_2082;
wire n_678;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_5415;
wire n_5419;
wire n_3805;
wire n_1990;
wire n_2943;
wire n_5205;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_6130;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_5976;
wire n_3128;
wire n_1527;
wire n_5732;
wire n_5372;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_5690;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_5801;
wire n_6047;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5347;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_6021;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_5656;
wire n_1469;
wire n_5125;
wire n_5857;
wire n_2650;
wire n_5652;
wire n_987;
wire n_5499;
wire n_720;
wire n_3348;
wire n_3229;
wire n_1707;
wire n_656;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_684;
wire n_5507;
wire n_1809;
wire n_5569;
wire n_4280;
wire n_1181;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_5455;
wire n_5442;
wire n_5948;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_5511;
wire n_2898;
wire n_5295;
wire n_2368;
wire n_4175;
wire n_5490;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_5836;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_5834;
wire n_3191;
wire n_5584;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_5707;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_5497;
wire n_880;
wire n_3505;
wire n_3540;
wire n_3577;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_1363;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_5481;
wire n_3590;
wire n_2435;
wire n_5344;
wire n_954;
wire n_4419;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_5794;
wire n_1382;
wire n_5408;
wire n_1736;
wire n_4053;
wire n_3848;
wire n_1483;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_5271;
wire n_5964;
wire n_6004;
wire n_2323;
wire n_2784;
wire n_5494;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_3755;
wire n_4042;
wire n_1125;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_5467;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5827;
wire n_5199;
wire n_3407;
wire n_5992;
wire n_5313;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_5513;
wire n_5614;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_3243;
wire n_2462;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_5835;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_5846;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_5592;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_5278;
wire n_3525;
wire n_3314;
wire n_2100;
wire n_5157;
wire n_2993;
wire n_4754;
wire n_3016;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_5708;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_5474;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_5649;
wire n_1905;
wire n_3466;
wire n_762;
wire n_5704;
wire n_4983;
wire n_1778;
wire n_5956;
wire n_5287;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_6007;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_6144;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_5516;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_5698;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_5771;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_5538;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_3141;
wire n_2755;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_5428;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_5677;
wire n_4124;
wire n_5570;
wire n_785;
wire n_5153;
wire n_4611;
wire n_5927;
wire n_5435;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_5566;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_5487;
wire n_5486;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_5889;
wire n_3217;
wire n_1983;
wire n_5391;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_5849;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_6092;
wire n_5951;
wire n_1692;
wire n_1084;
wire n_5912;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_5574;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_6165;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_5469;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_5910;
wire n_5895;
wire n_1041;
wire n_5804;
wire n_3134;
wire n_5965;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_5682;
wire n_5387;
wire n_654;
wire n_5557;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_5681;
wire n_6119;
wire n_1271;
wire n_4901;
wire n_4145;
wire n_4821;
wire n_1545;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_2141;
wire n_5316;
wire n_5703;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_5564;
wire n_5620;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_5406;
wire n_2125;
wire n_2561;
wire n_652;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_5724;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_5806;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_5738;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_5710;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_5979;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_6044;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_5517;
wire n_3207;
wire n_5605;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_6125;
wire n_655;
wire n_4726;
wire n_1045;
wire n_5907;
wire n_786;
wire n_1559;
wire n_6045;
wire n_1872;
wire n_5040;
wire n_6063;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_1727;
wire n_6154;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_5977;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_6003;
wire n_3843;
wire n_1098;
wire n_5746;
wire n_2045;
wire n_817;
wire n_5451;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_3543;
wire n_3621;
wire n_6031;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_6060;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_5417;
wire n_2587;
wire n_3199;
wire n_680;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_5864;
wire n_1953;
wire n_4741;
wire n_6172;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_5432;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_5453;
wire n_3658;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_5842;
wire n_5814;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_5699;
wire n_5531;
wire n_5765;
wire n_2953;
wire n_4295;
wire n_5943;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_6088;
wire n_5777;
wire n_4225;
wire n_747;
wire n_2565;
wire n_5495;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5655;
wire n_5064;
wire n_5610;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_5759;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_6035;
wire n_957;
wire n_1994;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_6114;
wire n_4568;
wire n_1205;
wire n_6061;
wire n_5559;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_5786;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_5737;
wire n_3604;
wire n_1501;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_5768;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_3811;
wire n_2022;
wire n_910;
wire n_1721;
wire n_3494;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_5350;
wire n_5470;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_5872;
wire n_5858;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_5700;
wire n_1500;
wire n_6037;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_5874;
wire n_904;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_5873;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_5588;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_5736;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_5928;
wire n_4089;
wire n_5478;
wire n_6016;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_6176;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_6080;
wire n_4865;
wire n_1039;
wire n_6078;
wire n_2043;
wire n_1480;
wire n_6056;
wire n_5832;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_5812;
wire n_2540;
wire n_973;
wire n_5743;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_679;
wire n_1629;
wire n_5368;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_5971;
wire n_812;
wire n_6145;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_5933;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_670;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_6030;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_5996;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_5903;
wire n_5986;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_5782;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_6050;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_5563;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_5840;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_2647;
wire n_883;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_5717;
wire n_6017;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_5720;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_5871;
wire n_1285;
wire n_1985;
wire n_5898;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_5896;
wire n_1649;
wire n_4555;
wire n_5882;
wire n_5940;
wire n_6089;
wire n_5650;
wire n_4969;
wire n_6057;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_5567;
wire n_1344;
wire n_6174;
wire n_2730;
wire n_2495;
wire n_6087;
wire n_5249;
wire n_2603;
wire n_2090;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_5625;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_5969;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_5022;
wire n_5670;
wire n_1280;
wire n_6041;
wire n_3296;
wire n_5276;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_5879;
wire n_4403;
wire n_5238;
wire n_6166;
wire n_5855;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_6081;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_5429;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_5535;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_6002;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_821;
wire n_4372;
wire n_1068;
wire n_982;
wire n_5640;
wire n_2831;
wire n_932;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_5560;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_5544;
wire n_6108;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_5744;
wire n_4013;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_5841;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_6086;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_5941;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_5611;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_3734;
wire n_1014;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_5701;
wire n_3746;
wire n_6067;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_4478;
wire n_1662;
wire n_2818;
wire n_1359;
wire n_5367;
wire n_3794;
wire n_674;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5970;
wire n_5202;
wire n_702;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_6111;
wire n_3058;
wire n_3861;
wire n_675;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_6011;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_5502;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_5850;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_5876;
wire n_5521;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_697;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_5856;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_5837;
wire n_4675;
wire n_2663;
wire n_5825;
wire n_4018;
wire n_5491;
wire n_2987;
wire n_694;
wire n_2938;
wire n_3780;
wire n_5496;
wire n_5802;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_5547;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_5596;
wire n_6074;
wire n_2684;
wire n_5983;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_5604;
wire n_1756;
wire n_1128;
wire n_5411;
wire n_673;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_5815;
wire n_4191;
wire n_5695;
wire n_6027;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_6095;
wire n_5331;
wire n_4330;
wire n_5311;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_5797;
wire n_4240;
wire n_3491;
wire n_5572;
wire n_1488;
wire n_704;
wire n_2148;
wire n_4162;
wire n_5565;
wire n_2339;
wire n_2861;
wire n_5520;
wire n_2731;
wire n_1999;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_5800;
wire n_5984;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_5888;
wire n_5669;
wire n_5772;
wire n_2208;
wire n_4775;
wire n_5884;
wire n_4864;
wire n_5758;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_5603;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_5763;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_6128;
wire n_2489;
wire n_6029;
wire n_1087;
wire n_657;
wire n_5751;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_5924;
wire n_1505;
wire n_5712;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_4871;
wire n_2403;
wire n_1070;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_6005;
wire n_4453;
wire n_3559;
wire n_5449;
wire n_4005;
wire n_6169;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_2424;
wire n_745;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_5926;
wire n_716;
wire n_1475;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_5398;
wire n_5860;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_6106;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_5919;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_6098;
wire n_6014;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_5043;
wire n_1755;
wire n_2025;
wire n_2357;
wire n_5583;
wire n_4654;
wire n_3640;
wire n_1159;
wire n_3481;
wire n_995;
wire n_2250;
wire n_3033;
wire n_6142;
wire n_5775;
wire n_2374;
wire n_1681;
wire n_6034;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_6071;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_6143;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_5483;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_5785;
wire n_2343;
wire n_793;
wire n_5967;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_5780;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_6084;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_5966;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_994;
wire n_5735;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_5752;
wire n_1661;
wire n_5360;
wire n_6104;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_6082;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_667;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_5877;
wire n_6018;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_5869;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_5632;
wire n_5582;
wire n_5425;
wire n_5886;
wire n_1216;
wire n_2716;
wire n_6032;
wire n_2452;
wire n_3650;
wire n_5446;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_5678;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_6122;
wire n_2790;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_3784;
wire n_5437;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_5454;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_5407;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_5913;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_5944;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_6000;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_5974;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_6046;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_6118;
wire n_5810;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_5991;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_5702;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_5914;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_5590;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_5809;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_5349;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_6146;
wire n_5813;
wire n_790;
wire n_5833;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_5616;
wire n_5805;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_5816;
wire n_3156;
wire n_672;
wire n_1941;
wire n_3483;
wire n_5416;
wire n_706;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_6102;
wire n_3097;
wire n_660;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_6072;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_5167;
wire n_5661;
wire n_5830;
wire n_5932;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_1476;
wire n_841;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_5558;
wire n_1826;
wire n_5687;
wire n_5383;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5587;
wire n_5236;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_661;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5954;
wire n_6156;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_5651;
wire n_4630;
wire n_1217;
wire n_5645;
wire n_3990;
wire n_1628;
wire n_5766;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_5878;
wire n_5671;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_5412;
wire n_2380;
wire n_769;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_669;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_5733;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_5791;
wire n_5727;
wire n_761;
wire n_5946;
wire n_5997;
wire n_2492;
wire n_3778;
wire n_5328;
wire n_5657;
wire n_1173;
wire n_4974;
wire n_5975;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_5938;
wire n_5602;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_5579;
wire n_1922;
wire n_5750;
wire n_4823;
wire n_5831;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_4243;
wire n_2205;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_5666;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_4142;
wire n_3671;
wire n_2015;
wire n_3982;
wire n_6103;
wire n_2609;
wire n_1161;
wire n_5546;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_5994;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_5626;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_5633;
wire n_1218;
wire n_5664;
wire n_5921;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_6159;
wire n_2429;
wire n_985;
wire n_2440;
wire n_6054;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_6152;
wire n_4075;
wire n_5340;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_5280;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_5925;
wire n_2909;
wire n_754;
wire n_6138;
wire n_5369;
wire n_975;
wire n_5730;
wire n_5576;
wire n_3359;
wire n_5272;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_5646;
wire n_5624;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_730;
wire n_5817;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_5586;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_6038;
wire n_5861;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_5619;
wire n_6112;
wire n_3965;
wire n_5859;
wire n_5380;
wire n_4500;
wire n_5065;
wire n_862;
wire n_5776;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_5606;
wire n_5644;
wire n_2813;
wire n_1935;
wire n_5826;
wire n_2027;
wire n_2091;
wire n_5920;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_6180;
wire n_5683;
wire n_2677;
wire n_3182;
wire n_5756;
wire n_3283;
wire n_5527;
wire n_1742;
wire n_4030;

INVx1_ASAP7_75t_L g652 ( 
.A(n_292),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_160),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_282),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_222),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_382),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_464),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_328),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_248),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_217),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_422),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_320),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_553),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_642),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_212),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_99),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_55),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_136),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_467),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_103),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_608),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_598),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_250),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_552),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_195),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_584),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_414),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_78),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_249),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_576),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_385),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_249),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_578),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_53),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_528),
.Y(n_685)
);

CKINVDCx16_ASAP7_75t_R g686 ( 
.A(n_310),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_56),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_650),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_502),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_516),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_193),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_56),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_2),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_644),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_533),
.Y(n_695)
);

BUFx10_ASAP7_75t_L g696 ( 
.A(n_500),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_137),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_635),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_340),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_211),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_77),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_460),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_4),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_176),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_3),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_461),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_328),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_634),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_398),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_66),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_419),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_314),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_514),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_285),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_433),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_10),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_140),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_135),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_270),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_395),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_349),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_178),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_393),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_451),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_109),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_223),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_323),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_476),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_67),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_217),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_434),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_413),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_18),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_105),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_214),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_93),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_625),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_243),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_624),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_129),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_513),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_500),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_497),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_534),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_254),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_613),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_305),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_589),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_379),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_469),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_195),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_48),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_533),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_265),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_504),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_625),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_172),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_516),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_1),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_99),
.Y(n_760)
);

CKINVDCx16_ASAP7_75t_R g761 ( 
.A(n_103),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_407),
.Y(n_762)
);

INVxp33_ASAP7_75t_SL g763 ( 
.A(n_419),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_16),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_622),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_63),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_171),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_77),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_544),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_288),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_101),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_612),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_153),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_479),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_550),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_168),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_642),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_568),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_14),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_505),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_492),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_132),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_214),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_385),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_600),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_595),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_648),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_471),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_263),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_605),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_221),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_22),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_228),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_581),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_339),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_279),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_614),
.Y(n_797)
);

CKINVDCx16_ASAP7_75t_R g798 ( 
.A(n_517),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_312),
.Y(n_799)
);

INVx1_ASAP7_75t_SL g800 ( 
.A(n_609),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_590),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_192),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_486),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_323),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_601),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_52),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_535),
.Y(n_807)
);

CKINVDCx16_ASAP7_75t_R g808 ( 
.A(n_596),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_544),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_396),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_371),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_109),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_114),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_503),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_213),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_458),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_355),
.Y(n_817)
);

BUFx8_ASAP7_75t_SL g818 ( 
.A(n_436),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_372),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_289),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_317),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_588),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_72),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_327),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_288),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_144),
.Y(n_826)
);

CKINVDCx16_ASAP7_75t_R g827 ( 
.A(n_180),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_276),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_639),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_202),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_122),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_227),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_514),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_483),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_286),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_626),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_526),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_517),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_307),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_519),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_496),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_320),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_352),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_149),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_488),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_162),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_96),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_291),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_62),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_293),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_315),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_643),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_100),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_593),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_189),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_151),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_510),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_477),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_133),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_540),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_295),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_422),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_253),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_312),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_572),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_10),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_243),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_325),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_185),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_480),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_527),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_55),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_156),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_98),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_61),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_105),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_373),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_178),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_403),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_508),
.Y(n_880)
);

CKINVDCx16_ASAP7_75t_R g881 ( 
.A(n_383),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_381),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_493),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_78),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_31),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_615),
.Y(n_886)
);

BUFx10_ASAP7_75t_L g887 ( 
.A(n_259),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_280),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_621),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_16),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_128),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_276),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_135),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_578),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_114),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_534),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_545),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_201),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_187),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_482),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_405),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_30),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_449),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_627),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_336),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_258),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_466),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_602),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_2),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_459),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_357),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_31),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_224),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_645),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_237),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_449),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_205),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_194),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_628),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_610),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_368),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_535),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_83),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_506),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_85),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_512),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_645),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_30),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_363),
.Y(n_929)
);

BUFx5_ASAP7_75t_L g930 ( 
.A(n_82),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_395),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_247),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_429),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_159),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_162),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_613),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_632),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_266),
.Y(n_938)
);

BUFx5_ASAP7_75t_L g939 ( 
.A(n_110),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_6),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_11),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_441),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_67),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_280),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_3),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_158),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_334),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_608),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_79),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_141),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_204),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_364),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_569),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_573),
.Y(n_954)
);

BUFx10_ASAP7_75t_L g955 ( 
.A(n_377),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_370),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_400),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_403),
.Y(n_958)
);

CKINVDCx16_ASAP7_75t_R g959 ( 
.A(n_125),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_355),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_397),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_405),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_6),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_46),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_571),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_397),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_181),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_529),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_111),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_70),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_628),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_191),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_345),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_155),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_111),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_618),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_432),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_45),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_284),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_120),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_54),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_336),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_481),
.Y(n_983)
);

CKINVDCx16_ASAP7_75t_R g984 ( 
.A(n_425),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_340),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_475),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_42),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_329),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_69),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_539),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_68),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_39),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_246),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_57),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_614),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_96),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_40),
.Y(n_997)
);

BUFx5_ASAP7_75t_L g998 ( 
.A(n_485),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_215),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_574),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_478),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_651),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_327),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_453),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_261),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_151),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_412),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_637),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_330),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_191),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_193),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_400),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_361),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_651),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_647),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_163),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_371),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_240),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_225),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_523),
.Y(n_1020)
);

BUFx10_ASAP7_75t_L g1021 ( 
.A(n_26),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_250),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_427),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_329),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_583),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_82),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_66),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_8),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_456),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_542),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_636),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_175),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_484),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_278),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_21),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_166),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_221),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_281),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_546),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_524),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_393),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_424),
.Y(n_1042)
);

BUFx8_ASAP7_75t_SL g1043 ( 
.A(n_199),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_24),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_284),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_89),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_379),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_599),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_545),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_157),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_277),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_406),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_251),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_386),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_93),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_369),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_154),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_41),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_515),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_121),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_442),
.Y(n_1061)
);

BUFx5_ASAP7_75t_L g1062 ( 
.A(n_637),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_331),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_555),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_81),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_238),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_554),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_21),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_48),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_520),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_251),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_313),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_587),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_603),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_165),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_498),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_58),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_456),
.Y(n_1078)
);

BUFx5_ASAP7_75t_L g1079 ( 
.A(n_181),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_287),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_321),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_76),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_231),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_570),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_623),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_52),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_252),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_473),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_431),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_201),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_620),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_593),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_468),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_156),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_509),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_53),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_261),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_307),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_560),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_530),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_347),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_52),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_170),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_501),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_283),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_478),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_599),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_184),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_406),
.Y(n_1110)
);

INVx4_ASAP7_75t_R g1111 ( 
.A(n_399),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_33),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_509),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_62),
.Y(n_1114)
);

BUFx10_ASAP7_75t_L g1115 ( 
.A(n_164),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_290),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_586),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_360),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_15),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_227),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_7),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_84),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_300),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_390),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_115),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_363),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_352),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_218),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_125),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_479),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_604),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_31),
.Y(n_1132)
);

INVxp67_ASAP7_75t_L g1133 ( 
.A(n_357),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_409),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_91),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_390),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_523),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_278),
.Y(n_1138)
);

CKINVDCx16_ASAP7_75t_R g1139 ( 
.A(n_686),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_818),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_818),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1128),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1043),
.Y(n_1143)
);

CKINVDCx14_ASAP7_75t_R g1144 ( 
.A(n_684),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_930),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_930),
.Y(n_1146)
);

INVxp33_ASAP7_75t_SL g1147 ( 
.A(n_1137),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1043),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_684),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_930),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_930),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_930),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_930),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_930),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_675),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_930),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_930),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_930),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_939),
.Y(n_1159)
);

INVxp33_ASAP7_75t_SL g1160 ( 
.A(n_1137),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_686),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_761),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_939),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_939),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_902),
.Y(n_1165)
);

NOR2xp67_ASAP7_75t_L g1166 ( 
.A(n_690),
.B(n_0),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_939),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_755),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_761),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_939),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_902),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_939),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_939),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_832),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_939),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_939),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_939),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_798),
.Y(n_1178)
);

BUFx10_ASAP7_75t_L g1179 ( 
.A(n_779),
.Y(n_1179)
);

INVxp33_ASAP7_75t_SL g1180 ( 
.A(n_690),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_998),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_798),
.Y(n_1182)
);

INVxp67_ASAP7_75t_L g1183 ( 
.A(n_987),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_998),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_998),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_998),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_998),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_998),
.Y(n_1188)
);

CKINVDCx16_ASAP7_75t_R g1189 ( 
.A(n_808),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_998),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_998),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_998),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_998),
.Y(n_1193)
);

INVxp33_ASAP7_75t_SL g1194 ( 
.A(n_743),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1062),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1062),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1062),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1062),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_763),
.B(n_0),
.Y(n_1199)
);

INVxp67_ASAP7_75t_L g1200 ( 
.A(n_987),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1062),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1062),
.Y(n_1202)
);

INVx4_ASAP7_75t_R g1203 ( 
.A(n_928),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_808),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_827),
.Y(n_1205)
);

CKINVDCx16_ASAP7_75t_R g1206 ( 
.A(n_827),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1062),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1062),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1062),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1062),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1079),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1079),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1079),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_881),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1079),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1079),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_779),
.Y(n_1217)
);

INVxp67_ASAP7_75t_SL g1218 ( 
.A(n_779),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1079),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1079),
.Y(n_1220)
);

CKINVDCx20_ASAP7_75t_R g1221 ( 
.A(n_833),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1079),
.Y(n_1222)
);

CKINVDCx16_ASAP7_75t_R g1223 ( 
.A(n_881),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1079),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1079),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_744),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_1087),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_744),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_744),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_744),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_744),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_1106),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_744),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_744),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_779),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_886),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_R g1237 ( 
.A(n_1131),
.B(n_0),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_959),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_886),
.Y(n_1239)
);

INVxp67_ASAP7_75t_SL g1240 ( 
.A(n_779),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_886),
.Y(n_1241)
);

CKINVDCx16_ASAP7_75t_R g1242 ( 
.A(n_959),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_984),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_984),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_656),
.Y(n_1245)
);

INVxp33_ASAP7_75t_SL g1246 ( 
.A(n_743),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_886),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_779),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_779),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_992),
.Y(n_1250)
);

CKINVDCx16_ASAP7_75t_R g1251 ( 
.A(n_705),
.Y(n_1251)
);

INVxp67_ASAP7_75t_SL g1252 ( 
.A(n_992),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_886),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_992),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1087),
.Y(n_1255)
);

INVxp67_ASAP7_75t_SL g1256 ( 
.A(n_992),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_880),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_992),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_886),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_886),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_656),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_919),
.Y(n_1262)
);

CKINVDCx16_ASAP7_75t_R g1263 ( 
.A(n_705),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_919),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_919),
.Y(n_1265)
);

INVxp33_ASAP7_75t_SL g1266 ( 
.A(n_880),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_992),
.Y(n_1267)
);

INVxp67_ASAP7_75t_SL g1268 ( 
.A(n_992),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_653),
.Y(n_1269)
);

INVxp67_ASAP7_75t_SL g1270 ( 
.A(n_928),
.Y(n_1270)
);

INVxp67_ASAP7_75t_SL g1271 ( 
.A(n_928),
.Y(n_1271)
);

INVxp33_ASAP7_75t_SL g1272 ( 
.A(n_933),
.Y(n_1272)
);

INVxp67_ASAP7_75t_SL g1273 ( 
.A(n_919),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_707),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_933),
.Y(n_1275)
);

BUFx2_ASAP7_75t_SL g1276 ( 
.A(n_768),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_654),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_655),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_707),
.Y(n_1279)
);

CKINVDCx16_ASAP7_75t_R g1280 ( 
.A(n_705),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_919),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_919),
.Y(n_1282)
);

INVxp33_ASAP7_75t_L g1283 ( 
.A(n_787),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_787),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_736),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_919),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_929),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_929),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_929),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_929),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_929),
.B(n_1),
.Y(n_1291)
);

INVxp33_ASAP7_75t_L g1292 ( 
.A(n_852),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_964),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_964),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_964),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_736),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_718),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_978),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_978),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_978),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1097),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_929),
.Y(n_1302)
);

INVxp33_ASAP7_75t_SL g1303 ( 
.A(n_716),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1097),
.Y(n_1304)
);

INVxp33_ASAP7_75t_SL g1305 ( 
.A(n_733),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1097),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_718),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_718),
.Y(n_1308)
);

INVxp33_ASAP7_75t_L g1309 ( 
.A(n_852),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_734),
.Y(n_1310)
);

CKINVDCx14_ASAP7_75t_R g1311 ( 
.A(n_705),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_929),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_936),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_734),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_936),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_734),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_815),
.Y(n_1317)
);

CKINVDCx14_ASAP7_75t_R g1318 ( 
.A(n_1021),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_936),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_815),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_815),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_942),
.Y(n_1322)
);

INVxp33_ASAP7_75t_SL g1323 ( 
.A(n_759),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_942),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_942),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1004),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_956),
.Y(n_1327)
);

INVxp33_ASAP7_75t_SL g1328 ( 
.A(n_764),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_657),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_956),
.Y(n_1330)
);

INVxp33_ASAP7_75t_L g1331 ( 
.A(n_1004),
.Y(n_1331)
);

CKINVDCx14_ASAP7_75t_R g1332 ( 
.A(n_1021),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_658),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_956),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1084),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1029),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_760),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1029),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1029),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1067),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1084),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1067),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_936),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1067),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1100),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1076),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1076),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_936),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1076),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_936),
.Y(n_1350)
);

CKINVDCx16_ASAP7_75t_R g1351 ( 
.A(n_1021),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_760),
.Y(n_1352)
);

NOR2xp67_ASAP7_75t_L g1353 ( 
.A(n_669),
.B(n_2),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1138),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1138),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1138),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_659),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_991),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_693),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_772),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_991),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_693),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_703),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_991),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_752),
.Y(n_1365)
);

CKINVDCx16_ASAP7_75t_R g1366 ( 
.A(n_1021),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_752),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_885),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_885),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_772),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_991),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_912),
.Y(n_1372)
);

CKINVDCx16_ASAP7_75t_R g1373 ( 
.A(n_696),
.Y(n_1373)
);

BUFx8_ASAP7_75t_SL g1374 ( 
.A(n_1109),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_660),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_941),
.Y(n_1376)
);

INVxp33_ASAP7_75t_SL g1377 ( 
.A(n_792),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_945),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_991),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_945),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_963),
.Y(n_1381)
);

INVxp33_ASAP7_75t_SL g1382 ( 
.A(n_806),
.Y(n_1382)
);

INVxp67_ASAP7_75t_SL g1383 ( 
.A(n_991),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_991),
.Y(n_1384)
);

CKINVDCx16_ASAP7_75t_R g1385 ( 
.A(n_696),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_661),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1031),
.Y(n_1387)
);

CKINVDCx14_ASAP7_75t_R g1388 ( 
.A(n_1109),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_963),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1031),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1035),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1031),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1035),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1080),
.B(n_3),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1080),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1031),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1031),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1031),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1031),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1055),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1055),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_774),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1129),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1055),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1055),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1055),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1055),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1055),
.Y(n_1408)
);

CKINVDCx16_ASAP7_75t_R g1409 ( 
.A(n_696),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1085),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_1085),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_774),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1129),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1085),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1085),
.Y(n_1415)
);

INVxp67_ASAP7_75t_SL g1416 ( 
.A(n_1085),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1085),
.Y(n_1417)
);

INVxp67_ASAP7_75t_SL g1418 ( 
.A(n_1085),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1128),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1128),
.Y(n_1420)
);

INVxp33_ASAP7_75t_SL g1421 ( 
.A(n_866),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1128),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1128),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_664),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1128),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_652),
.Y(n_1426)
);

CKINVDCx14_ASAP7_75t_R g1427 ( 
.A(n_696),
.Y(n_1427)
);

CKINVDCx14_ASAP7_75t_R g1428 ( 
.A(n_887),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_665),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_887),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_662),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_890),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_666),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_666),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_668),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_672),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_674),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_674),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1069),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_676),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_676),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_681),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_887),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_887),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_681),
.Y(n_1445)
);

INVxp67_ASAP7_75t_SL g1446 ( 
.A(n_663),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_663),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_688),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_955),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_688),
.Y(n_1450)
);

INVxp67_ASAP7_75t_SL g1451 ( 
.A(n_663),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_691),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_691),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_692),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_670),
.Y(n_1455)
);

CKINVDCx16_ASAP7_75t_R g1456 ( 
.A(n_955),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_692),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_671),
.Y(n_1458)
);

CKINVDCx16_ASAP7_75t_R g1459 ( 
.A(n_955),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_702),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_702),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_704),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_683),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_704),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_708),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_776),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_708),
.Y(n_1467)
);

INVxp67_ASAP7_75t_SL g1468 ( 
.A(n_683),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_711),
.Y(n_1469)
);

INVxp33_ASAP7_75t_SL g1470 ( 
.A(n_909),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_711),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_776),
.Y(n_1472)
);

INVxp33_ASAP7_75t_SL g1473 ( 
.A(n_940),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_673),
.Y(n_1474)
);

CKINVDCx14_ASAP7_75t_R g1475 ( 
.A(n_955),
.Y(n_1475)
);

INVxp67_ASAP7_75t_SL g1476 ( 
.A(n_683),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_712),
.Y(n_1477)
);

INVxp67_ASAP7_75t_SL g1478 ( 
.A(n_709),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_712),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_678),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_715),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_709),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_715),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_679),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_731),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_680),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_731),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_735),
.Y(n_1488)
);

CKINVDCx14_ASAP7_75t_R g1489 ( 
.A(n_1115),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_682),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_735),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_844),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_685),
.Y(n_1493)
);

INVxp33_ASAP7_75t_SL g1494 ( 
.A(n_981),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_844),
.Y(n_1495)
);

INVxp33_ASAP7_75t_L g1496 ( 
.A(n_740),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1069),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_740),
.Y(n_1498)
);

INVxp33_ASAP7_75t_L g1499 ( 
.A(n_741),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_687),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_741),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_709),
.Y(n_1502)
);

INVxp33_ASAP7_75t_SL g1503 ( 
.A(n_997),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_762),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_762),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_762),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_689),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_748),
.Y(n_1508)
);

CKINVDCx16_ASAP7_75t_R g1509 ( 
.A(n_1115),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_765),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1115),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_765),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_765),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_778),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_748),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_778),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_778),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_790),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_790),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_790),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_796),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_796),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_796),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_921),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_1132),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_921),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_921),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_922),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_922),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_750),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_922),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_924),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_924),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1115),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_924),
.Y(n_1535)
);

INVxp33_ASAP7_75t_SL g1536 ( 
.A(n_1028),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_948),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_694),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_948),
.Y(n_1539)
);

CKINVDCx16_ASAP7_75t_R g1540 ( 
.A(n_850),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_948),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_962),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_962),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_962),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_985),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_985),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_985),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1010),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1010),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1010),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1050),
.Y(n_1551)
);

INVxp67_ASAP7_75t_SL g1552 ( 
.A(n_1050),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1050),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1051),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1051),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_695),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1051),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1057),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1057),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_697),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1057),
.Y(n_1561)
);

INVxp67_ASAP7_75t_SL g1562 ( 
.A(n_1063),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1140),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1226),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1161),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1226),
.Y(n_1566)
);

CKINVDCx6p67_ASAP7_75t_R g1567 ( 
.A(n_1139),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1228),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1270),
.B(n_768),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1217),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1156),
.A2(n_1077),
.B(n_1063),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1217),
.Y(n_1572)
);

INVx5_ASAP7_75t_L g1573 ( 
.A(n_1217),
.Y(n_1573)
);

OAI22x1_ASAP7_75t_SL g1574 ( 
.A1(n_1245),
.A2(n_850),
.B1(n_855),
.B2(n_853),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1217),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1218),
.B(n_1063),
.Y(n_1576)
);

INVx5_ASAP7_75t_L g1577 ( 
.A(n_1217),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1250),
.Y(n_1578)
);

BUFx12f_ASAP7_75t_L g1579 ( 
.A(n_1140),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1147),
.A2(n_1058),
.B1(n_1068),
.B2(n_1044),
.Y(n_1580)
);

BUFx12f_ASAP7_75t_L g1581 ( 
.A(n_1141),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1250),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1161),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1155),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1228),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_1250),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1235),
.Y(n_1587)
);

INVx4_ASAP7_75t_L g1588 ( 
.A(n_1302),
.Y(n_1588)
);

BUFx8_ASAP7_75t_SL g1589 ( 
.A(n_1374),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1240),
.B(n_1077),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1252),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1256),
.B(n_1077),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1268),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1250),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1250),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1162),
.Y(n_1596)
);

INVx5_ASAP7_75t_L g1597 ( 
.A(n_1258),
.Y(n_1597)
);

BUFx8_ASAP7_75t_L g1598 ( 
.A(n_1165),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1258),
.Y(n_1599)
);

BUFx12f_ASAP7_75t_L g1600 ( 
.A(n_1141),
.Y(n_1600)
);

BUFx12f_ASAP7_75t_L g1601 ( 
.A(n_1143),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1297),
.Y(n_1602)
);

NOR2x1_ASAP7_75t_L g1603 ( 
.A(n_1398),
.B(n_757),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1271),
.B(n_1123),
.Y(n_1604)
);

OA21x2_ASAP7_75t_L g1605 ( 
.A1(n_1229),
.A2(n_1130),
.B(n_1124),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1258),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1261),
.Y(n_1607)
);

BUFx12f_ASAP7_75t_L g1608 ( 
.A(n_1143),
.Y(n_1608)
);

BUFx8_ASAP7_75t_SL g1609 ( 
.A(n_1274),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1430),
.Y(n_1610)
);

BUFx12f_ASAP7_75t_L g1611 ( 
.A(n_1148),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_SL g1612 ( 
.A1(n_1244),
.A2(n_855),
.B1(n_862),
.B2(n_853),
.Y(n_1612)
);

CKINVDCx16_ASAP7_75t_R g1613 ( 
.A(n_1189),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1258),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1235),
.Y(n_1615)
);

INVx5_ASAP7_75t_L g1616 ( 
.A(n_1258),
.Y(n_1616)
);

BUFx8_ASAP7_75t_L g1617 ( 
.A(n_1165),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1229),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1302),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1273),
.B(n_768),
.Y(n_1620)
);

BUFx8_ASAP7_75t_SL g1621 ( 
.A(n_1279),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1302),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1230),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1302),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1342),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_1302),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1142),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1430),
.Y(n_1628)
);

INVx5_ASAP7_75t_L g1629 ( 
.A(n_1312),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1147),
.A2(n_1119),
.B1(n_1121),
.B2(n_1112),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1248),
.Y(n_1631)
);

BUFx8_ASAP7_75t_SL g1632 ( 
.A(n_1285),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1251),
.B(n_789),
.Y(n_1633)
);

INVx4_ASAP7_75t_L g1634 ( 
.A(n_1312),
.Y(n_1634)
);

INVx5_ASAP7_75t_L g1635 ( 
.A(n_1312),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1160),
.A2(n_699),
.B1(n_700),
.B2(n_698),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1312),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1162),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1446),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_L g1640 ( 
.A(n_1312),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1142),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1148),
.Y(n_1642)
);

BUFx6f_ASAP7_75t_L g1643 ( 
.A(n_1319),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1248),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1160),
.A2(n_706),
.B1(n_710),
.B2(n_701),
.Y(n_1645)
);

CKINVDCx6p67_ASAP7_75t_R g1646 ( 
.A(n_1206),
.Y(n_1646)
);

XOR2xp5_ASAP7_75t_L g1647 ( 
.A(n_1296),
.B(n_937),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1169),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1379),
.B(n_789),
.Y(n_1649)
);

INVx3_ASAP7_75t_L g1650 ( 
.A(n_1142),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1249),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1451),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1383),
.B(n_789),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1443),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1411),
.B(n_793),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1230),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1254),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1443),
.Y(n_1658)
);

BUFx8_ASAP7_75t_SL g1659 ( 
.A(n_1337),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_1319),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1231),
.Y(n_1661)
);

INVx5_ASAP7_75t_L g1662 ( 
.A(n_1319),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1267),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_SL g1664 ( 
.A1(n_1180),
.A2(n_875),
.B1(n_901),
.B2(n_862),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1231),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1233),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1416),
.B(n_793),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1233),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1319),
.Y(n_1669)
);

BUFx6f_ASAP7_75t_L g1670 ( 
.A(n_1319),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1371),
.Y(n_1671)
);

BUFx8_ASAP7_75t_SL g1672 ( 
.A(n_1352),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1178),
.Y(n_1673)
);

INVx4_ASAP7_75t_L g1674 ( 
.A(n_1371),
.Y(n_1674)
);

OA21x2_ASAP7_75t_L g1675 ( 
.A1(n_1234),
.A2(n_1130),
.B(n_1124),
.Y(n_1675)
);

BUFx12f_ASAP7_75t_L g1676 ( 
.A(n_1178),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1234),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1182),
.Y(n_1678)
);

INVx4_ASAP7_75t_L g1679 ( 
.A(n_1371),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1236),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1418),
.B(n_1123),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1276),
.B(n_1123),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1371),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1342),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1387),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1267),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_1360),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1182),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1387),
.Y(n_1689)
);

BUFx12f_ASAP7_75t_L g1690 ( 
.A(n_1204),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1313),
.Y(n_1691)
);

BUFx12f_ASAP7_75t_L g1692 ( 
.A(n_1204),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_SL g1693 ( 
.A(n_1284),
.B(n_910),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1236),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1307),
.B(n_793),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1239),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1387),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1179),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1303),
.B(n_817),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1404),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1404),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1239),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1388),
.A2(n_714),
.B1(n_717),
.B2(n_713),
.Y(n_1703)
);

OAI21x1_ASAP7_75t_L g1704 ( 
.A1(n_1156),
.A2(n_775),
.B(n_770),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1205),
.Y(n_1705)
);

BUFx8_ASAP7_75t_L g1706 ( 
.A(n_1171),
.Y(n_1706)
);

CKINVDCx20_ASAP7_75t_R g1707 ( 
.A(n_1370),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1468),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1179),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1398),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1476),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1313),
.Y(n_1712)
);

OA21x2_ASAP7_75t_L g1713 ( 
.A1(n_1241),
.A2(n_1134),
.B(n_775),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1315),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1179),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1315),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1157),
.A2(n_777),
.B(n_770),
.Y(n_1717)
);

NOR2xp67_ASAP7_75t_L g1718 ( 
.A(n_1269),
.B(n_669),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1241),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_1343),
.Y(n_1720)
);

OAI22x1_ASAP7_75t_SL g1721 ( 
.A1(n_1402),
.A2(n_990),
.B1(n_1015),
.B2(n_937),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1247),
.Y(n_1722)
);

INVx4_ASAP7_75t_L g1723 ( 
.A(n_1157),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1180),
.A2(n_720),
.B1(n_723),
.B2(n_719),
.Y(n_1724)
);

AOI22x1_ASAP7_75t_SL g1725 ( 
.A1(n_1412),
.A2(n_1122),
.B1(n_1015),
.B2(n_1016),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1247),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1348),
.Y(n_1727)
);

OAI21x1_ASAP7_75t_L g1728 ( 
.A1(n_1150),
.A2(n_781),
.B(n_777),
.Y(n_1728)
);

OA21x2_ASAP7_75t_L g1729 ( 
.A1(n_1253),
.A2(n_1134),
.B(n_1120),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1308),
.B(n_817),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1310),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1432),
.Y(n_1732)
);

BUFx12f_ASAP7_75t_L g1733 ( 
.A(n_1205),
.Y(n_1733)
);

BUFx8_ASAP7_75t_L g1734 ( 
.A(n_1171),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1348),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_1444),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1350),
.Y(n_1737)
);

OAI21x1_ASAP7_75t_L g1738 ( 
.A1(n_1151),
.A2(n_782),
.B(n_781),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_SL g1739 ( 
.A(n_1335),
.B(n_990),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1358),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1358),
.Y(n_1741)
);

OA21x2_ASAP7_75t_L g1742 ( 
.A1(n_1253),
.A2(n_797),
.B(n_782),
.Y(n_1742)
);

OAI21x1_ASAP7_75t_L g1743 ( 
.A1(n_1152),
.A2(n_801),
.B(n_797),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1364),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1364),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1269),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1259),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1314),
.B(n_817),
.Y(n_1748)
);

BUFx3_ASAP7_75t_L g1749 ( 
.A(n_1316),
.Y(n_1749)
);

INVx3_ASAP7_75t_L g1750 ( 
.A(n_1384),
.Y(n_1750)
);

BUFx12f_ASAP7_75t_L g1751 ( 
.A(n_1214),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1317),
.B(n_1320),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1478),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1259),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1390),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1390),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1276),
.B(n_821),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1260),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1214),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1552),
.B(n_821),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1392),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1303),
.B(n_821),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1260),
.Y(n_1763)
);

BUFx6f_ASAP7_75t_L g1764 ( 
.A(n_1400),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1321),
.B(n_839),
.Y(n_1765)
);

OA21x2_ASAP7_75t_L g1766 ( 
.A1(n_1262),
.A2(n_805),
.B(n_801),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1400),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1262),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1322),
.Y(n_1769)
);

BUFx12f_ASAP7_75t_L g1770 ( 
.A(n_1238),
.Y(n_1770)
);

BUFx3_ASAP7_75t_L g1771 ( 
.A(n_1324),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1264),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1444),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1264),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1562),
.B(n_839),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1238),
.Y(n_1776)
);

BUFx6f_ASAP7_75t_L g1777 ( 
.A(n_1293),
.Y(n_1777)
);

CKINVDCx11_ASAP7_75t_R g1778 ( 
.A(n_1466),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1265),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1243),
.Y(n_1780)
);

BUFx6f_ASAP7_75t_L g1781 ( 
.A(n_1293),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1265),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1301),
.Y(n_1783)
);

INVx4_ASAP7_75t_L g1784 ( 
.A(n_1301),
.Y(n_1784)
);

OAI22x1_ASAP7_75t_R g1785 ( 
.A1(n_1540),
.A2(n_1017),
.B1(n_1052),
.B2(n_1016),
.Y(n_1785)
);

BUFx3_ASAP7_75t_L g1786 ( 
.A(n_1325),
.Y(n_1786)
);

BUFx12f_ASAP7_75t_L g1787 ( 
.A(n_1243),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1281),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1281),
.Y(n_1789)
);

OAI21x1_ASAP7_75t_L g1790 ( 
.A1(n_1153),
.A2(n_809),
.B(n_805),
.Y(n_1790)
);

INVx5_ASAP7_75t_L g1791 ( 
.A(n_1447),
.Y(n_1791)
);

INVxp33_ASAP7_75t_SL g1792 ( 
.A(n_1199),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1447),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1327),
.Y(n_1794)
);

INVx4_ASAP7_75t_L g1795 ( 
.A(n_1463),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1277),
.Y(n_1796)
);

BUFx8_ASAP7_75t_SL g1797 ( 
.A(n_1472),
.Y(n_1797)
);

OAI21x1_ASAP7_75t_L g1798 ( 
.A1(n_1154),
.A2(n_811),
.B(n_809),
.Y(n_1798)
);

INVx5_ASAP7_75t_L g1799 ( 
.A(n_1463),
.Y(n_1799)
);

BUFx8_ASAP7_75t_L g1800 ( 
.A(n_1341),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1330),
.B(n_839),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1482),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1282),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1482),
.Y(n_1804)
);

INVx4_ASAP7_75t_L g1805 ( 
.A(n_1502),
.Y(n_1805)
);

AOI22x1_ASAP7_75t_SL g1806 ( 
.A1(n_1492),
.A2(n_1122),
.B1(n_1052),
.B2(n_1053),
.Y(n_1806)
);

BUFx8_ASAP7_75t_L g1807 ( 
.A(n_1341),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1305),
.B(n_847),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1502),
.Y(n_1809)
);

AOI22x1_ASAP7_75t_SL g1810 ( 
.A1(n_1495),
.A2(n_1053),
.B1(n_1056),
.B2(n_1017),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1282),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1334),
.B(n_847),
.Y(n_1812)
);

BUFx3_ASAP7_75t_L g1813 ( 
.A(n_1336),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1286),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1277),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1286),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1287),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1522),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1278),
.Y(n_1819)
);

AOI22x1_ASAP7_75t_SL g1820 ( 
.A1(n_1168),
.A2(n_1083),
.B1(n_1056),
.B2(n_1103),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1287),
.Y(n_1821)
);

BUFx3_ASAP7_75t_L g1822 ( 
.A(n_1338),
.Y(n_1822)
);

BUFx3_ASAP7_75t_L g1823 ( 
.A(n_1339),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1288),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1288),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1340),
.B(n_847),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1144),
.A2(n_725),
.B1(n_726),
.B2(n_724),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1278),
.Y(n_1828)
);

BUFx12f_ASAP7_75t_L g1829 ( 
.A(n_1329),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1329),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1333),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1344),
.B(n_1346),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1289),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_SL g1834 ( 
.A1(n_1223),
.A2(n_1083),
.B1(n_1103),
.B2(n_677),
.Y(n_1834)
);

INVx6_ASAP7_75t_L g1835 ( 
.A(n_1394),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1290),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1290),
.Y(n_1837)
);

BUFx6f_ASAP7_75t_L g1838 ( 
.A(n_1522),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1194),
.A2(n_728),
.B1(n_729),
.B2(n_727),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1333),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1361),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1361),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1535),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1194),
.A2(n_1266),
.B1(n_1272),
.B2(n_1246),
.Y(n_1844)
);

INVx5_ASAP7_75t_L g1845 ( 
.A(n_1535),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1347),
.B(n_854),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_1542),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_1542),
.Y(n_1848)
);

BUFx12f_ASAP7_75t_L g1849 ( 
.A(n_1357),
.Y(n_1849)
);

CKINVDCx20_ASAP7_75t_R g1850 ( 
.A(n_1174),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1349),
.B(n_854),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1396),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1397),
.Y(n_1853)
);

OA21x2_ASAP7_75t_L g1854 ( 
.A1(n_1291),
.A2(n_813),
.B(n_811),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1357),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1354),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1543),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1355),
.B(n_854),
.Y(n_1858)
);

BUFx6f_ASAP7_75t_L g1859 ( 
.A(n_1543),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1555),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1375),
.Y(n_1861)
);

BUFx8_ASAP7_75t_SL g1862 ( 
.A(n_1221),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1399),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1401),
.Y(n_1864)
);

BUFx6f_ASAP7_75t_L g1865 ( 
.A(n_1555),
.Y(n_1865)
);

AOI22x1_ASAP7_75t_SL g1866 ( 
.A1(n_1232),
.A2(n_677),
.B1(n_721),
.B2(n_667),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1557),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1405),
.Y(n_1868)
);

BUFx3_ASAP7_75t_L g1869 ( 
.A(n_1356),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1496),
.B(n_870),
.Y(n_1870)
);

OAI22x1_ASAP7_75t_SL g1871 ( 
.A1(n_1246),
.A2(n_771),
.B1(n_730),
.B2(n_721),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1499),
.B(n_870),
.Y(n_1872)
);

BUFx6f_ASAP7_75t_L g1873 ( 
.A(n_1557),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1406),
.Y(n_1874)
);

INVx5_ASAP7_75t_L g1875 ( 
.A(n_1449),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1407),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_1375),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1386),
.Y(n_1878)
);

BUFx2_ASAP7_75t_L g1879 ( 
.A(n_1386),
.Y(n_1879)
);

BUFx6f_ASAP7_75t_L g1880 ( 
.A(n_1408),
.Y(n_1880)
);

INVx6_ASAP7_75t_L g1881 ( 
.A(n_1394),
.Y(n_1881)
);

BUFx12f_ASAP7_75t_L g1882 ( 
.A(n_1424),
.Y(n_1882)
);

CKINVDCx20_ASAP7_75t_R g1883 ( 
.A(n_1242),
.Y(n_1883)
);

INVx6_ASAP7_75t_L g1884 ( 
.A(n_1449),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1410),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1511),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1414),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1415),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1417),
.B(n_870),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1266),
.A2(n_737),
.B1(n_738),
.B2(n_732),
.Y(n_1890)
);

INVx4_ASAP7_75t_L g1891 ( 
.A(n_1158),
.Y(n_1891)
);

INVx3_ASAP7_75t_L g1892 ( 
.A(n_1419),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1420),
.B(n_954),
.Y(n_1893)
);

INVxp67_ASAP7_75t_SL g1894 ( 
.A(n_1511),
.Y(n_1894)
);

OAI22x1_ASAP7_75t_R g1895 ( 
.A1(n_1373),
.A2(n_754),
.B1(n_766),
.B2(n_739),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1422),
.Y(n_1896)
);

BUFx12f_ASAP7_75t_L g1897 ( 
.A(n_1424),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1423),
.B(n_954),
.Y(n_1898)
);

BUFx6f_ASAP7_75t_L g1899 ( 
.A(n_1425),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1159),
.Y(n_1900)
);

BUFx8_ASAP7_75t_L g1901 ( 
.A(n_1403),
.Y(n_1901)
);

OAI22x1_ASAP7_75t_SL g1902 ( 
.A1(n_1272),
.A2(n_722),
.B1(n_730),
.B2(n_667),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1429),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1145),
.Y(n_1904)
);

BUFx8_ASAP7_75t_L g1905 ( 
.A(n_1403),
.Y(n_1905)
);

NOR2x1_ASAP7_75t_L g1906 ( 
.A(n_1698),
.B(n_1145),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1619),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1777),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1777),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1576),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1576),
.B(n_1504),
.Y(n_1911)
);

BUFx6f_ASAP7_75t_L g1912 ( 
.A(n_1619),
.Y(n_1912)
);

INVx3_ASAP7_75t_L g1913 ( 
.A(n_1723),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1591),
.B(n_1163),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1777),
.Y(n_1915)
);

AND2x6_ASAP7_75t_L g1916 ( 
.A(n_1682),
.B(n_1146),
.Y(n_1916)
);

OAI21x1_ASAP7_75t_L g1917 ( 
.A1(n_1571),
.A2(n_1167),
.B(n_1164),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1862),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1704),
.Y(n_1919)
);

INVx3_ASAP7_75t_L g1920 ( 
.A(n_1723),
.Y(n_1920)
);

BUFx6f_ASAP7_75t_L g1921 ( 
.A(n_1619),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1704),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1576),
.B(n_1504),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1777),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1792),
.B(n_1305),
.Y(n_1925)
);

BUFx2_ASAP7_75t_L g1926 ( 
.A(n_1602),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1593),
.B(n_1170),
.Y(n_1927)
);

INVx3_ASAP7_75t_L g1928 ( 
.A(n_1723),
.Y(n_1928)
);

HB1xp67_ASAP7_75t_L g1929 ( 
.A(n_1602),
.Y(n_1929)
);

BUFx2_ASAP7_75t_L g1930 ( 
.A(n_1625),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1717),
.Y(n_1931)
);

XNOR2xp5_ASAP7_75t_L g1932 ( 
.A(n_1664),
.B(n_1574),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1792),
.A2(n_1166),
.B1(n_1353),
.B2(n_1227),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1717),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1571),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1777),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1781),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1904),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1781),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1639),
.B(n_1323),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1781),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1904),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1728),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1781),
.Y(n_1944)
);

INVx3_ASAP7_75t_L g1945 ( 
.A(n_1572),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1781),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_L g1947 ( 
.A(n_1619),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1682),
.B(n_1294),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1620),
.B(n_1172),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1757),
.B(n_1295),
.Y(n_1950)
);

INVxp67_ASAP7_75t_L g1951 ( 
.A(n_1693),
.Y(n_1951)
);

BUFx6f_ASAP7_75t_L g1952 ( 
.A(n_1619),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1728),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1783),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1620),
.B(n_1173),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1783),
.Y(n_1956)
);

BUFx2_ASAP7_75t_L g1957 ( 
.A(n_1625),
.Y(n_1957)
);

INVx5_ASAP7_75t_L g1958 ( 
.A(n_1716),
.Y(n_1958)
);

INVx3_ASAP7_75t_L g1959 ( 
.A(n_1622),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1783),
.Y(n_1960)
);

CKINVDCx16_ASAP7_75t_R g1961 ( 
.A(n_1613),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1738),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1783),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1590),
.B(n_1505),
.Y(n_1964)
);

NAND2xp33_ASAP7_75t_SL g1965 ( 
.A(n_1633),
.B(n_1283),
.Y(n_1965)
);

OAI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1835),
.A2(n_1318),
.B1(n_1332),
.B2(n_1311),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1757),
.B(n_1298),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1783),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1793),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1738),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1743),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1743),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1590),
.B(n_1505),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1590),
.B(n_1506),
.Y(n_1974)
);

XNOR2xp5_ASAP7_75t_L g1975 ( 
.A(n_1721),
.B(n_1439),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1569),
.B(n_1604),
.Y(n_1976)
);

BUFx6f_ASAP7_75t_L g1977 ( 
.A(n_1622),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1793),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1790),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1793),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1622),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1620),
.B(n_1175),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1790),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1681),
.B(n_1176),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1699),
.A2(n_1275),
.B1(n_1413),
.B2(n_771),
.Y(n_1985)
);

CKINVDCx20_ASAP7_75t_R g1986 ( 
.A(n_1850),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1798),
.Y(n_1987)
);

BUFx2_ASAP7_75t_L g1988 ( 
.A(n_1684),
.Y(n_1988)
);

HB1xp67_ASAP7_75t_L g1989 ( 
.A(n_1684),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1793),
.Y(n_1990)
);

INVx2_ASAP7_75t_SL g1991 ( 
.A(n_1835),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1681),
.B(n_1177),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1681),
.B(n_1181),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1622),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1793),
.Y(n_1995)
);

INVx3_ASAP7_75t_L g1996 ( 
.A(n_1572),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_L g1997 ( 
.A(n_1652),
.B(n_1323),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1891),
.B(n_1184),
.Y(n_1998)
);

BUFx6f_ASAP7_75t_L g1999 ( 
.A(n_1622),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1798),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1592),
.B(n_1506),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1900),
.Y(n_2002)
);

AND2x6_ASAP7_75t_L g2003 ( 
.A(n_1592),
.B(n_1146),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1900),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1627),
.Y(n_2005)
);

BUFx6f_ASAP7_75t_L g2006 ( 
.A(n_1624),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1802),
.Y(n_2007)
);

OAI21x1_ASAP7_75t_L g2008 ( 
.A1(n_1854),
.A2(n_1186),
.B(n_1185),
.Y(n_2008)
);

OAI22xp5_ASAP7_75t_SL g2009 ( 
.A1(n_1612),
.A2(n_1834),
.B1(n_1525),
.B2(n_1497),
.Y(n_2009)
);

NAND2xp33_ASAP7_75t_L g2010 ( 
.A(n_1569),
.B(n_1429),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1627),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1718),
.B(n_1263),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1891),
.B(n_1187),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1627),
.Y(n_2014)
);

BUFx6f_ASAP7_75t_L g2015 ( 
.A(n_1624),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1604),
.B(n_1299),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1641),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1641),
.Y(n_2018)
);

INVx5_ASAP7_75t_L g2019 ( 
.A(n_1716),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1802),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1641),
.Y(n_2021)
);

INVx3_ASAP7_75t_L g2022 ( 
.A(n_1575),
.Y(n_2022)
);

OAI21x1_ASAP7_75t_L g2023 ( 
.A1(n_1854),
.A2(n_1190),
.B(n_1188),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1802),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1650),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1802),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_L g2027 ( 
.A(n_1624),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1802),
.Y(n_2028)
);

INVx4_ASAP7_75t_L g2029 ( 
.A(n_1715),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1650),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1575),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1804),
.Y(n_2032)
);

OA21x2_ASAP7_75t_L g2033 ( 
.A1(n_1564),
.A2(n_1190),
.B(n_1188),
.Y(n_2033)
);

BUFx12f_ASAP7_75t_L g2034 ( 
.A(n_1778),
.Y(n_2034)
);

OA21x2_ASAP7_75t_L g2035 ( 
.A1(n_1564),
.A2(n_1192),
.B(n_1191),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1891),
.B(n_1191),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1870),
.B(n_1300),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1870),
.B(n_1304),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1760),
.B(n_1192),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1872),
.B(n_1306),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1650),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1874),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1872),
.B(n_1510),
.Y(n_2043)
);

NAND2x1_ASAP7_75t_L g2044 ( 
.A(n_1715),
.B(n_1111),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1610),
.B(n_1280),
.Y(n_2045)
);

BUFx6f_ASAP7_75t_L g2046 ( 
.A(n_1624),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1760),
.B(n_1193),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1760),
.B(n_1193),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1775),
.B(n_1510),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1566),
.Y(n_2050)
);

BUFx6f_ASAP7_75t_L g2051 ( 
.A(n_1624),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1566),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1568),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1804),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1804),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1568),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_SL g2057 ( 
.A(n_1829),
.B(n_1351),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1775),
.B(n_1592),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_1732),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1804),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1804),
.Y(n_2061)
);

BUFx6f_ASAP7_75t_L g2062 ( 
.A(n_1626),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1775),
.B(n_1715),
.Y(n_2063)
);

OAI21x1_ASAP7_75t_L g2064 ( 
.A1(n_1854),
.A2(n_1196),
.B(n_1195),
.Y(n_2064)
);

AND2x6_ASAP7_75t_L g2065 ( 
.A(n_1715),
.B(n_1195),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_L g2066 ( 
.A(n_1708),
.B(n_1328),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1585),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1715),
.B(n_1196),
.Y(n_2068)
);

BUFx2_ASAP7_75t_L g2069 ( 
.A(n_1883),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1585),
.Y(n_2070)
);

BUFx3_ASAP7_75t_L g2071 ( 
.A(n_1854),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1832),
.B(n_1512),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1618),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1618),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1623),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_1711),
.B(n_1328),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1623),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1832),
.B(n_1512),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1809),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1832),
.B(n_1513),
.Y(n_2080)
);

INVxp67_ASAP7_75t_SL g2081 ( 
.A(n_1710),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1809),
.Y(n_2082)
);

BUFx2_ASAP7_75t_L g2083 ( 
.A(n_1883),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1656),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1835),
.B(n_1881),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1656),
.Y(n_2086)
);

OA21x2_ASAP7_75t_L g2087 ( 
.A1(n_1661),
.A2(n_1198),
.B(n_1197),
.Y(n_2087)
);

BUFx6f_ASAP7_75t_L g2088 ( 
.A(n_1626),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1661),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1809),
.Y(n_2090)
);

NAND2xp33_ASAP7_75t_L g2091 ( 
.A(n_1610),
.B(n_1455),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1698),
.B(n_1197),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1665),
.Y(n_2093)
);

BUFx6f_ASAP7_75t_L g2094 ( 
.A(n_1626),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_1626),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1809),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1628),
.B(n_1366),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_1835),
.B(n_1513),
.Y(n_2098)
);

XOR2xp5_ASAP7_75t_L g2099 ( 
.A(n_1725),
.B(n_1427),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1709),
.B(n_1753),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1665),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_L g2102 ( 
.A(n_1626),
.Y(n_2102)
);

OR2x6_ASAP7_75t_L g2103 ( 
.A(n_1829),
.B(n_954),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_1889),
.B(n_1514),
.Y(n_2104)
);

AO21x2_ASAP7_75t_L g2105 ( 
.A1(n_1649),
.A2(n_1237),
.B(n_1201),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1809),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1709),
.B(n_1198),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1818),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_1637),
.Y(n_2109)
);

OAI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_1881),
.A2(n_1475),
.B1(n_1489),
.B2(n_1428),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1666),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_SL g2112 ( 
.A(n_1628),
.B(n_1385),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1666),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1653),
.B(n_1201),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1668),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1668),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1677),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1881),
.B(n_1514),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1677),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1818),
.Y(n_2120)
);

OAI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_1881),
.A2(n_1382),
.B1(n_1421),
.B2(n_1377),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1680),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1637),
.Y(n_2123)
);

HB1xp67_ASAP7_75t_L g2124 ( 
.A(n_1565),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1680),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1818),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_1583),
.Y(n_2127)
);

BUFx6f_ASAP7_75t_L g2128 ( 
.A(n_1637),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1694),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1655),
.B(n_1202),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1818),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1694),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1696),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1696),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1838),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1838),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1702),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1838),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1838),
.Y(n_2139)
);

BUFx4f_ASAP7_75t_L g2140 ( 
.A(n_1605),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1702),
.Y(n_2141)
);

INVx3_ASAP7_75t_L g2142 ( 
.A(n_1578),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1719),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_SL g2144 ( 
.A(n_1654),
.B(n_1409),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1889),
.B(n_1516),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1838),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_1578),
.Y(n_2147)
);

OAI21x1_ASAP7_75t_L g2148 ( 
.A1(n_1667),
.A2(n_1207),
.B(n_1202),
.Y(n_2148)
);

BUFx3_ASAP7_75t_L g2149 ( 
.A(n_1710),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1843),
.Y(n_2150)
);

HB1xp67_ASAP7_75t_L g2151 ( 
.A(n_1596),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1719),
.Y(n_2152)
);

INVx4_ASAP7_75t_L g2153 ( 
.A(n_1843),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1722),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1894),
.B(n_1207),
.Y(n_2155)
);

BUFx6f_ASAP7_75t_L g2156 ( 
.A(n_1637),
.Y(n_2156)
);

INVx3_ASAP7_75t_L g2157 ( 
.A(n_1578),
.Y(n_2157)
);

BUFx8_ASAP7_75t_L g2158 ( 
.A(n_1579),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1722),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1843),
.Y(n_2160)
);

BUFx6f_ASAP7_75t_L g2161 ( 
.A(n_1637),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1726),
.Y(n_2162)
);

INVxp67_ASAP7_75t_L g2163 ( 
.A(n_1739),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1843),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1843),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1726),
.Y(n_2166)
);

BUFx3_ASAP7_75t_L g2167 ( 
.A(n_1710),
.Y(n_2167)
);

HB1xp67_ASAP7_75t_L g2168 ( 
.A(n_1638),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1747),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1747),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_1889),
.B(n_1516),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1654),
.B(n_1208),
.Y(n_2172)
);

AND2x4_ASAP7_75t_L g2173 ( 
.A(n_1893),
.B(n_1517),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1754),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_1658),
.B(n_1736),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1754),
.Y(n_2176)
);

INVx3_ASAP7_75t_L g2177 ( 
.A(n_1578),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1758),
.Y(n_2178)
);

INVx6_ASAP7_75t_L g2179 ( 
.A(n_1710),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1658),
.B(n_1208),
.Y(n_2180)
);

BUFx8_ASAP7_75t_L g2181 ( 
.A(n_1579),
.Y(n_2181)
);

INVx3_ASAP7_75t_L g2182 ( 
.A(n_1582),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1847),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1758),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1847),
.Y(n_2185)
);

BUFx3_ASAP7_75t_L g2186 ( 
.A(n_1710),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1736),
.B(n_1209),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1763),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_1893),
.B(n_1898),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1763),
.Y(n_2190)
);

CKINVDCx8_ASAP7_75t_R g2191 ( 
.A(n_1673),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_1609),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1768),
.Y(n_2193)
);

BUFx3_ASAP7_75t_L g2194 ( 
.A(n_1731),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_SL g2195 ( 
.A(n_1849),
.B(n_1456),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1847),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1768),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1772),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1772),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1774),
.Y(n_2200)
);

AND2x4_ASAP7_75t_L g2201 ( 
.A(n_1893),
.B(n_1517),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1774),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1847),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1773),
.B(n_1210),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_1640),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_1640),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_1898),
.B(n_1518),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1848),
.Y(n_2208)
);

OAI22xp5_ASAP7_75t_SL g2209 ( 
.A1(n_1647),
.A2(n_795),
.B1(n_800),
.B2(n_722),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1779),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_1898),
.B(n_1518),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1779),
.Y(n_2212)
);

AND2x4_ASAP7_75t_L g2213 ( 
.A(n_1603),
.B(n_1519),
.Y(n_2213)
);

CKINVDCx6p67_ASAP7_75t_R g2214 ( 
.A(n_1567),
.Y(n_2214)
);

BUFx6f_ASAP7_75t_L g2215 ( 
.A(n_1640),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1782),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_1731),
.B(n_1749),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1782),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_1848),
.Y(n_2219)
);

AND2x4_ASAP7_75t_L g2220 ( 
.A(n_1851),
.B(n_1519),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_SL g2221 ( 
.A(n_1886),
.B(n_1459),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1811),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_1582),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1848),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_1749),
.B(n_1520),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_1640),
.Y(n_2226)
);

AND2x4_ASAP7_75t_L g2227 ( 
.A(n_1851),
.B(n_1520),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_1769),
.B(n_1521),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_1769),
.B(n_1521),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1811),
.Y(n_2230)
);

AND2x6_ASAP7_75t_L g2231 ( 
.A(n_1762),
.B(n_1210),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1814),
.Y(n_2232)
);

AND2x6_ASAP7_75t_L g2233 ( 
.A(n_1808),
.B(n_1211),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1848),
.Y(n_2234)
);

HB1xp67_ASAP7_75t_L g2235 ( 
.A(n_1648),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_1771),
.B(n_1523),
.Y(n_2236)
);

AND2x4_ASAP7_75t_L g2237 ( 
.A(n_1851),
.B(n_1523),
.Y(n_2237)
);

AND2x4_ASAP7_75t_L g2238 ( 
.A(n_1858),
.B(n_1524),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1814),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1816),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1848),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_1640),
.Y(n_2242)
);

NAND2xp33_ASAP7_75t_L g2243 ( 
.A(n_1886),
.B(n_1455),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_1858),
.B(n_1524),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1816),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1859),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1859),
.Y(n_2247)
);

OAI22xp5_ASAP7_75t_SL g2248 ( 
.A1(n_1647),
.A2(n_795),
.B1(n_807),
.B2(n_800),
.Y(n_2248)
);

NOR2xp33_ASAP7_75t_L g2249 ( 
.A(n_1703),
.B(n_1377),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1817),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_1858),
.B(n_1526),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_1771),
.B(n_1526),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1817),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1821),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_1859),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1821),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1784),
.B(n_1211),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1859),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1833),
.Y(n_2259)
);

OAI22xp5_ASAP7_75t_L g2260 ( 
.A1(n_1580),
.A2(n_1421),
.B1(n_1470),
.B2(n_1382),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1833),
.Y(n_2261)
);

INVx3_ASAP7_75t_L g2262 ( 
.A(n_1582),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_1643),
.Y(n_2263)
);

BUFx2_ASAP7_75t_L g2264 ( 
.A(n_1598),
.Y(n_2264)
);

CKINVDCx5p33_ASAP7_75t_R g2265 ( 
.A(n_1621),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_1784),
.B(n_1212),
.Y(n_2266)
);

INVx4_ASAP7_75t_L g2267 ( 
.A(n_1859),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1836),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_1865),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1836),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1865),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1837),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1837),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1841),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_1786),
.B(n_1527),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1841),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1784),
.B(n_1212),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_1643),
.Y(n_2278)
);

AND2x6_ASAP7_75t_L g2279 ( 
.A(n_1786),
.B(n_1213),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_L g2280 ( 
.A(n_1827),
.B(n_1470),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1865),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_1865),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1865),
.Y(n_2283)
);

BUFx6f_ASAP7_75t_L g2284 ( 
.A(n_1643),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1788),
.Y(n_2285)
);

AND2x4_ASAP7_75t_L g2286 ( 
.A(n_1794),
.B(n_1527),
.Y(n_2286)
);

BUFx6f_ASAP7_75t_L g2287 ( 
.A(n_1643),
.Y(n_2287)
);

BUFx2_ASAP7_75t_L g2288 ( 
.A(n_1598),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_1795),
.B(n_1215),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1788),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1788),
.Y(n_2291)
);

INVx4_ASAP7_75t_L g2292 ( 
.A(n_1873),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_1873),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1789),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1795),
.B(n_1805),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_1789),
.Y(n_2296)
);

AND2x4_ASAP7_75t_L g2297 ( 
.A(n_1794),
.B(n_1528),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_1813),
.B(n_1822),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_1805),
.B(n_1215),
.Y(n_2299)
);

AND2x4_ASAP7_75t_L g2300 ( 
.A(n_1813),
.B(n_1528),
.Y(n_2300)
);

XNOR2x2_ASAP7_75t_L g2301 ( 
.A(n_1844),
.B(n_807),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1873),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_1822),
.B(n_1529),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1803),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_1805),
.B(n_1216),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1803),
.Y(n_2306)
);

HB1xp67_ASAP7_75t_L g2307 ( 
.A(n_1678),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_1823),
.B(n_1529),
.Y(n_2308)
);

INVx3_ASAP7_75t_L g2309 ( 
.A(n_1586),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1803),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1910),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2033),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_2085),
.B(n_1875),
.Y(n_2313)
);

OAI21xp33_ASAP7_75t_SL g2314 ( 
.A1(n_1976),
.A2(n_976),
.B(n_972),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2231),
.B(n_1875),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1910),
.Y(n_2316)
);

INVx2_ASAP7_75t_SL g2317 ( 
.A(n_2085),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2033),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2231),
.B(n_1875),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2033),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2033),
.Y(n_2321)
);

BUFx2_ASAP7_75t_L g2322 ( 
.A(n_1951),
.Y(n_2322)
);

INVx5_ASAP7_75t_L g2323 ( 
.A(n_2003),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1910),
.Y(n_2324)
);

INVx2_ASAP7_75t_SL g2325 ( 
.A(n_2098),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_1976),
.B(n_1875),
.Y(n_2326)
);

CKINVDCx6p67_ASAP7_75t_R g2327 ( 
.A(n_2034),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_1938),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2035),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2035),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2035),
.Y(n_2331)
);

HB1xp67_ASAP7_75t_L g2332 ( 
.A(n_1926),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1938),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2035),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2087),
.Y(n_2335)
);

BUFx4f_ASAP7_75t_L g2336 ( 
.A(n_2231),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_1942),
.Y(n_2337)
);

INVx6_ASAP7_75t_L g2338 ( 
.A(n_2179),
.Y(n_2338)
);

BUFx10_ASAP7_75t_L g2339 ( 
.A(n_1925),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2087),
.Y(n_2340)
);

NOR3xp33_ASAP7_75t_L g2341 ( 
.A(n_2260),
.B(n_1815),
.C(n_1796),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2087),
.Y(n_2342)
);

NAND2xp33_ASAP7_75t_L g2343 ( 
.A(n_1916),
.B(n_1746),
.Y(n_2343)
);

INVx1_ASAP7_75t_SL g2344 ( 
.A(n_1986),
.Y(n_2344)
);

INVx3_ASAP7_75t_L g2345 ( 
.A(n_2087),
.Y(n_2345)
);

BUFx6f_ASAP7_75t_L g2346 ( 
.A(n_2003),
.Y(n_2346)
);

INVx2_ASAP7_75t_SL g2347 ( 
.A(n_2098),
.Y(n_2347)
);

INVx2_ASAP7_75t_SL g2348 ( 
.A(n_2118),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1942),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_1991),
.B(n_1819),
.Y(n_2350)
);

INVxp67_ASAP7_75t_L g2351 ( 
.A(n_2059),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2049),
.B(n_1823),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2050),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2050),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2052),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2049),
.B(n_1856),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2052),
.Y(n_2357)
);

XNOR2x2_ASAP7_75t_L g2358 ( 
.A(n_2301),
.B(n_897),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_SL g2359 ( 
.A(n_1991),
.B(n_1819),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2053),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2053),
.Y(n_2361)
);

BUFx3_ASAP7_75t_L g2362 ( 
.A(n_2003),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2056),
.Y(n_2363)
);

BUFx6f_ASAP7_75t_L g2364 ( 
.A(n_2003),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2043),
.B(n_2016),
.Y(n_2365)
);

BUFx3_ASAP7_75t_L g2366 ( 
.A(n_2003),
.Y(n_2366)
);

INVx3_ASAP7_75t_L g2367 ( 
.A(n_1919),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2056),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_1940),
.B(n_1746),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2067),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2067),
.Y(n_2371)
);

BUFx3_ASAP7_75t_L g2372 ( 
.A(n_2003),
.Y(n_2372)
);

INVx2_ASAP7_75t_SL g2373 ( 
.A(n_2118),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_1935),
.Y(n_2374)
);

OAI22xp33_ASAP7_75t_L g2375 ( 
.A1(n_1933),
.A2(n_1636),
.B1(n_1724),
.B2(n_1645),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_1935),
.Y(n_2376)
);

BUFx4f_ASAP7_75t_L g2377 ( 
.A(n_2231),
.Y(n_2377)
);

OAI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_2058),
.A2(n_1855),
.B1(n_1861),
.B2(n_1840),
.Y(n_2378)
);

INVx1_ASAP7_75t_SL g2379 ( 
.A(n_2069),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2043),
.B(n_1856),
.Y(n_2380)
);

AND2x4_ASAP7_75t_L g2381 ( 
.A(n_2189),
.B(n_1869),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_1919),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2070),
.Y(n_2383)
);

OR2x2_ASAP7_75t_L g2384 ( 
.A(n_1933),
.B(n_1673),
.Y(n_2384)
);

OR2x6_ASAP7_75t_L g2385 ( 
.A(n_2189),
.B(n_1849),
.Y(n_2385)
);

BUFx2_ASAP7_75t_L g2386 ( 
.A(n_2163),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2070),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_1922),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2073),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_1922),
.Y(n_2390)
);

BUFx10_ASAP7_75t_L g2391 ( 
.A(n_2249),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2231),
.B(n_1605),
.Y(n_2392)
);

BUFx3_ASAP7_75t_L g2393 ( 
.A(n_2003),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2073),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2231),
.B(n_1605),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_1931),
.Y(n_2396)
);

INVx1_ASAP7_75t_SL g2397 ( 
.A(n_2069),
.Y(n_2397)
);

HB1xp67_ASAP7_75t_L g2398 ( 
.A(n_1926),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2074),
.Y(n_2399)
);

INVx3_ASAP7_75t_L g2400 ( 
.A(n_1931),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_SL g2401 ( 
.A(n_1997),
.B(n_1830),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2074),
.Y(n_2402)
);

BUFx3_ASAP7_75t_L g2403 ( 
.A(n_1916),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2075),
.Y(n_2404)
);

NOR2x1p5_ASAP7_75t_L g2405 ( 
.A(n_2214),
.B(n_1567),
.Y(n_2405)
);

INVx4_ASAP7_75t_L g2406 ( 
.A(n_1913),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2075),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_SL g2408 ( 
.A(n_2066),
.B(n_1828),
.Y(n_2408)
);

NAND2xp33_ASAP7_75t_R g2409 ( 
.A(n_2083),
.B(n_1828),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2077),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2077),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2084),
.Y(n_2412)
);

INVx3_ASAP7_75t_L g2413 ( 
.A(n_1934),
.Y(n_2413)
);

INVx3_ASAP7_75t_L g2414 ( 
.A(n_1934),
.Y(n_2414)
);

BUFx6f_ASAP7_75t_L g2415 ( 
.A(n_2071),
.Y(n_2415)
);

INVx3_ASAP7_75t_L g2416 ( 
.A(n_1917),
.Y(n_2416)
);

INVx3_ASAP7_75t_L g2417 ( 
.A(n_1917),
.Y(n_2417)
);

NOR2xp33_ASAP7_75t_R g2418 ( 
.A(n_1918),
.B(n_1903),
.Y(n_2418)
);

BUFx6f_ASAP7_75t_L g2419 ( 
.A(n_2071),
.Y(n_2419)
);

INVxp67_ASAP7_75t_SL g2420 ( 
.A(n_1913),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2084),
.Y(n_2421)
);

INVx4_ASAP7_75t_L g2422 ( 
.A(n_1913),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2086),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2233),
.B(n_1605),
.Y(n_2424)
);

INVx2_ASAP7_75t_SL g2425 ( 
.A(n_2217),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2233),
.B(n_1675),
.Y(n_2426)
);

BUFx6f_ASAP7_75t_L g2427 ( 
.A(n_2071),
.Y(n_2427)
);

NOR2xp33_ASAP7_75t_L g2428 ( 
.A(n_2076),
.B(n_1830),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2233),
.B(n_1675),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2086),
.Y(n_2430)
);

BUFx3_ASAP7_75t_L g2431 ( 
.A(n_1916),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2089),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2089),
.Y(n_2433)
);

NAND2xp33_ASAP7_75t_SL g2434 ( 
.A(n_1966),
.B(n_1877),
.Y(n_2434)
);

OAI22xp33_ASAP7_75t_L g2435 ( 
.A1(n_1985),
.A2(n_1839),
.B1(n_1890),
.B2(n_1630),
.Y(n_2435)
);

BUFx3_ASAP7_75t_L g2436 ( 
.A(n_1916),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2093),
.Y(n_2437)
);

BUFx3_ASAP7_75t_L g2438 ( 
.A(n_1916),
.Y(n_2438)
);

OR2x6_ASAP7_75t_L g2439 ( 
.A(n_2103),
.B(n_1882),
.Y(n_2439)
);

INVx5_ASAP7_75t_L g2440 ( 
.A(n_2065),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2093),
.Y(n_2441)
);

AOI22xp5_ASAP7_75t_L g2442 ( 
.A1(n_2233),
.A2(n_1713),
.B1(n_1729),
.B2(n_1675),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2101),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2016),
.B(n_1869),
.Y(n_2444)
);

AND3x2_ASAP7_75t_L g2445 ( 
.A(n_2264),
.B(n_1133),
.C(n_758),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2101),
.Y(n_2446)
);

INVxp33_ASAP7_75t_L g2447 ( 
.A(n_2209),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2111),
.Y(n_2448)
);

AOI21x1_ASAP7_75t_L g2449 ( 
.A1(n_1943),
.A2(n_1713),
.B(n_1675),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_2121),
.B(n_1877),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2233),
.B(n_1713),
.Y(n_2451)
);

CKINVDCx5p33_ASAP7_75t_R g2452 ( 
.A(n_2192),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_1948),
.B(n_1796),
.Y(n_2453)
);

OR2x2_ASAP7_75t_L g2454 ( 
.A(n_1985),
.B(n_1705),
.Y(n_2454)
);

INVx3_ASAP7_75t_L g2455 ( 
.A(n_1911),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2023),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2111),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2233),
.B(n_1713),
.Y(n_2458)
);

BUFx6f_ASAP7_75t_L g2459 ( 
.A(n_2140),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2113),
.Y(n_2460)
);

BUFx3_ASAP7_75t_L g2461 ( 
.A(n_1916),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2023),
.Y(n_2462)
);

AOI22xp33_ASAP7_75t_L g2463 ( 
.A1(n_2233),
.A2(n_1916),
.B1(n_1923),
.B2(n_1911),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2113),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_SL g2465 ( 
.A(n_2110),
.B(n_1878),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_2192),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2064),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2115),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2115),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2116),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2064),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2005),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2116),
.Y(n_2473)
);

INVx1_ASAP7_75t_SL g2474 ( 
.A(n_2083),
.Y(n_2474)
);

AOI22xp33_ASAP7_75t_L g2475 ( 
.A1(n_1911),
.A2(n_1742),
.B1(n_1766),
.B2(n_1729),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2005),
.Y(n_2476)
);

NAND2xp33_ASAP7_75t_SL g2477 ( 
.A(n_2012),
.B(n_1878),
.Y(n_2477)
);

BUFx8_ASAP7_75t_SL g2478 ( 
.A(n_2034),
.Y(n_2478)
);

BUFx10_ASAP7_75t_L g2479 ( 
.A(n_2280),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2011),
.Y(n_2480)
);

AND3x2_ASAP7_75t_L g2481 ( 
.A(n_2264),
.B(n_1133),
.C(n_758),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2117),
.Y(n_2482)
);

INVx2_ASAP7_75t_SL g2483 ( 
.A(n_2217),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_2100),
.B(n_1903),
.Y(n_2484)
);

OR2x6_ASAP7_75t_L g2485 ( 
.A(n_2103),
.B(n_1882),
.Y(n_2485)
);

INVx8_ASAP7_75t_L g2486 ( 
.A(n_2279),
.Y(n_2486)
);

INVx4_ASAP7_75t_L g2487 ( 
.A(n_1920),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_SL g2488 ( 
.A(n_2194),
.B(n_1815),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2011),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2014),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2117),
.Y(n_2491)
);

BUFx10_ASAP7_75t_L g2492 ( 
.A(n_2265),
.Y(n_2492)
);

AND2x6_ASAP7_75t_L g2493 ( 
.A(n_1943),
.B(n_813),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2119),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_SL g2495 ( 
.A(n_2194),
.B(n_1831),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2119),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2122),
.Y(n_2497)
);

CKINVDCx11_ASAP7_75t_R g2498 ( 
.A(n_2214),
.Y(n_2498)
);

INVx4_ASAP7_75t_L g2499 ( 
.A(n_1928),
.Y(n_2499)
);

AND3x2_ASAP7_75t_L g2500 ( 
.A(n_2288),
.B(n_1776),
.C(n_1705),
.Y(n_2500)
);

INVx2_ASAP7_75t_SL g2501 ( 
.A(n_2298),
.Y(n_2501)
);

OAI22x1_ASAP7_75t_L g2502 ( 
.A1(n_1932),
.A2(n_1183),
.B1(n_1200),
.B2(n_1149),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_SL g2503 ( 
.A(n_1961),
.B(n_1897),
.Y(n_2503)
);

INVx2_ASAP7_75t_SL g2504 ( 
.A(n_2298),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_1928),
.B(n_1742),
.Y(n_2505)
);

OAI21xp33_ASAP7_75t_SL g2506 ( 
.A1(n_2039),
.A2(n_976),
.B(n_972),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2122),
.Y(n_2507)
);

BUFx6f_ASAP7_75t_L g2508 ( 
.A(n_2140),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2125),
.Y(n_2509)
);

INVx4_ASAP7_75t_L g2510 ( 
.A(n_1928),
.Y(n_2510)
);

INVx1_ASAP7_75t_SL g2511 ( 
.A(n_2124),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2125),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2129),
.Y(n_2513)
);

INVx2_ASAP7_75t_SL g2514 ( 
.A(n_1948),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2129),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_SL g2516 ( 
.A(n_2194),
.B(n_1831),
.Y(n_2516)
);

AOI22xp33_ASAP7_75t_L g2517 ( 
.A1(n_1911),
.A2(n_1766),
.B1(n_1742),
.B2(n_1494),
.Y(n_2517)
);

OA22x2_ASAP7_75t_L g2518 ( 
.A1(n_2009),
.A2(n_1255),
.B1(n_1345),
.B2(n_1326),
.Y(n_2518)
);

BUFx2_ASAP7_75t_L g2519 ( 
.A(n_2127),
.Y(n_2519)
);

INVx3_ASAP7_75t_L g2520 ( 
.A(n_1923),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2132),
.Y(n_2521)
);

AOI22xp5_ASAP7_75t_L g2522 ( 
.A1(n_2105),
.A2(n_1766),
.B1(n_1742),
.B2(n_1902),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2132),
.Y(n_2523)
);

BUFx3_ASAP7_75t_L g2524 ( 
.A(n_2279),
.Y(n_2524)
);

BUFx6f_ASAP7_75t_SL g2525 ( 
.A(n_2103),
.Y(n_2525)
);

INVx8_ASAP7_75t_L g2526 ( 
.A(n_2279),
.Y(n_2526)
);

CKINVDCx5p33_ASAP7_75t_R g2527 ( 
.A(n_2265),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2133),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2133),
.Y(n_2529)
);

OR2x6_ASAP7_75t_L g2530 ( 
.A(n_2103),
.B(n_1897),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2134),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2172),
.B(n_1766),
.Y(n_2532)
);

NOR2xp33_ASAP7_75t_L g2533 ( 
.A(n_1930),
.B(n_1879),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2134),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2137),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2137),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2141),
.Y(n_2537)
);

BUFx2_ASAP7_75t_L g2538 ( 
.A(n_2151),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2141),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2143),
.Y(n_2540)
);

AOI22xp5_ASAP7_75t_L g2541 ( 
.A1(n_2105),
.A2(n_1871),
.B1(n_1473),
.B2(n_1503),
.Y(n_2541)
);

INVx5_ASAP7_75t_L g2542 ( 
.A(n_2065),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2143),
.Y(n_2543)
);

BUFx6f_ASAP7_75t_L g2544 ( 
.A(n_2140),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2152),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2152),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2154),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2154),
.Y(n_2548)
);

NAND2xp33_ASAP7_75t_SL g2549 ( 
.A(n_2112),
.B(n_1879),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2159),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2180),
.B(n_2187),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2159),
.Y(n_2552)
);

INVx4_ASAP7_75t_L g2553 ( 
.A(n_2029),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_1950),
.B(n_1884),
.Y(n_2554)
);

CKINVDCx5p33_ASAP7_75t_R g2555 ( 
.A(n_1961),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_1950),
.B(n_1884),
.Y(n_2556)
);

INVx3_ASAP7_75t_L g2557 ( 
.A(n_1923),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2162),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_SL g2559 ( 
.A(n_1930),
.B(n_1509),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2162),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2166),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2166),
.Y(n_2562)
);

INVx1_ASAP7_75t_SL g2563 ( 
.A(n_2168),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_SL g2564 ( 
.A(n_1957),
.B(n_1776),
.Y(n_2564)
);

INVxp67_ASAP7_75t_SL g2565 ( 
.A(n_2063),
.Y(n_2565)
);

AOI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2105),
.A2(n_1473),
.B1(n_1503),
.B2(n_1494),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2169),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_1957),
.B(n_1780),
.Y(n_2568)
);

CKINVDCx6p67_ASAP7_75t_R g2569 ( 
.A(n_2288),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2169),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2170),
.Y(n_2571)
);

INVx5_ASAP7_75t_L g2572 ( 
.A(n_2065),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2170),
.Y(n_2573)
);

CKINVDCx6p67_ASAP7_75t_R g2574 ( 
.A(n_2103),
.Y(n_2574)
);

CKINVDCx20_ASAP7_75t_R g2575 ( 
.A(n_2158),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2204),
.B(n_1588),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2174),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_SL g2578 ( 
.A(n_1988),
.B(n_1780),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2174),
.Y(n_2579)
);

BUFx2_ASAP7_75t_L g2580 ( 
.A(n_2235),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2176),
.Y(n_2581)
);

INVx11_ASAP7_75t_L g2582 ( 
.A(n_2158),
.Y(n_2582)
);

NAND2xp33_ASAP7_75t_SL g2583 ( 
.A(n_2144),
.B(n_1688),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2176),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2155),
.B(n_1588),
.Y(n_2585)
);

INVxp33_ASAP7_75t_SL g2586 ( 
.A(n_2195),
.Y(n_2586)
);

NOR2x1p5_ASAP7_75t_L g2587 ( 
.A(n_2044),
.B(n_1646),
.Y(n_2587)
);

AOI22xp33_ASAP7_75t_L g2588 ( 
.A1(n_1923),
.A2(n_1536),
.B1(n_976),
.B2(n_994),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2047),
.B(n_1634),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2178),
.Y(n_2590)
);

BUFx3_ASAP7_75t_L g2591 ( 
.A(n_2279),
.Y(n_2591)
);

OAI22xp5_ASAP7_75t_L g2592 ( 
.A1(n_2048),
.A2(n_1759),
.B1(n_1474),
.B2(n_1480),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2178),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2184),
.Y(n_2594)
);

OR2x2_ASAP7_75t_L g2595 ( 
.A(n_1965),
.B(n_1584),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2184),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_SL g2597 ( 
.A(n_1988),
.B(n_1458),
.Y(n_2597)
);

AND2x4_ASAP7_75t_L g2598 ( 
.A(n_1964),
.B(n_1973),
.Y(n_2598)
);

INVxp33_ASAP7_75t_L g2599 ( 
.A(n_2209),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_SL g2600 ( 
.A(n_1967),
.B(n_1458),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_1964),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2014),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2188),
.Y(n_2603)
);

NOR2xp33_ASAP7_75t_L g2604 ( 
.A(n_2221),
.B(n_1536),
.Y(n_2604)
);

NOR3xp33_ASAP7_75t_L g2605 ( 
.A(n_2009),
.B(n_1642),
.C(n_1563),
.Y(n_2605)
);

NAND2xp33_ASAP7_75t_SL g2606 ( 
.A(n_2045),
.B(n_1474),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2092),
.B(n_1634),
.Y(n_2607)
);

AND2x6_ASAP7_75t_L g2608 ( 
.A(n_1953),
.B(n_822),
.Y(n_2608)
);

INVxp67_ASAP7_75t_SL g2609 ( 
.A(n_2295),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2188),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2017),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2107),
.B(n_1634),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2017),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2018),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2190),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_1964),
.B(n_1674),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_SL g2617 ( 
.A(n_1967),
.B(n_1480),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_SL g2618 ( 
.A(n_1964),
.B(n_1973),
.Y(n_2618)
);

OAI22xp33_ASAP7_75t_SL g2619 ( 
.A1(n_1949),
.A2(n_898),
.B1(n_1039),
.B2(n_897),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2018),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2021),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_1973),
.B(n_1674),
.Y(n_2622)
);

AO21x2_ASAP7_75t_L g2623 ( 
.A1(n_1953),
.A2(n_1730),
.B(n_1695),
.Y(n_2623)
);

NOR2xp33_ASAP7_75t_SL g2624 ( 
.A(n_2057),
.B(n_1581),
.Y(n_2624)
);

BUFx10_ASAP7_75t_L g2625 ( 
.A(n_2279),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2021),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2190),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2025),
.Y(n_2628)
);

INVx3_ASAP7_75t_L g2629 ( 
.A(n_1973),
.Y(n_2629)
);

AOI21x1_ASAP7_75t_L g2630 ( 
.A1(n_1962),
.A2(n_1825),
.B(n_1824),
.Y(n_2630)
);

AND2x6_ASAP7_75t_L g2631 ( 
.A(n_1962),
.B(n_822),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2193),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2193),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2197),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2197),
.Y(n_2635)
);

BUFx6f_ASAP7_75t_L g2636 ( 
.A(n_2149),
.Y(n_2636)
);

INVx2_ASAP7_75t_SL g2637 ( 
.A(n_2037),
.Y(n_2637)
);

CKINVDCx5p33_ASAP7_75t_R g2638 ( 
.A(n_2158),
.Y(n_2638)
);

BUFx6f_ASAP7_75t_L g2639 ( 
.A(n_2149),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2198),
.Y(n_2640)
);

BUFx3_ASAP7_75t_L g2641 ( 
.A(n_2279),
.Y(n_2641)
);

BUFx6f_ASAP7_75t_L g2642 ( 
.A(n_2149),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2198),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2199),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2199),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2200),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_SL g2647 ( 
.A(n_1974),
.B(n_1484),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2200),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_1974),
.B(n_1674),
.Y(n_2649)
);

NAND2xp33_ASAP7_75t_L g2650 ( 
.A(n_2279),
.B(n_1484),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_2158),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2202),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2202),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2210),
.Y(n_2654)
);

BUFx2_ASAP7_75t_L g2655 ( 
.A(n_2307),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2210),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2212),
.Y(n_2657)
);

INVx3_ASAP7_75t_L g2658 ( 
.A(n_1974),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2212),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_SL g2660 ( 
.A(n_2001),
.B(n_1486),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2216),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2216),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2218),
.Y(n_2663)
);

INVx2_ASAP7_75t_SL g2664 ( 
.A(n_2037),
.Y(n_2664)
);

BUFx6f_ASAP7_75t_L g2665 ( 
.A(n_2167),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2025),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2030),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_SL g2668 ( 
.A(n_2001),
.B(n_1486),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2218),
.Y(n_2669)
);

INVx3_ASAP7_75t_L g2670 ( 
.A(n_2001),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2222),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2030),
.Y(n_2672)
);

INVx3_ASAP7_75t_L g2673 ( 
.A(n_2001),
.Y(n_2673)
);

BUFx6f_ASAP7_75t_SL g2674 ( 
.A(n_2213),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2114),
.B(n_1679),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_SL g2676 ( 
.A(n_2220),
.B(n_2227),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2041),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2130),
.B(n_1679),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2038),
.B(n_1884),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2041),
.Y(n_2680)
);

INVxp67_ASAP7_75t_SL g2681 ( 
.A(n_2068),
.Y(n_2681)
);

INVxp33_ASAP7_75t_L g2682 ( 
.A(n_2248),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2008),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2008),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_1955),
.B(n_1679),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2222),
.Y(n_2686)
);

INVx4_ASAP7_75t_L g2687 ( 
.A(n_2029),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2230),
.Y(n_2688)
);

BUFx4f_ASAP7_75t_L g2689 ( 
.A(n_2213),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2038),
.B(n_1884),
.Y(n_2690)
);

INVx3_ASAP7_75t_L g2691 ( 
.A(n_2104),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2230),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2232),
.Y(n_2693)
);

AOI22xp33_ASAP7_75t_L g2694 ( 
.A1(n_1982),
.A2(n_1074),
.B1(n_994),
.B2(n_1257),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2232),
.Y(n_2695)
);

INVx4_ASAP7_75t_L g2696 ( 
.A(n_2029),
.Y(n_2696)
);

NAND2xp33_ASAP7_75t_L g2697 ( 
.A(n_1906),
.B(n_1490),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_SL g2698 ( 
.A(n_2220),
.B(n_2227),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2239),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2239),
.Y(n_2700)
);

OR2x2_ASAP7_75t_L g2701 ( 
.A(n_2301),
.B(n_1493),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2240),
.Y(n_2702)
);

AND2x6_ASAP7_75t_L g2703 ( 
.A(n_1970),
.B(n_824),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2240),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_SL g2705 ( 
.A(n_2220),
.B(n_2227),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_SL g2706 ( 
.A(n_2227),
.B(n_2237),
.Y(n_2706)
);

NOR2xp33_ASAP7_75t_L g2707 ( 
.A(n_2097),
.B(n_1493),
.Y(n_2707)
);

BUFx2_ASAP7_75t_L g2708 ( 
.A(n_1929),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2245),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2245),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_SL g2711 ( 
.A(n_2237),
.B(n_1500),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2250),
.Y(n_2712)
);

CKINVDCx5p33_ASAP7_75t_R g2713 ( 
.A(n_2181),
.Y(n_2713)
);

INVx2_ASAP7_75t_SL g2714 ( 
.A(n_2040),
.Y(n_2714)
);

INVx3_ASAP7_75t_L g2715 ( 
.A(n_2104),
.Y(n_2715)
);

NOR2xp33_ASAP7_75t_L g2716 ( 
.A(n_1989),
.B(n_1500),
.Y(n_2716)
);

INVx3_ASAP7_75t_L g2717 ( 
.A(n_2104),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_1984),
.B(n_1570),
.Y(n_2718)
);

INVxp33_ASAP7_75t_L g2719 ( 
.A(n_2248),
.Y(n_2719)
);

INVx1_ASAP7_75t_SL g2720 ( 
.A(n_2040),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2072),
.B(n_1292),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_1992),
.B(n_1993),
.Y(n_2722)
);

NAND2xp33_ASAP7_75t_L g2723 ( 
.A(n_1906),
.B(n_1507),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2250),
.Y(n_2724)
);

NAND2xp33_ASAP7_75t_L g2725 ( 
.A(n_2065),
.B(n_1507),
.Y(n_2725)
);

NAND3xp33_ASAP7_75t_L g2726 ( 
.A(n_2010),
.B(n_1765),
.C(n_1748),
.Y(n_2726)
);

AND2x2_ASAP7_75t_L g2727 ( 
.A(n_2072),
.B(n_1309),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2253),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2181),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2253),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2254),
.Y(n_2731)
);

AOI21x1_ASAP7_75t_L g2732 ( 
.A1(n_1970),
.A2(n_1825),
.B(n_1824),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_1914),
.B(n_1570),
.Y(n_2733)
);

BUFx3_ASAP7_75t_L g2734 ( 
.A(n_2104),
.Y(n_2734)
);

INVx5_ASAP7_75t_L g2735 ( 
.A(n_2065),
.Y(n_2735)
);

AND2x6_ASAP7_75t_L g2736 ( 
.A(n_1971),
.B(n_824),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2254),
.Y(n_2737)
);

BUFx3_ASAP7_75t_L g2738 ( 
.A(n_2171),
.Y(n_2738)
);

INVx2_ASAP7_75t_SL g2739 ( 
.A(n_2145),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_2478),
.Y(n_2740)
);

BUFx6f_ASAP7_75t_L g2741 ( 
.A(n_2415),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2311),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2311),
.Y(n_2743)
);

BUFx3_ASAP7_75t_L g2744 ( 
.A(n_2708),
.Y(n_2744)
);

INVx4_ASAP7_75t_L g2745 ( 
.A(n_2415),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_SL g2746 ( 
.A(n_2336),
.B(n_2029),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2686),
.Y(n_2747)
);

INVx4_ASAP7_75t_L g2748 ( 
.A(n_2415),
.Y(n_2748)
);

AND2x4_ASAP7_75t_L g2749 ( 
.A(n_2734),
.B(n_2738),
.Y(n_2749)
);

INVx1_ASAP7_75t_SL g2750 ( 
.A(n_2511),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2365),
.B(n_2720),
.Y(n_2751)
);

INVx4_ASAP7_75t_L g2752 ( 
.A(n_2415),
.Y(n_2752)
);

INVx1_ASAP7_75t_SL g2753 ( 
.A(n_2563),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2316),
.Y(n_2754)
);

INVx4_ASAP7_75t_L g2755 ( 
.A(n_2415),
.Y(n_2755)
);

INVx4_ASAP7_75t_SL g2756 ( 
.A(n_2493),
.Y(n_2756)
);

AOI22xp33_ASAP7_75t_L g2757 ( 
.A1(n_2455),
.A2(n_2171),
.B1(n_2201),
.B2(n_2173),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2316),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2325),
.B(n_2347),
.Y(n_2759)
);

AOI22xp33_ASAP7_75t_L g2760 ( 
.A1(n_2455),
.A2(n_2171),
.B1(n_2201),
.B2(n_2173),
.Y(n_2760)
);

BUFx2_ASAP7_75t_L g2761 ( 
.A(n_2519),
.Y(n_2761)
);

INVx4_ASAP7_75t_L g2762 ( 
.A(n_2419),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2324),
.Y(n_2763)
);

AND2x4_ASAP7_75t_SL g2764 ( 
.A(n_2385),
.B(n_1646),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2686),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2324),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2472),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2472),
.Y(n_2768)
);

NAND2x1p5_ASAP7_75t_L g2769 ( 
.A(n_2362),
.B(n_2171),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2472),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2354),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2369),
.B(n_2191),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2476),
.Y(n_2773)
);

AND2x4_ASAP7_75t_L g2774 ( 
.A(n_2734),
.B(n_2237),
.Y(n_2774)
);

AND2x4_ASAP7_75t_L g2775 ( 
.A(n_2734),
.B(n_2237),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2476),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2325),
.B(n_1927),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2476),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2354),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2480),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2480),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2355),
.Y(n_2782)
);

OAI221xp5_ASAP7_75t_L g2783 ( 
.A1(n_2588),
.A2(n_2243),
.B1(n_2091),
.B2(n_1752),
.C(n_1812),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2355),
.Y(n_2784)
);

BUFx3_ASAP7_75t_L g2785 ( 
.A(n_2708),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2480),
.Y(n_2786)
);

INVxp67_ASAP7_75t_L g2787 ( 
.A(n_2721),
.Y(n_2787)
);

INVx2_ASAP7_75t_SL g2788 ( 
.A(n_2554),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2489),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2357),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2489),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2489),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2490),
.Y(n_2793)
);

AO21x2_ASAP7_75t_L g2794 ( 
.A1(n_2392),
.A2(n_1972),
.B(n_1971),
.Y(n_2794)
);

BUFx6f_ASAP7_75t_L g2795 ( 
.A(n_2419),
.Y(n_2795)
);

INVxp67_ASAP7_75t_L g2796 ( 
.A(n_2721),
.Y(n_2796)
);

AND2x4_ASAP7_75t_L g2797 ( 
.A(n_2738),
.B(n_2238),
.Y(n_2797)
);

INVx4_ASAP7_75t_L g2798 ( 
.A(n_2419),
.Y(n_2798)
);

NOR2xp33_ASAP7_75t_L g2799 ( 
.A(n_2428),
.B(n_2191),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2490),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2347),
.B(n_2348),
.Y(n_2801)
);

BUFx2_ASAP7_75t_L g2802 ( 
.A(n_2519),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2365),
.B(n_2145),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2490),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2602),
.Y(n_2805)
);

NOR2xp33_ASAP7_75t_L g2806 ( 
.A(n_2384),
.B(n_2175),
.Y(n_2806)
);

AND2x4_ASAP7_75t_L g2807 ( 
.A(n_2738),
.B(n_2238),
.Y(n_2807)
);

BUFx3_ASAP7_75t_L g2808 ( 
.A(n_2598),
.Y(n_2808)
);

AND2x4_ASAP7_75t_L g2809 ( 
.A(n_2598),
.B(n_2238),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2602),
.Y(n_2810)
);

BUFx3_ASAP7_75t_L g2811 ( 
.A(n_2598),
.Y(n_2811)
);

AND2x4_ASAP7_75t_L g2812 ( 
.A(n_2598),
.B(n_2238),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2357),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2361),
.Y(n_2814)
);

INVx4_ASAP7_75t_SL g2815 ( 
.A(n_2493),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2514),
.B(n_2211),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_SL g2817 ( 
.A(n_2336),
.B(n_1972),
.Y(n_2817)
);

OAI21xp5_ASAP7_75t_L g2818 ( 
.A1(n_2395),
.A2(n_2148),
.B(n_1983),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_SL g2819 ( 
.A(n_2336),
.B(n_1979),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2514),
.B(n_2211),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2602),
.Y(n_2821)
);

AO22x2_ASAP7_75t_L g2822 ( 
.A1(n_2701),
.A2(n_1820),
.B1(n_1725),
.B2(n_1810),
.Y(n_2822)
);

INVx2_ASAP7_75t_SL g2823 ( 
.A(n_2554),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2611),
.Y(n_2824)
);

NAND2x1p5_ASAP7_75t_L g2825 ( 
.A(n_2362),
.B(n_2173),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2611),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2611),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2613),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2613),
.Y(n_2829)
);

HB1xp67_ASAP7_75t_L g2830 ( 
.A(n_2332),
.Y(n_2830)
);

AOI22xp33_ASAP7_75t_L g2831 ( 
.A1(n_2455),
.A2(n_2173),
.B1(n_2207),
.B2(n_2201),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2348),
.B(n_1998),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2613),
.Y(n_2833)
);

OAI21xp33_ASAP7_75t_SL g2834 ( 
.A1(n_2406),
.A2(n_1983),
.B(n_1979),
.Y(n_2834)
);

INVx5_ASAP7_75t_L g2835 ( 
.A(n_2486),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2614),
.Y(n_2836)
);

BUFx3_ASAP7_75t_L g2837 ( 
.A(n_2381),
.Y(n_2837)
);

INVx8_ASAP7_75t_L g2838 ( 
.A(n_2486),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2614),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2373),
.B(n_2013),
.Y(n_2840)
);

AOI22xp33_ASAP7_75t_L g2841 ( 
.A1(n_2455),
.A2(n_2201),
.B1(n_2207),
.B2(n_2244),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2614),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2620),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2453),
.B(n_2637),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2363),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2620),
.Y(n_2846)
);

BUFx6f_ASAP7_75t_L g2847 ( 
.A(n_2419),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2620),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2621),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2621),
.Y(n_2850)
);

INVx6_ASAP7_75t_L g2851 ( 
.A(n_2492),
.Y(n_2851)
);

AND2x6_ASAP7_75t_L g2852 ( 
.A(n_2403),
.B(n_1987),
.Y(n_2852)
);

BUFx4_ASAP7_75t_L g2853 ( 
.A(n_2327),
.Y(n_2853)
);

NOR2xp33_ASAP7_75t_L g2854 ( 
.A(n_2384),
.B(n_1538),
.Y(n_2854)
);

AND2x4_ASAP7_75t_L g2855 ( 
.A(n_2425),
.B(n_2244),
.Y(n_2855)
);

BUFx6f_ASAP7_75t_L g2856 ( 
.A(n_2427),
.Y(n_2856)
);

INVxp67_ASAP7_75t_L g2857 ( 
.A(n_2727),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2621),
.Y(n_2858)
);

AOI22xp33_ASAP7_75t_L g2859 ( 
.A1(n_2520),
.A2(n_2601),
.B1(n_2629),
.B2(n_2557),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2368),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2368),
.Y(n_2861)
);

BUFx3_ASAP7_75t_L g2862 ( 
.A(n_2381),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2626),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2370),
.Y(n_2864)
);

AO22x2_ASAP7_75t_L g2865 ( 
.A1(n_2701),
.A2(n_2358),
.B1(n_2454),
.B2(n_2341),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2626),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2373),
.B(n_2042),
.Y(n_2867)
);

CKINVDCx5p33_ASAP7_75t_R g2868 ( 
.A(n_2418),
.Y(n_2868)
);

AND2x2_ASAP7_75t_L g2869 ( 
.A(n_2453),
.B(n_2637),
.Y(n_2869)
);

AND2x6_ASAP7_75t_L g2870 ( 
.A(n_2403),
.B(n_1987),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2626),
.Y(n_2871)
);

INVx3_ASAP7_75t_L g2872 ( 
.A(n_2427),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2628),
.Y(n_2873)
);

NOR2xp33_ASAP7_75t_L g2874 ( 
.A(n_2454),
.B(n_1538),
.Y(n_2874)
);

AND2x4_ASAP7_75t_L g2875 ( 
.A(n_2425),
.B(n_2244),
.Y(n_2875)
);

AND2x2_ASAP7_75t_L g2876 ( 
.A(n_2664),
.B(n_2078),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2628),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2565),
.B(n_2420),
.Y(n_2878)
);

INVxp67_ASAP7_75t_L g2879 ( 
.A(n_2727),
.Y(n_2879)
);

INVx2_ASAP7_75t_L g2880 ( 
.A(n_2370),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2664),
.B(n_2714),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_L g2882 ( 
.A(n_2322),
.B(n_2386),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2407),
.Y(n_2883)
);

AND2x2_ASAP7_75t_L g2884 ( 
.A(n_2714),
.B(n_2078),
.Y(n_2884)
);

BUFx3_ASAP7_75t_L g2885 ( 
.A(n_2381),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2666),
.Y(n_2886)
);

BUFx4f_ASAP7_75t_L g2887 ( 
.A(n_2346),
.Y(n_2887)
);

AND2x4_ASAP7_75t_L g2888 ( 
.A(n_2483),
.B(n_2501),
.Y(n_2888)
);

OR2x2_ASAP7_75t_L g2889 ( 
.A(n_2538),
.B(n_2580),
.Y(n_2889)
);

INVx2_ASAP7_75t_L g2890 ( 
.A(n_2407),
.Y(n_2890)
);

AND3x4_ASAP7_75t_L g2891 ( 
.A(n_2605),
.B(n_1785),
.C(n_1806),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2410),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2444),
.B(n_2080),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2666),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2410),
.Y(n_2895)
);

BUFx2_ASAP7_75t_L g2896 ( 
.A(n_2580),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2667),
.Y(n_2897)
);

NOR2xp33_ASAP7_75t_L g2898 ( 
.A(n_2322),
.B(n_1556),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2422),
.B(n_2256),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_L g2900 ( 
.A(n_2386),
.B(n_1556),
.Y(n_2900)
);

INVx5_ASAP7_75t_L g2901 ( 
.A(n_2486),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2421),
.Y(n_2902)
);

NOR2xp33_ASAP7_75t_L g2903 ( 
.A(n_2401),
.B(n_1560),
.Y(n_2903)
);

NOR2xp33_ASAP7_75t_L g2904 ( 
.A(n_2408),
.B(n_1560),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2667),
.Y(n_2905)
);

AOI22xp33_ASAP7_75t_L g2906 ( 
.A1(n_2520),
.A2(n_2207),
.B1(n_2251),
.B2(n_2244),
.Y(n_2906)
);

INVx4_ASAP7_75t_L g2907 ( 
.A(n_2427),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2667),
.Y(n_2908)
);

NOR2x1p5_ASAP7_75t_L g2909 ( 
.A(n_2327),
.B(n_1676),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2421),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2423),
.Y(n_2911)
);

INVx1_ASAP7_75t_SL g2912 ( 
.A(n_2655),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2672),
.Y(n_2913)
);

INVx4_ASAP7_75t_L g2914 ( 
.A(n_2427),
.Y(n_2914)
);

AND2x6_ASAP7_75t_L g2915 ( 
.A(n_2403),
.B(n_2000),
.Y(n_2915)
);

BUFx6f_ASAP7_75t_L g2916 ( 
.A(n_2427),
.Y(n_2916)
);

INVxp67_ASAP7_75t_L g2917 ( 
.A(n_2533),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2672),
.Y(n_2918)
);

BUFx3_ASAP7_75t_L g2919 ( 
.A(n_2381),
.Y(n_2919)
);

BUFx6f_ASAP7_75t_L g2920 ( 
.A(n_2346),
.Y(n_2920)
);

AND2x2_ASAP7_75t_L g2921 ( 
.A(n_2444),
.B(n_2080),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2672),
.Y(n_2922)
);

BUFx6f_ASAP7_75t_L g2923 ( 
.A(n_2346),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2423),
.Y(n_2924)
);

XNOR2x2_ASAP7_75t_L g2925 ( 
.A(n_2358),
.B(n_898),
.Y(n_2925)
);

INVx2_ASAP7_75t_SL g2926 ( 
.A(n_2556),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2677),
.Y(n_2927)
);

AOI22xp5_ASAP7_75t_L g2928 ( 
.A1(n_2317),
.A2(n_2213),
.B1(n_2036),
.B2(n_2207),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2483),
.B(n_2251),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2380),
.B(n_2251),
.Y(n_2930)
);

CKINVDCx5p33_ASAP7_75t_R g2931 ( 
.A(n_2452),
.Y(n_2931)
);

BUFx6f_ASAP7_75t_L g2932 ( 
.A(n_2346),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2380),
.B(n_2251),
.Y(n_2933)
);

AOI22xp33_ASAP7_75t_L g2934 ( 
.A1(n_2520),
.A2(n_2213),
.B1(n_2002),
.B2(n_2004),
.Y(n_2934)
);

AOI22xp33_ASAP7_75t_L g2935 ( 
.A1(n_2520),
.A2(n_2002),
.B1(n_2004),
.B2(n_2256),
.Y(n_2935)
);

AND2x4_ASAP7_75t_L g2936 ( 
.A(n_2501),
.B(n_2286),
.Y(n_2936)
);

NOR2xp33_ASAP7_75t_L g2937 ( 
.A(n_2566),
.B(n_1676),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2677),
.Y(n_2938)
);

BUFx3_ASAP7_75t_L g2939 ( 
.A(n_2655),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_SL g2940 ( 
.A(n_2377),
.B(n_2000),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2677),
.Y(n_2941)
);

BUFx3_ASAP7_75t_L g2942 ( 
.A(n_2679),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2680),
.Y(n_2943)
);

NOR2xp33_ASAP7_75t_L g2944 ( 
.A(n_2566),
.B(n_1690),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2680),
.Y(n_2945)
);

INVx3_ASAP7_75t_L g2946 ( 
.A(n_2422),
.Y(n_2946)
);

AOI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2317),
.A2(n_2689),
.B1(n_2557),
.B2(n_2629),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2680),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_SL g2949 ( 
.A(n_2377),
.B(n_2310),
.Y(n_2949)
);

NOR2xp33_ASAP7_75t_L g2950 ( 
.A(n_2375),
.B(n_1690),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2432),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2432),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_SL g2953 ( 
.A(n_2466),
.B(n_1589),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2433),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2433),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2443),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2422),
.B(n_2259),
.Y(n_2957)
);

INVx2_ASAP7_75t_SL g2958 ( 
.A(n_2556),
.Y(n_2958)
);

INVx2_ASAP7_75t_SL g2959 ( 
.A(n_2679),
.Y(n_2959)
);

AND2x2_ASAP7_75t_L g2960 ( 
.A(n_2352),
.B(n_2225),
.Y(n_2960)
);

INVx3_ASAP7_75t_L g2961 ( 
.A(n_2422),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2443),
.Y(n_2962)
);

BUFx2_ASAP7_75t_L g2963 ( 
.A(n_2398),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2446),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2446),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2507),
.Y(n_2966)
);

INVx4_ASAP7_75t_L g2967 ( 
.A(n_2486),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2435),
.B(n_1692),
.Y(n_2968)
);

INVx4_ASAP7_75t_L g2969 ( 
.A(n_2486),
.Y(n_2969)
);

INVx3_ASAP7_75t_L g2970 ( 
.A(n_2487),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2507),
.Y(n_2971)
);

BUFx6f_ASAP7_75t_L g2972 ( 
.A(n_2346),
.Y(n_2972)
);

CKINVDCx20_ASAP7_75t_R g2973 ( 
.A(n_2555),
.Y(n_2973)
);

AOI22xp33_ASAP7_75t_L g2974 ( 
.A1(n_2557),
.A2(n_2261),
.B1(n_2268),
.B2(n_2259),
.Y(n_2974)
);

BUFx6f_ASAP7_75t_L g2975 ( 
.A(n_2364),
.Y(n_2975)
);

NAND3xp33_ASAP7_75t_L g2976 ( 
.A(n_2716),
.B(n_1807),
.C(n_1800),
.Y(n_2976)
);

AND2x4_ASAP7_75t_L g2977 ( 
.A(n_2504),
.B(n_2286),
.Y(n_2977)
);

BUFx2_ASAP7_75t_L g2978 ( 
.A(n_2379),
.Y(n_2978)
);

BUFx2_ASAP7_75t_L g2979 ( 
.A(n_2397),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2352),
.B(n_2225),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2509),
.Y(n_2981)
);

AND2x4_ASAP7_75t_L g2982 ( 
.A(n_2504),
.B(n_2286),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2509),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2512),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2512),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2515),
.Y(n_2986)
);

INVx4_ASAP7_75t_L g2987 ( 
.A(n_2526),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2515),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2523),
.Y(n_2989)
);

AND2x4_ASAP7_75t_L g2990 ( 
.A(n_2691),
.B(n_2286),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2523),
.Y(n_2991)
);

AND2x6_ASAP7_75t_L g2992 ( 
.A(n_2431),
.B(n_2304),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2528),
.Y(n_2993)
);

INVx4_ASAP7_75t_L g2994 ( 
.A(n_2526),
.Y(n_2994)
);

AND2x6_ASAP7_75t_L g2995 ( 
.A(n_2431),
.B(n_2304),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2528),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2537),
.Y(n_2997)
);

INVxp67_ASAP7_75t_SL g2998 ( 
.A(n_2487),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2537),
.Y(n_2999)
);

AND2x4_ASAP7_75t_L g3000 ( 
.A(n_2691),
.B(n_2297),
.Y(n_3000)
);

BUFx6f_ASAP7_75t_L g3001 ( 
.A(n_2364),
.Y(n_3001)
);

BUFx6f_ASAP7_75t_L g3002 ( 
.A(n_2364),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2539),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2539),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2487),
.B(n_2261),
.Y(n_3005)
);

BUFx2_ASAP7_75t_L g3006 ( 
.A(n_2474),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2545),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2545),
.Y(n_3008)
);

INVx2_ASAP7_75t_SL g3009 ( 
.A(n_2690),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2548),
.Y(n_3010)
);

AND2x4_ASAP7_75t_L g3011 ( 
.A(n_2691),
.B(n_2715),
.Y(n_3011)
);

NOR2xp33_ASAP7_75t_L g3012 ( 
.A(n_2595),
.B(n_2391),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2548),
.Y(n_3013)
);

AND2x2_ASAP7_75t_L g3014 ( 
.A(n_2356),
.B(n_2303),
.Y(n_3014)
);

BUFx6f_ASAP7_75t_L g3015 ( 
.A(n_2364),
.Y(n_3015)
);

BUFx4f_ASAP7_75t_L g3016 ( 
.A(n_2364),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_2595),
.B(n_1692),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2550),
.Y(n_3018)
);

INVx1_ASAP7_75t_SL g3019 ( 
.A(n_2344),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2550),
.Y(n_3020)
);

AND2x4_ASAP7_75t_L g3021 ( 
.A(n_2691),
.B(n_2297),
.Y(n_3021)
);

AND2x4_ASAP7_75t_L g3022 ( 
.A(n_2715),
.B(n_2297),
.Y(n_3022)
);

OAI221xp5_ASAP7_75t_L g3023 ( 
.A1(n_2694),
.A2(n_1846),
.B1(n_1826),
.B2(n_1801),
.C(n_1096),
.Y(n_3023)
);

BUFx6f_ASAP7_75t_L g3024 ( 
.A(n_2636),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2552),
.Y(n_3025)
);

CKINVDCx20_ASAP7_75t_R g3026 ( 
.A(n_2575),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2552),
.Y(n_3027)
);

NOR2xp33_ASAP7_75t_L g3028 ( 
.A(n_2391),
.B(n_1733),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_2356),
.B(n_2303),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2558),
.Y(n_3030)
);

BUFx6f_ASAP7_75t_L g3031 ( 
.A(n_2636),
.Y(n_3031)
);

INVx3_ASAP7_75t_L g3032 ( 
.A(n_2487),
.Y(n_3032)
);

AND2x6_ASAP7_75t_L g3033 ( 
.A(n_2431),
.B(n_2306),
.Y(n_3033)
);

BUFx10_ASAP7_75t_L g3034 ( 
.A(n_2527),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2558),
.Y(n_3035)
);

BUFx2_ASAP7_75t_L g3036 ( 
.A(n_2351),
.Y(n_3036)
);

AOI22x1_ASAP7_75t_L g3037 ( 
.A1(n_2382),
.A2(n_2310),
.B1(n_2306),
.B2(n_2290),
.Y(n_3037)
);

AND2x2_ASAP7_75t_L g3038 ( 
.A(n_2739),
.B(n_2308),
.Y(n_3038)
);

INVx3_ASAP7_75t_L g3039 ( 
.A(n_2499),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2560),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2560),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2561),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2561),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2567),
.Y(n_3044)
);

NAND2x1p5_ASAP7_75t_L g3045 ( 
.A(n_2362),
.B(n_2167),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_L g3046 ( 
.A(n_2391),
.B(n_1733),
.Y(n_3046)
);

INVx3_ASAP7_75t_L g3047 ( 
.A(n_2499),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2567),
.Y(n_3048)
);

NOR2xp33_ASAP7_75t_L g3049 ( 
.A(n_2391),
.B(n_1751),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2570),
.Y(n_3050)
);

BUFx10_ASAP7_75t_L g3051 ( 
.A(n_2604),
.Y(n_3051)
);

INVx3_ASAP7_75t_L g3052 ( 
.A(n_2499),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2570),
.Y(n_3053)
);

INVx8_ASAP7_75t_L g3054 ( 
.A(n_2526),
.Y(n_3054)
);

CKINVDCx5p33_ASAP7_75t_R g3055 ( 
.A(n_2498),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2571),
.Y(n_3056)
);

AOI22xp33_ASAP7_75t_L g3057 ( 
.A1(n_2557),
.A2(n_2270),
.B1(n_2272),
.B2(n_2268),
.Y(n_3057)
);

BUFx6f_ASAP7_75t_L g3058 ( 
.A(n_2636),
.Y(n_3058)
);

AND2x4_ASAP7_75t_L g3059 ( 
.A(n_2715),
.B(n_2297),
.Y(n_3059)
);

AND2x4_ASAP7_75t_L g3060 ( 
.A(n_2715),
.B(n_2300),
.Y(n_3060)
);

INVx4_ASAP7_75t_SL g3061 ( 
.A(n_2493),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2499),
.B(n_2270),
.Y(n_3062)
);

BUFx6f_ASAP7_75t_L g3063 ( 
.A(n_2636),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2571),
.Y(n_3064)
);

AND2x2_ASAP7_75t_L g3065 ( 
.A(n_2739),
.B(n_2228),
.Y(n_3065)
);

BUFx3_ASAP7_75t_L g3066 ( 
.A(n_2690),
.Y(n_3066)
);

BUFx6f_ASAP7_75t_L g3067 ( 
.A(n_2636),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2579),
.Y(n_3068)
);

NOR2xp33_ASAP7_75t_L g3069 ( 
.A(n_2479),
.B(n_1751),
.Y(n_3069)
);

OR2x6_ASAP7_75t_L g3070 ( 
.A(n_2526),
.B(n_2300),
.Y(n_3070)
);

NOR2xp33_ASAP7_75t_L g3071 ( 
.A(n_2479),
.B(n_1770),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2579),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2581),
.Y(n_3073)
);

BUFx3_ASAP7_75t_L g3074 ( 
.A(n_2492),
.Y(n_3074)
);

INVxp67_ASAP7_75t_SL g3075 ( 
.A(n_2510),
.Y(n_3075)
);

INVx3_ASAP7_75t_L g3076 ( 
.A(n_2510),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2581),
.Y(n_3077)
);

AND2x4_ASAP7_75t_L g3078 ( 
.A(n_2717),
.B(n_2300),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2593),
.Y(n_3079)
);

BUFx3_ASAP7_75t_L g3080 ( 
.A(n_2492),
.Y(n_3080)
);

NOR2xp33_ASAP7_75t_L g3081 ( 
.A(n_2479),
.B(n_2600),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2593),
.Y(n_3082)
);

CKINVDCx20_ASAP7_75t_R g3083 ( 
.A(n_2569),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2594),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2594),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2633),
.Y(n_3086)
);

NOR2xp33_ASAP7_75t_L g3087 ( 
.A(n_2479),
.B(n_1770),
.Y(n_3087)
);

AND2x2_ASAP7_75t_L g3088 ( 
.A(n_2328),
.B(n_2308),
.Y(n_3088)
);

INVx8_ASAP7_75t_L g3089 ( 
.A(n_2526),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2510),
.B(n_2722),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2635),
.Y(n_3091)
);

OAI22xp5_ASAP7_75t_L g3092 ( 
.A1(n_2463),
.A2(n_2044),
.B1(n_2273),
.B2(n_2272),
.Y(n_3092)
);

INVx4_ASAP7_75t_L g3093 ( 
.A(n_2459),
.Y(n_3093)
);

BUFx6f_ASAP7_75t_L g3094 ( 
.A(n_2639),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2643),
.Y(n_3095)
);

INVx2_ASAP7_75t_SL g3096 ( 
.A(n_2689),
.Y(n_3096)
);

AOI22xp33_ASAP7_75t_L g3097 ( 
.A1(n_2601),
.A2(n_2274),
.B1(n_2276),
.B2(n_2273),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2645),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2645),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_2646),
.Y(n_3100)
);

INVx4_ASAP7_75t_SL g3101 ( 
.A(n_2493),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_SL g3102 ( 
.A(n_2638),
.B(n_1632),
.Y(n_3102)
);

INVxp67_ASAP7_75t_L g3103 ( 
.A(n_2617),
.Y(n_3103)
);

NAND2x1p5_ASAP7_75t_L g3104 ( 
.A(n_2366),
.B(n_2167),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2646),
.Y(n_3105)
);

BUFx8_ASAP7_75t_SL g3106 ( 
.A(n_2651),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_SL g3107 ( 
.A(n_2377),
.B(n_2285),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_SL g3108 ( 
.A(n_2323),
.B(n_2285),
.Y(n_3108)
);

OAI221xp5_ASAP7_75t_L g3109 ( 
.A1(n_2541),
.A2(n_1096),
.B1(n_1099),
.B2(n_1039),
.C(n_1431),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2656),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2656),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2551),
.B(n_2276),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2659),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_2659),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_2328),
.B(n_2228),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2681),
.B(n_2257),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2688),
.Y(n_3117)
);

NAND3xp33_ASAP7_75t_L g3118 ( 
.A(n_2592),
.B(n_1807),
.C(n_1800),
.Y(n_3118)
);

INVx4_ASAP7_75t_L g3119 ( 
.A(n_2459),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_L g3120 ( 
.A(n_2541),
.B(n_1787),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2688),
.Y(n_3121)
);

AND2x4_ASAP7_75t_L g3122 ( 
.A(n_2717),
.B(n_2300),
.Y(n_3122)
);

CKINVDCx5p33_ASAP7_75t_R g3123 ( 
.A(n_2409),
.Y(n_3123)
);

AND2x4_ASAP7_75t_L g3124 ( 
.A(n_2717),
.B(n_2229),
.Y(n_3124)
);

INVx4_ASAP7_75t_L g3125 ( 
.A(n_2459),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2692),
.Y(n_3126)
);

BUFx2_ASAP7_75t_L g3127 ( 
.A(n_2385),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2693),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2693),
.Y(n_3129)
);

INVx4_ASAP7_75t_L g3130 ( 
.A(n_2459),
.Y(n_3130)
);

AND2x2_ASAP7_75t_SL g3131 ( 
.A(n_2689),
.B(n_826),
.Y(n_3131)
);

BUFx4f_ASAP7_75t_L g3132 ( 
.A(n_2459),
.Y(n_3132)
);

NOR2xp33_ASAP7_75t_L g3133 ( 
.A(n_2339),
.B(n_1787),
.Y(n_3133)
);

BUFx3_ASAP7_75t_L g3134 ( 
.A(n_2717),
.Y(n_3134)
);

AO22x2_ASAP7_75t_L g3135 ( 
.A1(n_2450),
.A2(n_1820),
.B1(n_1806),
.B2(n_1810),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2695),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2333),
.B(n_2266),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2695),
.Y(n_3138)
);

AND2x2_ASAP7_75t_L g3139 ( 
.A(n_2333),
.B(n_2229),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2699),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2337),
.B(n_2236),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2699),
.Y(n_3142)
);

INVx1_ASAP7_75t_SL g3143 ( 
.A(n_2564),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2702),
.Y(n_3144)
);

NOR2xp33_ASAP7_75t_L g3145 ( 
.A(n_2339),
.B(n_1642),
.Y(n_3145)
);

NOR2xp33_ASAP7_75t_L g3146 ( 
.A(n_2339),
.B(n_2277),
.Y(n_3146)
);

CKINVDCx5p33_ASAP7_75t_R g3147 ( 
.A(n_2582),
.Y(n_3147)
);

AND2x2_ASAP7_75t_SL g3148 ( 
.A(n_2343),
.B(n_826),
.Y(n_3148)
);

OR2x2_ASAP7_75t_L g3149 ( 
.A(n_2568),
.B(n_1331),
.Y(n_3149)
);

BUFx3_ASAP7_75t_L g3150 ( 
.A(n_2385),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_SL g3151 ( 
.A(n_2323),
.B(n_2290),
.Y(n_3151)
);

OAI22xp5_ASAP7_75t_L g3152 ( 
.A1(n_2436),
.A2(n_2461),
.B1(n_2438),
.B2(n_2366),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2702),
.Y(n_3153)
);

AND2x4_ASAP7_75t_L g3154 ( 
.A(n_2601),
.B(n_2236),
.Y(n_3154)
);

AND2x2_ASAP7_75t_L g3155 ( 
.A(n_2349),
.B(n_2252),
.Y(n_3155)
);

AND2x2_ASAP7_75t_L g3156 ( 
.A(n_2349),
.B(n_2252),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2724),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2728),
.Y(n_3158)
);

OR2x6_ASAP7_75t_L g3159 ( 
.A(n_2385),
.B(n_2275),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2728),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2731),
.Y(n_3161)
);

NOR2xp33_ASAP7_75t_SL g3162 ( 
.A(n_2713),
.B(n_1659),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_L g3163 ( 
.A(n_2339),
.B(n_2289),
.Y(n_3163)
);

BUFx6f_ASAP7_75t_L g3164 ( 
.A(n_2639),
.Y(n_3164)
);

NOR3xp33_ASAP7_75t_L g3165 ( 
.A(n_2378),
.B(n_2275),
.C(n_1481),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2731),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2601),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2629),
.Y(n_3168)
);

NOR2xp33_ASAP7_75t_L g3169 ( 
.A(n_2484),
.B(n_2578),
.Y(n_3169)
);

OAI22xp5_ASAP7_75t_L g3170 ( 
.A1(n_2436),
.A2(n_2294),
.B1(n_2296),
.B2(n_2291),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_2630),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2629),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2658),
.Y(n_3173)
);

INVx6_ASAP7_75t_L g3174 ( 
.A(n_2587),
.Y(n_3174)
);

AND2x4_ASAP7_75t_L g3175 ( 
.A(n_2658),
.B(n_2186),
.Y(n_3175)
);

NOR2xp33_ASAP7_75t_L g3176 ( 
.A(n_2707),
.B(n_2299),
.Y(n_3176)
);

INVx2_ASAP7_75t_SL g3177 ( 
.A(n_2658),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2353),
.B(n_2305),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_3176),
.B(n_2353),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2771),
.Y(n_3180)
);

OAI22xp5_ASAP7_75t_L g3181 ( 
.A1(n_3090),
.A2(n_2438),
.B1(n_2461),
.B2(n_2436),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_3176),
.B(n_2360),
.Y(n_3182)
);

NOR2xp33_ASAP7_75t_L g3183 ( 
.A(n_2917),
.B(n_2447),
.Y(n_3183)
);

NOR2xp67_ASAP7_75t_L g3184 ( 
.A(n_2931),
.B(n_2726),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_3112),
.B(n_2360),
.Y(n_3185)
);

INVx2_ASAP7_75t_SL g3186 ( 
.A(n_2939),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_SL g3187 ( 
.A(n_3132),
.B(n_2508),
.Y(n_3187)
);

OR2x2_ASAP7_75t_L g3188 ( 
.A(n_2889),
.B(n_2597),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2960),
.B(n_2371),
.Y(n_3189)
);

AND2x4_ASAP7_75t_SL g3190 ( 
.A(n_3034),
.B(n_2569),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2771),
.Y(n_3191)
);

O2A1O1Ixp5_ASAP7_75t_L g3192 ( 
.A1(n_2817),
.A2(n_2465),
.B(n_2326),
.C(n_2434),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_2772),
.B(n_2599),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_SL g3194 ( 
.A(n_2751),
.B(n_2508),
.Y(n_3194)
);

INVx3_ASAP7_75t_L g3195 ( 
.A(n_2745),
.Y(n_3195)
);

NOR2xp33_ASAP7_75t_L g3196 ( 
.A(n_2772),
.B(n_2682),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2960),
.B(n_2371),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2980),
.B(n_2383),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_2980),
.B(n_2383),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_SL g3200 ( 
.A(n_2749),
.B(n_2508),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2946),
.A2(n_2687),
.B(n_2553),
.Y(n_3201)
);

AOI22xp33_ASAP7_75t_L g3202 ( 
.A1(n_2925),
.A2(n_2518),
.B1(n_2719),
.B2(n_2522),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_3014),
.B(n_2387),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2779),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_SL g3205 ( 
.A(n_2749),
.B(n_2508),
.Y(n_3205)
);

NOR2xp33_ASAP7_75t_L g3206 ( 
.A(n_2799),
.B(n_2586),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_3014),
.B(n_2387),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_3029),
.B(n_2389),
.Y(n_3208)
);

INVx4_ASAP7_75t_L g3209 ( 
.A(n_2741),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_3029),
.B(n_2389),
.Y(n_3210)
);

NOR2xp33_ASAP7_75t_L g3211 ( 
.A(n_2799),
.B(n_2488),
.Y(n_3211)
);

NOR2xp33_ASAP7_75t_L g3212 ( 
.A(n_2787),
.B(n_2495),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_2747),
.Y(n_3213)
);

AND2x4_ASAP7_75t_L g3214 ( 
.A(n_2808),
.B(n_2587),
.Y(n_3214)
);

AOI22xp33_ASAP7_75t_L g3215 ( 
.A1(n_2925),
.A2(n_2518),
.B1(n_2522),
.B2(n_2658),
.Y(n_3215)
);

OAI22xp33_ASAP7_75t_SL g3216 ( 
.A1(n_3109),
.A2(n_2624),
.B1(n_2503),
.B2(n_2485),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_SL g3217 ( 
.A(n_3132),
.B(n_2544),
.Y(n_3217)
);

AOI22xp33_ASAP7_75t_L g3218 ( 
.A1(n_2865),
.A2(n_2518),
.B1(n_2673),
.B2(n_2670),
.Y(n_3218)
);

NOR2xp33_ASAP7_75t_L g3219 ( 
.A(n_2796),
.B(n_2516),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_2747),
.Y(n_3220)
);

INVxp67_ASAP7_75t_L g3221 ( 
.A(n_2978),
.Y(n_3221)
);

INVxp67_ASAP7_75t_L g3222 ( 
.A(n_2979),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2893),
.B(n_2394),
.Y(n_3223)
);

INVxp67_ASAP7_75t_SL g3224 ( 
.A(n_2741),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2893),
.B(n_2394),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2921),
.B(n_2803),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_2782),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_2921),
.B(n_2399),
.Y(n_3228)
);

AOI22xp33_ASAP7_75t_L g3229 ( 
.A1(n_2865),
.A2(n_2673),
.B1(n_2670),
.B2(n_2402),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2803),
.B(n_2399),
.Y(n_3230)
);

BUFx8_ASAP7_75t_L g3231 ( 
.A(n_3006),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_3038),
.B(n_2402),
.Y(n_3232)
);

OAI22xp5_ASAP7_75t_L g3233 ( 
.A1(n_2859),
.A2(n_2461),
.B1(n_2438),
.B2(n_2544),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_3038),
.B(n_2404),
.Y(n_3234)
);

OAI22xp5_ASAP7_75t_L g3235 ( 
.A1(n_2998),
.A2(n_2544),
.B1(n_2366),
.B2(n_2393),
.Y(n_3235)
);

AOI22xp33_ASAP7_75t_L g3236 ( 
.A1(n_2865),
.A2(n_2673),
.B1(n_2670),
.B2(n_2411),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_3065),
.B(n_2404),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_3065),
.B(n_2411),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2765),
.Y(n_3239)
);

NAND2xp33_ASAP7_75t_L g3240 ( 
.A(n_2835),
.B(n_2544),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_3088),
.B(n_3115),
.Y(n_3241)
);

NOR2xp33_ASAP7_75t_L g3242 ( 
.A(n_2857),
.B(n_2647),
.Y(n_3242)
);

INVx2_ASAP7_75t_L g3243 ( 
.A(n_2784),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_2844),
.B(n_2660),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2784),
.Y(n_3245)
);

NAND2x1p5_ASAP7_75t_L g3246 ( 
.A(n_3132),
.B(n_2372),
.Y(n_3246)
);

NOR2xp33_ASAP7_75t_L g3247 ( 
.A(n_2879),
.B(n_2668),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_3088),
.B(n_2412),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2790),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_3115),
.B(n_2412),
.Y(n_3250)
);

AOI22xp33_ASAP7_75t_L g3251 ( 
.A1(n_3148),
.A2(n_2673),
.B1(n_2670),
.B2(n_2437),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3139),
.B(n_2430),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3139),
.B(n_2430),
.Y(n_3253)
);

AOI22xp5_ASAP7_75t_L g3254 ( 
.A1(n_2950),
.A2(n_2697),
.B1(n_2723),
.B2(n_2674),
.Y(n_3254)
);

INVx2_ASAP7_75t_L g3255 ( 
.A(n_2813),
.Y(n_3255)
);

NOR2xp33_ASAP7_75t_L g3256 ( 
.A(n_3012),
.B(n_2559),
.Y(n_3256)
);

AOI22xp5_ASAP7_75t_L g3257 ( 
.A1(n_2950),
.A2(n_2549),
.B1(n_2477),
.B2(n_2618),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_SL g3258 ( 
.A(n_2749),
.B(n_2774),
.Y(n_3258)
);

AOI22xp33_ASAP7_75t_L g3259 ( 
.A1(n_3148),
.A2(n_2441),
.B1(n_2448),
.B2(n_2437),
.Y(n_3259)
);

OR2x2_ASAP7_75t_L g3260 ( 
.A(n_2750),
.B(n_2711),
.Y(n_3260)
);

BUFx2_ASAP7_75t_L g3261 ( 
.A(n_2761),
.Y(n_3261)
);

NAND3xp33_ASAP7_75t_L g3262 ( 
.A(n_2874),
.B(n_1617),
.C(n_1598),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3141),
.B(n_2441),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_SL g3264 ( 
.A(n_2774),
.B(n_2544),
.Y(n_3264)
);

AOI22xp5_ASAP7_75t_L g3265 ( 
.A1(n_2968),
.A2(n_2676),
.B1(n_2705),
.B2(n_2698),
.Y(n_3265)
);

NOR2xp33_ASAP7_75t_L g3266 ( 
.A(n_3012),
.B(n_2350),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3141),
.B(n_2448),
.Y(n_3267)
);

NOR2xp33_ASAP7_75t_L g3268 ( 
.A(n_2874),
.B(n_2359),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_3155),
.B(n_3156),
.Y(n_3269)
);

BUFx2_ASAP7_75t_L g3270 ( 
.A(n_2802),
.Y(n_3270)
);

OAI22x1_ASAP7_75t_R g3271 ( 
.A1(n_2740),
.A2(n_1687),
.B1(n_1707),
.B2(n_1607),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_SL g3272 ( 
.A(n_2774),
.B(n_2323),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_SL g3273 ( 
.A(n_2775),
.B(n_2323),
.Y(n_3273)
);

INVx3_ASAP7_75t_L g3274 ( 
.A(n_2745),
.Y(n_3274)
);

AOI22xp33_ASAP7_75t_L g3275 ( 
.A1(n_3131),
.A2(n_2460),
.B1(n_2464),
.B2(n_2457),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_SL g3276 ( 
.A(n_2946),
.B(n_2323),
.Y(n_3276)
);

A2O1A1Ixp33_ASAP7_75t_SL g3277 ( 
.A1(n_3146),
.A2(n_2460),
.B(n_2464),
.C(n_2457),
.Y(n_3277)
);

BUFx8_ASAP7_75t_L g3278 ( 
.A(n_2896),
.Y(n_3278)
);

NOR2xp33_ASAP7_75t_SL g3279 ( 
.A(n_2953),
.B(n_2729),
.Y(n_3279)
);

AOI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_2946),
.A2(n_2687),
.B(n_2553),
.Y(n_3280)
);

OAI22xp5_ASAP7_75t_L g3281 ( 
.A1(n_3075),
.A2(n_2372),
.B1(n_2393),
.B2(n_2524),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2814),
.Y(n_3282)
);

OAI22xp33_ASAP7_75t_L g3283 ( 
.A1(n_2968),
.A2(n_2468),
.B1(n_2470),
.B2(n_2469),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2814),
.Y(n_3284)
);

NAND2xp33_ASAP7_75t_L g3285 ( 
.A(n_2835),
.B(n_2323),
.Y(n_3285)
);

HB1xp67_ASAP7_75t_L g3286 ( 
.A(n_2744),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3155),
.B(n_2468),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3156),
.B(n_2469),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2845),
.Y(n_3289)
);

NOR2xp33_ASAP7_75t_L g3290 ( 
.A(n_2854),
.B(n_2726),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2860),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_SL g3292 ( 
.A(n_2775),
.B(n_2553),
.Y(n_3292)
);

AOI22xp33_ASAP7_75t_L g3293 ( 
.A1(n_3131),
.A2(n_2473),
.B1(n_2482),
.B2(n_2470),
.Y(n_3293)
);

HB1xp67_ASAP7_75t_L g3294 ( 
.A(n_2785),
.Y(n_3294)
);

INVx4_ASAP7_75t_L g3295 ( 
.A(n_2741),
.Y(n_3295)
);

AND2x2_ASAP7_75t_L g3296 ( 
.A(n_2869),
.B(n_1534),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_2876),
.B(n_2884),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_2860),
.Y(n_3298)
);

INVxp67_ASAP7_75t_L g3299 ( 
.A(n_2830),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_SL g3300 ( 
.A(n_2775),
.B(n_2553),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_2876),
.B(n_2473),
.Y(n_3301)
);

AOI22xp33_ASAP7_75t_L g3302 ( 
.A1(n_2930),
.A2(n_2491),
.B1(n_2494),
.B2(n_2482),
.Y(n_3302)
);

INVx3_ASAP7_75t_L g3303 ( 
.A(n_2745),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_2797),
.B(n_2687),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_L g3305 ( 
.A(n_2884),
.B(n_2491),
.Y(n_3305)
);

NOR2xp33_ASAP7_75t_L g3306 ( 
.A(n_2854),
.B(n_2704),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_2881),
.B(n_2494),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_2898),
.B(n_2900),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_2881),
.B(n_2496),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_2816),
.B(n_2496),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_2861),
.Y(n_3311)
);

BUFx4_ASAP7_75t_L g3312 ( 
.A(n_2853),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2861),
.Y(n_3313)
);

AOI22xp5_ASAP7_75t_L g3314 ( 
.A1(n_3169),
.A2(n_2706),
.B1(n_2583),
.B2(n_2606),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_2864),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_SL g3316 ( 
.A(n_2961),
.B(n_2687),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_2816),
.B(n_2497),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_2864),
.Y(n_3318)
);

AOI22xp33_ASAP7_75t_L g3319 ( 
.A1(n_2930),
.A2(n_2497),
.B1(n_2521),
.B2(n_2513),
.Y(n_3319)
);

BUFx5_ASAP7_75t_L g3320 ( 
.A(n_2852),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_SL g3321 ( 
.A(n_2961),
.B(n_2696),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_2820),
.B(n_2513),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_SL g3323 ( 
.A(n_2961),
.B(n_2696),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_2820),
.B(n_2521),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_2880),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_SL g3326 ( 
.A(n_2970),
.B(n_2696),
.Y(n_3326)
);

BUFx3_ASAP7_75t_L g3327 ( 
.A(n_2963),
.Y(n_3327)
);

NAND3xp33_ASAP7_75t_L g3328 ( 
.A(n_2900),
.B(n_1706),
.C(n_1617),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_2933),
.B(n_2788),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_2933),
.B(n_2529),
.Y(n_3330)
);

BUFx4f_ASAP7_75t_L g3331 ( 
.A(n_2851),
.Y(n_3331)
);

AOI22xp33_ASAP7_75t_L g3332 ( 
.A1(n_2788),
.A2(n_2529),
.B1(n_2534),
.B2(n_2531),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2823),
.B(n_2531),
.Y(n_3333)
);

AOI21x1_ASAP7_75t_L g3334 ( 
.A1(n_2949),
.A2(n_2732),
.B(n_2630),
.Y(n_3334)
);

AND2x2_ASAP7_75t_L g3335 ( 
.A(n_2753),
.B(n_2502),
.Y(n_3335)
);

O2A1O1Ixp33_ASAP7_75t_L g3336 ( 
.A1(n_3103),
.A2(n_2619),
.B(n_2314),
.C(n_2506),
.Y(n_3336)
);

OAI22xp33_ASAP7_75t_L g3337 ( 
.A1(n_2867),
.A2(n_2536),
.B1(n_2540),
.B2(n_2535),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_2926),
.B(n_2535),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_2880),
.Y(n_3339)
);

INVx4_ASAP7_75t_L g3340 ( 
.A(n_2741),
.Y(n_3340)
);

AOI22x1_ASAP7_75t_L g3341 ( 
.A1(n_2883),
.A2(n_2540),
.B1(n_2543),
.B2(n_2536),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_2926),
.B(n_2543),
.Y(n_3342)
);

NOR2xp67_ASAP7_75t_SL g3343 ( 
.A(n_2835),
.B(n_2372),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_SL g3344 ( 
.A(n_2970),
.B(n_2696),
.Y(n_3344)
);

HB1xp67_ASAP7_75t_L g3345 ( 
.A(n_2912),
.Y(n_3345)
);

AOI22xp5_ASAP7_75t_L g3346 ( 
.A1(n_3169),
.A2(n_2650),
.B1(n_2725),
.B2(n_2609),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_2958),
.B(n_2546),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_2959),
.B(n_2546),
.Y(n_3348)
);

O2A1O1Ixp5_ASAP7_75t_L g3349 ( 
.A1(n_2817),
.A2(n_2562),
.B(n_2573),
.C(n_2547),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_3009),
.B(n_2547),
.Y(n_3350)
);

OAI22xp33_ASAP7_75t_L g3351 ( 
.A1(n_2759),
.A2(n_2573),
.B1(n_2577),
.B2(n_2562),
.Y(n_3351)
);

NAND2xp33_ASAP7_75t_L g3352 ( 
.A(n_2835),
.B(n_2736),
.Y(n_3352)
);

O2A1O1Ixp5_ASAP7_75t_L g3353 ( 
.A1(n_2819),
.A2(n_2584),
.B(n_2590),
.C(n_2577),
.Y(n_3353)
);

AOI22xp5_ASAP7_75t_L g3354 ( 
.A1(n_3081),
.A2(n_2737),
.B1(n_2584),
.B2(n_2596),
.Y(n_3354)
);

AOI21xp5_ASAP7_75t_L g3355 ( 
.A1(n_2970),
.A2(n_2426),
.B(n_2424),
.Y(n_3355)
);

NAND3xp33_ASAP7_75t_L g3356 ( 
.A(n_2903),
.B(n_1706),
.C(n_1617),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_SL g3357 ( 
.A(n_3032),
.B(n_2393),
.Y(n_3357)
);

CKINVDCx5p33_ASAP7_75t_R g3358 ( 
.A(n_2868),
.Y(n_3358)
);

AND2x2_ASAP7_75t_L g3359 ( 
.A(n_2882),
.B(n_2574),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_2890),
.Y(n_3360)
);

NOR2xp33_ASAP7_75t_L g3361 ( 
.A(n_2806),
.B(n_2709),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_SL g3362 ( 
.A(n_3032),
.B(n_2625),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_2890),
.Y(n_3363)
);

NOR2xp33_ASAP7_75t_L g3364 ( 
.A(n_2806),
.B(n_2709),
.Y(n_3364)
);

OAI22xp33_ASAP7_75t_L g3365 ( 
.A1(n_2801),
.A2(n_2596),
.B1(n_2603),
.B2(n_2590),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_SL g3366 ( 
.A(n_3032),
.B(n_2625),
.Y(n_3366)
);

NOR2xp33_ASAP7_75t_L g3367 ( 
.A(n_3149),
.B(n_2730),
.Y(n_3367)
);

INVx2_ASAP7_75t_L g3368 ( 
.A(n_2892),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_SL g3369 ( 
.A(n_3039),
.B(n_2625),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_SL g3370 ( 
.A(n_3039),
.B(n_2625),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_SL g3371 ( 
.A(n_3039),
.B(n_2603),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_2895),
.Y(n_3372)
);

AOI22xp5_ASAP7_75t_L g3373 ( 
.A1(n_3081),
.A2(n_2737),
.B1(n_2730),
.B2(n_2615),
.Y(n_3373)
);

INVx2_ASAP7_75t_SL g3374 ( 
.A(n_3036),
.Y(n_3374)
);

AND2x4_ASAP7_75t_L g3375 ( 
.A(n_2808),
.B(n_2439),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3009),
.B(n_2610),
.Y(n_3376)
);

INVx2_ASAP7_75t_L g3377 ( 
.A(n_2895),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_2902),
.Y(n_3378)
);

AOI22xp33_ASAP7_75t_L g3379 ( 
.A1(n_2902),
.A2(n_2911),
.B1(n_2924),
.B2(n_2910),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_2777),
.B(n_2610),
.Y(n_3380)
);

NAND3xp33_ASAP7_75t_L g3381 ( 
.A(n_2903),
.B(n_1734),
.C(n_1706),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_2910),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2911),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3146),
.B(n_2615),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3163),
.B(n_2627),
.Y(n_3385)
);

AOI22xp33_ASAP7_75t_L g3386 ( 
.A1(n_2951),
.A2(n_2632),
.B1(n_2634),
.B2(n_2627),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2951),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_2952),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3163),
.B(n_2632),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_2878),
.B(n_2634),
.Y(n_3390)
);

AOI22xp33_ASAP7_75t_SL g3391 ( 
.A1(n_2937),
.A2(n_2525),
.B1(n_1800),
.B2(n_1901),
.Y(n_3391)
);

BUFx3_ASAP7_75t_L g3392 ( 
.A(n_3034),
.Y(n_3392)
);

AOI21xp5_ASAP7_75t_L g3393 ( 
.A1(n_3047),
.A2(n_2451),
.B(n_2429),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_SL g3394 ( 
.A(n_2797),
.B(n_2704),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_2952),
.Y(n_3395)
);

NOR2xp33_ASAP7_75t_L g3396 ( 
.A(n_3051),
.B(n_2710),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_2888),
.B(n_2640),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_2888),
.B(n_2640),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_2954),
.Y(n_3399)
);

OR2x2_ASAP7_75t_L g3400 ( 
.A(n_3019),
.B(n_2644),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_2955),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_SL g3402 ( 
.A(n_2797),
.B(n_2710),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_2955),
.Y(n_3403)
);

NOR2xp33_ASAP7_75t_L g3404 ( 
.A(n_3051),
.B(n_2644),
.Y(n_3404)
);

BUFx6f_ASAP7_75t_L g3405 ( 
.A(n_2795),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_2888),
.B(n_2648),
.Y(n_3406)
);

BUFx6f_ASAP7_75t_L g3407 ( 
.A(n_2795),
.Y(n_3407)
);

NOR2xp33_ASAP7_75t_L g3408 ( 
.A(n_3051),
.B(n_2648),
.Y(n_3408)
);

NOR2xp33_ASAP7_75t_L g3409 ( 
.A(n_2942),
.B(n_2652),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_2832),
.B(n_2652),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_2840),
.B(n_2653),
.Y(n_3411)
);

NAND2x1p5_ASAP7_75t_L g3412 ( 
.A(n_3093),
.B(n_2524),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3116),
.B(n_2653),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_2956),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_L g3415 ( 
.A(n_2942),
.B(n_2654),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_L g3416 ( 
.A(n_3066),
.B(n_2654),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_2985),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_SL g3418 ( 
.A(n_2807),
.B(n_2657),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_SL g3419 ( 
.A(n_3047),
.B(n_2661),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3137),
.B(n_2661),
.Y(n_3420)
);

INVx4_ASAP7_75t_L g3421 ( 
.A(n_2795),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_3178),
.B(n_2662),
.Y(n_3422)
);

INVx2_ASAP7_75t_SL g3423 ( 
.A(n_3034),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_2985),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_SL g3425 ( 
.A(n_3047),
.B(n_2662),
.Y(n_3425)
);

INVxp33_ASAP7_75t_L g3426 ( 
.A(n_2904),
.Y(n_3426)
);

NOR2xp33_ASAP7_75t_L g3427 ( 
.A(n_3143),
.B(n_2700),
.Y(n_3427)
);

NOR2xp33_ASAP7_75t_L g3428 ( 
.A(n_3123),
.B(n_2700),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_SL g3429 ( 
.A(n_3052),
.B(n_2663),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3124),
.B(n_2669),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_2986),
.Y(n_3431)
);

INVx3_ASAP7_75t_L g3432 ( 
.A(n_2748),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3124),
.B(n_2669),
.Y(n_3433)
);

NAND2x1p5_ASAP7_75t_L g3434 ( 
.A(n_3093),
.B(n_2524),
.Y(n_3434)
);

INVx5_ASAP7_75t_L g3435 ( 
.A(n_2795),
.Y(n_3435)
);

AND2x6_ASAP7_75t_SL g3436 ( 
.A(n_3120),
.B(n_2439),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_2986),
.Y(n_3437)
);

O2A1O1Ixp33_ASAP7_75t_L g3438 ( 
.A1(n_2783),
.A2(n_2619),
.B(n_2314),
.C(n_2506),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_3124),
.B(n_2671),
.Y(n_3439)
);

NOR2xp33_ASAP7_75t_L g3440 ( 
.A(n_3123),
.B(n_2712),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3154),
.B(n_2671),
.Y(n_3441)
);

A2O1A1Ixp33_ASAP7_75t_L g3442 ( 
.A1(n_2904),
.A2(n_2712),
.B(n_2458),
.C(n_2641),
.Y(n_3442)
);

AND2x2_ASAP7_75t_SL g3443 ( 
.A(n_2937),
.B(n_2517),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_SL g3444 ( 
.A(n_2807),
.B(n_2809),
.Y(n_3444)
);

NOR2xp33_ASAP7_75t_L g3445 ( 
.A(n_3017),
.B(n_1866),
.Y(n_3445)
);

HB1xp67_ASAP7_75t_L g3446 ( 
.A(n_2837),
.Y(n_3446)
);

AOI22xp5_ASAP7_75t_L g3447 ( 
.A1(n_2944),
.A2(n_2525),
.B1(n_2622),
.B2(n_2616),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3154),
.B(n_2345),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3154),
.B(n_2345),
.Y(n_3449)
);

AOI22xp33_ASAP7_75t_L g3450 ( 
.A1(n_2989),
.A2(n_2493),
.B1(n_2631),
.B2(n_2608),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_2989),
.Y(n_3451)
);

CKINVDCx5p33_ASAP7_75t_R g3452 ( 
.A(n_2868),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_2855),
.B(n_2345),
.Y(n_3453)
);

AOI22xp33_ASAP7_75t_L g3454 ( 
.A1(n_2999),
.A2(n_2493),
.B1(n_2631),
.B2(n_2608),
.Y(n_3454)
);

NOR2xp33_ASAP7_75t_L g3455 ( 
.A(n_3145),
.B(n_1866),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_2999),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_2855),
.B(n_2345),
.Y(n_3457)
);

AOI22xp5_ASAP7_75t_L g3458 ( 
.A1(n_2944),
.A2(n_2525),
.B1(n_2649),
.B2(n_2608),
.Y(n_3458)
);

NAND2x1p5_ASAP7_75t_L g3459 ( 
.A(n_3093),
.B(n_2591),
.Y(n_3459)
);

NOR2xp33_ASAP7_75t_L g3460 ( 
.A(n_3145),
.B(n_2099),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3040),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_2855),
.B(n_2623),
.Y(n_3462)
);

AOI22xp33_ASAP7_75t_L g3463 ( 
.A1(n_3040),
.A2(n_2493),
.B1(n_2631),
.B2(n_2608),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_2875),
.B(n_2623),
.Y(n_3464)
);

AOI22xp33_ASAP7_75t_L g3465 ( 
.A1(n_3041),
.A2(n_2608),
.B1(n_2703),
.B2(n_2631),
.Y(n_3465)
);

AND2x2_ASAP7_75t_L g3466 ( 
.A(n_3165),
.B(n_2439),
.Y(n_3466)
);

NOR2xp33_ASAP7_75t_L g3467 ( 
.A(n_2837),
.B(n_2099),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3041),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3043),
.Y(n_3469)
);

OR2x2_ASAP7_75t_L g3470 ( 
.A(n_3159),
.B(n_1975),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_2875),
.B(n_2675),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_2929),
.B(n_2678),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3043),
.Y(n_3473)
);

NOR2xp33_ASAP7_75t_L g3474 ( 
.A(n_2862),
.B(n_2439),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_2929),
.B(n_2703),
.Y(n_3475)
);

O2A1O1Ixp33_ASAP7_75t_L g3476 ( 
.A1(n_3023),
.A2(n_1074),
.B(n_2718),
.C(n_2685),
.Y(n_3476)
);

INVx2_ASAP7_75t_SL g3477 ( 
.A(n_3174),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3072),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_3028),
.B(n_2439),
.Y(n_3479)
);

BUFx3_ASAP7_75t_L g3480 ( 
.A(n_2973),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_L g3481 ( 
.A(n_2862),
.B(n_2485),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3084),
.Y(n_3482)
);

NOR2xp33_ASAP7_75t_L g3483 ( 
.A(n_2885),
.B(n_2485),
.Y(n_3483)
);

INVx3_ASAP7_75t_L g3484 ( 
.A(n_2748),
.Y(n_3484)
);

AOI22xp33_ASAP7_75t_L g3485 ( 
.A1(n_3084),
.A2(n_2631),
.B1(n_2703),
.B2(n_2608),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3086),
.Y(n_3486)
);

NOR2xp33_ASAP7_75t_L g3487 ( 
.A(n_2885),
.B(n_2919),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_L g3488 ( 
.A1(n_3086),
.A2(n_2631),
.B1(n_2703),
.B2(n_2608),
.Y(n_3488)
);

A2O1A1Ixp33_ASAP7_75t_SL g3489 ( 
.A1(n_2818),
.A2(n_2400),
.B(n_2413),
.C(n_2367),
.Y(n_3489)
);

INVx8_ASAP7_75t_L g3490 ( 
.A(n_2809),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3091),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_SL g3492 ( 
.A(n_2807),
.B(n_2591),
.Y(n_3492)
);

AND2x4_ASAP7_75t_L g3493 ( 
.A(n_2811),
.B(n_2485),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_2929),
.B(n_2736),
.Y(n_3494)
);

NOR2xp33_ASAP7_75t_L g3495 ( 
.A(n_2919),
.B(n_2485),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3091),
.Y(n_3496)
);

OR2x2_ASAP7_75t_L g3497 ( 
.A(n_3159),
.B(n_1975),
.Y(n_3497)
);

NOR2xp33_ASAP7_75t_L g3498 ( 
.A(n_3028),
.B(n_2530),
.Y(n_3498)
);

OR2x6_ASAP7_75t_L g3499 ( 
.A(n_3159),
.B(n_2530),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_2936),
.B(n_2736),
.Y(n_3500)
);

OAI22xp5_ASAP7_75t_L g3501 ( 
.A1(n_2887),
.A2(n_2641),
.B1(n_2591),
.B2(n_2374),
.Y(n_3501)
);

AOI22xp5_ASAP7_75t_L g3502 ( 
.A1(n_2809),
.A2(n_2631),
.B1(n_2736),
.B2(n_2703),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_2936),
.B(n_2703),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_2936),
.B(n_2703),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3099),
.Y(n_3505)
);

AOI22xp5_ASAP7_75t_L g3506 ( 
.A1(n_2812),
.A2(n_2736),
.B1(n_2530),
.B2(n_2313),
.Y(n_3506)
);

INVx8_ASAP7_75t_L g3507 ( 
.A(n_2812),
.Y(n_3507)
);

AOI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_2812),
.A2(n_3000),
.B1(n_3021),
.B2(n_2990),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3099),
.Y(n_3509)
);

INVx3_ASAP7_75t_L g3510 ( 
.A(n_2748),
.Y(n_3510)
);

AOI22xp5_ASAP7_75t_L g3511 ( 
.A1(n_2990),
.A2(n_2736),
.B1(n_2530),
.B2(n_2641),
.Y(n_3511)
);

NOR2xp33_ASAP7_75t_L g3512 ( 
.A(n_3046),
.B(n_2500),
.Y(n_3512)
);

OR2x6_ASAP7_75t_L g3513 ( 
.A(n_3159),
.B(n_2851),
.Y(n_3513)
);

BUFx6f_ASAP7_75t_L g3514 ( 
.A(n_2847),
.Y(n_3514)
);

BUFx2_ASAP7_75t_L g3515 ( 
.A(n_2973),
.Y(n_3515)
);

NAND2xp33_ASAP7_75t_L g3516 ( 
.A(n_2835),
.B(n_2901),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_2977),
.B(n_2736),
.Y(n_3517)
);

AND2x6_ASAP7_75t_SL g3518 ( 
.A(n_3049),
.B(n_1672),
.Y(n_3518)
);

AOI22xp5_ASAP7_75t_L g3519 ( 
.A1(n_2990),
.A2(n_2338),
.B1(n_2589),
.B2(n_2639),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3100),
.Y(n_3520)
);

NOR2x1p5_ASAP7_75t_L g3521 ( 
.A(n_2976),
.B(n_1581),
.Y(n_3521)
);

BUFx3_ASAP7_75t_L g3522 ( 
.A(n_3083),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3105),
.Y(n_3523)
);

INVx1_ASAP7_75t_SL g3524 ( 
.A(n_3083),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3105),
.Y(n_3525)
);

CKINVDCx5p33_ASAP7_75t_R g3526 ( 
.A(n_3106),
.Y(n_3526)
);

INVx2_ASAP7_75t_L g3527 ( 
.A(n_3114),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_2977),
.B(n_2585),
.Y(n_3528)
);

BUFx3_ASAP7_75t_L g3529 ( 
.A(n_3327),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3213),
.Y(n_3530)
);

INVx3_ASAP7_75t_L g3531 ( 
.A(n_3195),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3220),
.Y(n_3532)
);

BUFx6f_ASAP7_75t_L g3533 ( 
.A(n_3331),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3180),
.Y(n_3534)
);

INVx2_ASAP7_75t_SL g3535 ( 
.A(n_3231),
.Y(n_3535)
);

INVx2_ASAP7_75t_SL g3536 ( 
.A(n_3231),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3179),
.B(n_3114),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3191),
.Y(n_3538)
);

BUFx6f_ASAP7_75t_L g3539 ( 
.A(n_3331),
.Y(n_3539)
);

AND2x4_ASAP7_75t_L g3540 ( 
.A(n_3214),
.B(n_2811),
.Y(n_3540)
);

OR2x2_ASAP7_75t_SL g3541 ( 
.A(n_3262),
.B(n_3118),
.Y(n_3541)
);

OR2x6_ASAP7_75t_L g3542 ( 
.A(n_3513),
.B(n_2851),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_3239),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3182),
.B(n_3126),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_SL g3545 ( 
.A(n_3290),
.B(n_3052),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3361),
.B(n_3126),
.Y(n_3546)
);

NOR2xp33_ASAP7_75t_L g3547 ( 
.A(n_3193),
.B(n_3069),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3361),
.B(n_3136),
.Y(n_3548)
);

NOR2xp33_ASAP7_75t_L g3549 ( 
.A(n_3193),
.B(n_3069),
.Y(n_3549)
);

AND2x4_ASAP7_75t_L g3550 ( 
.A(n_3214),
.B(n_3150),
.Y(n_3550)
);

CKINVDCx11_ASAP7_75t_R g3551 ( 
.A(n_3518),
.Y(n_3551)
);

INVx1_ASAP7_75t_SL g3552 ( 
.A(n_3261),
.Y(n_3552)
);

OR2x6_ASAP7_75t_L g3553 ( 
.A(n_3513),
.B(n_2838),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3364),
.B(n_3136),
.Y(n_3554)
);

CKINVDCx11_ASAP7_75t_R g3555 ( 
.A(n_3524),
.Y(n_3555)
);

NAND3xp33_ASAP7_75t_L g3556 ( 
.A(n_3290),
.B(n_1734),
.C(n_1807),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3204),
.Y(n_3557)
);

BUFx2_ASAP7_75t_L g3558 ( 
.A(n_3270),
.Y(n_3558)
);

INVx5_ASAP7_75t_L g3559 ( 
.A(n_3405),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3227),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3243),
.Y(n_3561)
);

AND2x4_ASAP7_75t_L g3562 ( 
.A(n_3375),
.B(n_3150),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3364),
.B(n_3142),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3249),
.Y(n_3564)
);

HB1xp67_ASAP7_75t_L g3565 ( 
.A(n_3345),
.Y(n_3565)
);

INVx4_ASAP7_75t_L g3566 ( 
.A(n_3435),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3245),
.Y(n_3567)
);

CKINVDCx20_ASAP7_75t_R g3568 ( 
.A(n_3278),
.Y(n_3568)
);

INVx3_ASAP7_75t_L g3569 ( 
.A(n_3195),
.Y(n_3569)
);

AOI22xp33_ASAP7_75t_L g3570 ( 
.A1(n_3443),
.A2(n_3135),
.B1(n_2822),
.B2(n_2891),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3185),
.B(n_3142),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_3255),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3420),
.B(n_3158),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3282),
.Y(n_3574)
);

INVx4_ASAP7_75t_L g3575 ( 
.A(n_3435),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3422),
.B(n_3158),
.Y(n_3576)
);

BUFx6f_ASAP7_75t_L g3577 ( 
.A(n_3405),
.Y(n_3577)
);

HB1xp67_ASAP7_75t_L g3578 ( 
.A(n_3345),
.Y(n_3578)
);

OR2x6_ASAP7_75t_L g3579 ( 
.A(n_3513),
.B(n_2838),
.Y(n_3579)
);

OR2x6_ASAP7_75t_L g3580 ( 
.A(n_3490),
.B(n_2838),
.Y(n_3580)
);

BUFx12f_ASAP7_75t_L g3581 ( 
.A(n_3278),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3284),
.Y(n_3582)
);

OR2x6_ASAP7_75t_L g3583 ( 
.A(n_3490),
.B(n_2838),
.Y(n_3583)
);

AOI22xp33_ASAP7_75t_L g3584 ( 
.A1(n_3443),
.A2(n_3268),
.B1(n_3211),
.B2(n_3306),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3289),
.Y(n_3585)
);

BUFx6f_ASAP7_75t_L g3586 ( 
.A(n_3405),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3291),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3311),
.Y(n_3588)
);

OR2x6_ASAP7_75t_L g3589 ( 
.A(n_3490),
.B(n_3054),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_SL g3590 ( 
.A(n_3306),
.B(n_3052),
.Y(n_3590)
);

AND2x4_ASAP7_75t_L g3591 ( 
.A(n_3375),
.B(n_3127),
.Y(n_3591)
);

OR2x6_ASAP7_75t_L g3592 ( 
.A(n_3507),
.B(n_3054),
.Y(n_3592)
);

BUFx3_ASAP7_75t_L g3593 ( 
.A(n_3374),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3313),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3325),
.Y(n_3595)
);

BUFx8_ASAP7_75t_SL g3596 ( 
.A(n_3312),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3226),
.B(n_2962),
.Y(n_3597)
);

NAND2xp33_ASAP7_75t_L g3598 ( 
.A(n_3320),
.B(n_2901),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3410),
.B(n_2964),
.Y(n_3599)
);

BUFx2_ASAP7_75t_L g3600 ( 
.A(n_3286),
.Y(n_3600)
);

AOI22xp5_ASAP7_75t_L g3601 ( 
.A1(n_3206),
.A2(n_3071),
.B1(n_3087),
.B2(n_3133),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3363),
.Y(n_3602)
);

AND2x4_ASAP7_75t_L g3603 ( 
.A(n_3493),
.B(n_3477),
.Y(n_3603)
);

INVx3_ASAP7_75t_SL g3604 ( 
.A(n_3358),
.Y(n_3604)
);

BUFx2_ASAP7_75t_L g3605 ( 
.A(n_3286),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3378),
.Y(n_3606)
);

NOR2xp33_ASAP7_75t_L g3607 ( 
.A(n_3196),
.B(n_3071),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3382),
.Y(n_3608)
);

INVx2_ASAP7_75t_SL g3609 ( 
.A(n_3294),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3383),
.Y(n_3610)
);

BUFx8_ASAP7_75t_L g3611 ( 
.A(n_3515),
.Y(n_3611)
);

AOI22xp5_ASAP7_75t_L g3612 ( 
.A1(n_3206),
.A2(n_3196),
.B1(n_3268),
.B2(n_3211),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3411),
.B(n_2965),
.Y(n_3613)
);

AOI22xp33_ASAP7_75t_L g3614 ( 
.A1(n_3308),
.A2(n_3135),
.B1(n_2822),
.B2(n_2971),
.Y(n_3614)
);

NAND2x1p5_ASAP7_75t_L g3615 ( 
.A(n_3435),
.B(n_3119),
.Y(n_3615)
);

BUFx2_ASAP7_75t_L g3616 ( 
.A(n_3221),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3387),
.Y(n_3617)
);

INVx4_ASAP7_75t_L g3618 ( 
.A(n_3435),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3380),
.B(n_2966),
.Y(n_3619)
);

NOR2xp33_ASAP7_75t_L g3620 ( 
.A(n_3426),
.B(n_3087),
.Y(n_3620)
);

INVx2_ASAP7_75t_L g3621 ( 
.A(n_3298),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3388),
.Y(n_3622)
);

INVx4_ASAP7_75t_L g3623 ( 
.A(n_3507),
.Y(n_3623)
);

BUFx2_ASAP7_75t_L g3624 ( 
.A(n_3222),
.Y(n_3624)
);

HB1xp67_ASAP7_75t_L g3625 ( 
.A(n_3400),
.Y(n_3625)
);

AOI22xp5_ASAP7_75t_L g3626 ( 
.A1(n_3183),
.A2(n_3133),
.B1(n_3162),
.B2(n_3102),
.Y(n_3626)
);

BUFx3_ASAP7_75t_L g3627 ( 
.A(n_3392),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_SL g3628 ( 
.A(n_3265),
.B(n_3076),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3395),
.Y(n_3629)
);

INVx3_ASAP7_75t_L g3630 ( 
.A(n_3274),
.Y(n_3630)
);

NOR2xp33_ASAP7_75t_L g3631 ( 
.A(n_3183),
.B(n_2977),
.Y(n_3631)
);

NOR2xp33_ASAP7_75t_L g3632 ( 
.A(n_3256),
.B(n_2982),
.Y(n_3632)
);

INVx2_ASAP7_75t_L g3633 ( 
.A(n_3315),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3399),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3318),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3413),
.B(n_2981),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3401),
.Y(n_3637)
);

INVx2_ASAP7_75t_L g3638 ( 
.A(n_3339),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_3230),
.B(n_3297),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3403),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3414),
.Y(n_3641)
);

INVxp67_ASAP7_75t_L g3642 ( 
.A(n_3427),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3189),
.B(n_2983),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3424),
.Y(n_3644)
);

AOI22xp33_ASAP7_75t_L g3645 ( 
.A1(n_3202),
.A2(n_3135),
.B1(n_2822),
.B2(n_2988),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3431),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3451),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3456),
.Y(n_3648)
);

INVx4_ASAP7_75t_L g3649 ( 
.A(n_3507),
.Y(n_3649)
);

OAI22xp5_ASAP7_75t_L g3650 ( 
.A1(n_3202),
.A2(n_3275),
.B1(n_3293),
.B2(n_3259),
.Y(n_3650)
);

BUFx6f_ASAP7_75t_L g3651 ( 
.A(n_3405),
.Y(n_3651)
);

INVx3_ASAP7_75t_L g3652 ( 
.A(n_3274),
.Y(n_3652)
);

BUFx3_ASAP7_75t_L g3653 ( 
.A(n_3186),
.Y(n_3653)
);

INVx3_ASAP7_75t_L g3654 ( 
.A(n_3303),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_3360),
.Y(n_3655)
);

AND2x4_ASAP7_75t_L g3656 ( 
.A(n_3493),
.B(n_3074),
.Y(n_3656)
);

INVx3_ASAP7_75t_L g3657 ( 
.A(n_3303),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3197),
.B(n_2984),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3198),
.B(n_2991),
.Y(n_3659)
);

BUFx4f_ASAP7_75t_L g3660 ( 
.A(n_3190),
.Y(n_3660)
);

BUFx2_ASAP7_75t_L g3661 ( 
.A(n_3299),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3468),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3199),
.B(n_3203),
.Y(n_3663)
);

AND2x4_ASAP7_75t_L g3664 ( 
.A(n_3499),
.B(n_3074),
.Y(n_3664)
);

AND2x2_ASAP7_75t_SL g3665 ( 
.A(n_3516),
.B(n_2764),
.Y(n_3665)
);

BUFx6f_ASAP7_75t_L g3666 ( 
.A(n_3407),
.Y(n_3666)
);

NOR2x1_ASAP7_75t_L g3667 ( 
.A(n_3480),
.B(n_3080),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_SL g3668 ( 
.A(n_3266),
.B(n_3011),
.Y(n_3668)
);

BUFx6f_ASAP7_75t_L g3669 ( 
.A(n_3407),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_3469),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3473),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3244),
.B(n_3080),
.Y(n_3672)
);

BUFx6f_ASAP7_75t_L g3673 ( 
.A(n_3407),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3207),
.B(n_2993),
.Y(n_3674)
);

AOI22xp33_ASAP7_75t_L g3675 ( 
.A1(n_3215),
.A2(n_2997),
.B1(n_3003),
.B2(n_2996),
.Y(n_3675)
);

CKINVDCx5p33_ASAP7_75t_R g3676 ( 
.A(n_3452),
.Y(n_3676)
);

NOR2xp33_ASAP7_75t_L g3677 ( 
.A(n_3428),
.B(n_1797),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_3208),
.B(n_3004),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3486),
.Y(n_3679)
);

CKINVDCx11_ASAP7_75t_R g3680 ( 
.A(n_3522),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3491),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3496),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_SL g3683 ( 
.A(n_3384),
.B(n_3076),
.Y(n_3683)
);

INVxp67_ASAP7_75t_SL g3684 ( 
.A(n_3240),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3505),
.Y(n_3685)
);

HB1xp67_ASAP7_75t_L g3686 ( 
.A(n_3446),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3210),
.B(n_3223),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3509),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3368),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_3225),
.B(n_3007),
.Y(n_3690)
);

INVx1_ASAP7_75t_SL g3691 ( 
.A(n_3260),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_SL g3692 ( 
.A(n_3385),
.B(n_3076),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_3228),
.B(n_3389),
.Y(n_3693)
);

INVx2_ASAP7_75t_L g3694 ( 
.A(n_3372),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3520),
.Y(n_3695)
);

CKINVDCx8_ASAP7_75t_R g3696 ( 
.A(n_3526),
.Y(n_3696)
);

INVx5_ASAP7_75t_L g3697 ( 
.A(n_3407),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3523),
.Y(n_3698)
);

AOI22xp33_ASAP7_75t_L g3699 ( 
.A1(n_3215),
.A2(n_3010),
.B1(n_3013),
.B2(n_3008),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3525),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_SL g3701 ( 
.A(n_3447),
.B(n_3119),
.Y(n_3701)
);

AOI22xp33_ASAP7_75t_L g3702 ( 
.A1(n_3367),
.A2(n_3020),
.B1(n_3025),
.B2(n_3018),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3377),
.Y(n_3703)
);

AND2x4_ASAP7_75t_L g3704 ( 
.A(n_3499),
.B(n_3096),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3417),
.Y(n_3705)
);

BUFx6f_ASAP7_75t_L g3706 ( 
.A(n_3514),
.Y(n_3706)
);

BUFx6f_ASAP7_75t_L g3707 ( 
.A(n_3514),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3241),
.B(n_3027),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3269),
.B(n_3030),
.Y(n_3709)
);

NOR2xp33_ASAP7_75t_L g3710 ( 
.A(n_3428),
.B(n_2742),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3437),
.Y(n_3711)
);

BUFx3_ASAP7_75t_L g3712 ( 
.A(n_3423),
.Y(n_3712)
);

NOR2xp67_ASAP7_75t_L g3713 ( 
.A(n_3356),
.B(n_3147),
.Y(n_3713)
);

AOI22xp5_ASAP7_75t_L g3714 ( 
.A1(n_3242),
.A2(n_1901),
.B1(n_1905),
.B2(n_3000),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3461),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3478),
.Y(n_3716)
);

BUFx4f_ASAP7_75t_L g3717 ( 
.A(n_3466),
.Y(n_3717)
);

AOI22xp5_ASAP7_75t_L g3718 ( 
.A1(n_3242),
.A2(n_1905),
.B1(n_3021),
.B2(n_3000),
.Y(n_3718)
);

INVx3_ASAP7_75t_L g3719 ( 
.A(n_3432),
.Y(n_3719)
);

AO22x1_ASAP7_75t_L g3720 ( 
.A1(n_3460),
.A2(n_1905),
.B1(n_1734),
.B2(n_3455),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3482),
.Y(n_3721)
);

HB1xp67_ASAP7_75t_L g3722 ( 
.A(n_3446),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3296),
.B(n_3021),
.Y(n_3723)
);

BUFx4f_ASAP7_75t_L g3724 ( 
.A(n_3479),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3527),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3397),
.Y(n_3726)
);

INVx3_ASAP7_75t_L g3727 ( 
.A(n_3432),
.Y(n_3727)
);

INVx3_ASAP7_75t_L g3728 ( 
.A(n_3484),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3330),
.B(n_3035),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_SL g3730 ( 
.A(n_3283),
.B(n_3119),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_SL g3731 ( 
.A(n_3283),
.B(n_3125),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_3232),
.B(n_3042),
.Y(n_3732)
);

HB1xp67_ASAP7_75t_L g3733 ( 
.A(n_3448),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3440),
.B(n_2743),
.Y(n_3734)
);

BUFx3_ASAP7_75t_L g3735 ( 
.A(n_3188),
.Y(n_3735)
);

BUFx6f_ASAP7_75t_L g3736 ( 
.A(n_3514),
.Y(n_3736)
);

AND2x4_ASAP7_75t_L g3737 ( 
.A(n_3258),
.B(n_3096),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3398),
.Y(n_3738)
);

NOR2xp33_ASAP7_75t_L g3739 ( 
.A(n_3440),
.B(n_2754),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_SL g3740 ( 
.A(n_3257),
.B(n_3125),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3406),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3333),
.Y(n_3742)
);

INVx5_ASAP7_75t_L g3743 ( 
.A(n_3514),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3234),
.B(n_3044),
.Y(n_3744)
);

BUFx3_ASAP7_75t_L g3745 ( 
.A(n_3335),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3237),
.B(n_3048),
.Y(n_3746)
);

AND2x4_ASAP7_75t_L g3747 ( 
.A(n_3444),
.B(n_3508),
.Y(n_3747)
);

CKINVDCx5p33_ASAP7_75t_R g3748 ( 
.A(n_3436),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3338),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3341),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3238),
.B(n_3050),
.Y(n_3751)
);

AND2x4_ASAP7_75t_L g3752 ( 
.A(n_3487),
.B(n_3022),
.Y(n_3752)
);

INVx3_ASAP7_75t_L g3753 ( 
.A(n_3484),
.Y(n_3753)
);

NOR2x1p5_ASAP7_75t_L g3754 ( 
.A(n_3381),
.B(n_2740),
.Y(n_3754)
);

INVx5_ASAP7_75t_L g3755 ( 
.A(n_3510),
.Y(n_3755)
);

BUFx4f_ASAP7_75t_L g3756 ( 
.A(n_3359),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_SL g3757 ( 
.A(n_3314),
.B(n_3125),
.Y(n_3757)
);

CKINVDCx5p33_ASAP7_75t_R g3758 ( 
.A(n_3467),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3342),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3347),
.Y(n_3760)
);

AOI22xp5_ASAP7_75t_L g3761 ( 
.A1(n_3247),
.A2(n_3059),
.B1(n_3060),
.B2(n_3022),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3348),
.Y(n_3762)
);

INVx3_ASAP7_75t_L g3763 ( 
.A(n_3510),
.Y(n_3763)
);

AND2x4_ASAP7_75t_L g3764 ( 
.A(n_3487),
.B(n_3059),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_3301),
.B(n_3305),
.Y(n_3765)
);

BUFx3_ASAP7_75t_L g3766 ( 
.A(n_3467),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3350),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3376),
.Y(n_3768)
);

HB1xp67_ASAP7_75t_L g3769 ( 
.A(n_3449),
.Y(n_3769)
);

AND2x2_ASAP7_75t_SL g3770 ( 
.A(n_3352),
.B(n_2764),
.Y(n_3770)
);

INVx3_ASAP7_75t_SL g3771 ( 
.A(n_3470),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3307),
.Y(n_3772)
);

AO22x1_ASAP7_75t_L g3773 ( 
.A1(n_3460),
.A2(n_3055),
.B1(n_1099),
.B2(n_2763),
.Y(n_3773)
);

OR2x2_ASAP7_75t_L g3774 ( 
.A(n_3329),
.B(n_2758),
.Y(n_3774)
);

INVx2_ASAP7_75t_SL g3775 ( 
.A(n_3271),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_SL g3776 ( 
.A(n_3254),
.B(n_3130),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3309),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3310),
.B(n_3053),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3317),
.B(n_3322),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3324),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3248),
.B(n_3056),
.Y(n_3781)
);

BUFx3_ASAP7_75t_L g3782 ( 
.A(n_3497),
.Y(n_3782)
);

INVx3_ASAP7_75t_L g3783 ( 
.A(n_3209),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3250),
.Y(n_3784)
);

AND2x4_ASAP7_75t_L g3785 ( 
.A(n_3184),
.B(n_3059),
.Y(n_3785)
);

INVx5_ASAP7_75t_L g3786 ( 
.A(n_3209),
.Y(n_3786)
);

INVx4_ASAP7_75t_L g3787 ( 
.A(n_3295),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3252),
.B(n_3253),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3263),
.Y(n_3789)
);

INVx2_ASAP7_75t_SL g3790 ( 
.A(n_3521),
.Y(n_3790)
);

BUFx3_ASAP7_75t_L g3791 ( 
.A(n_3474),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3267),
.Y(n_3792)
);

BUFx6f_ASAP7_75t_L g3793 ( 
.A(n_3295),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3430),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_3287),
.B(n_3064),
.Y(n_3795)
);

BUFx2_ASAP7_75t_R g3796 ( 
.A(n_3187),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3288),
.Y(n_3797)
);

AND2x4_ASAP7_75t_L g3798 ( 
.A(n_3474),
.B(n_3060),
.Y(n_3798)
);

HB1xp67_ASAP7_75t_L g3799 ( 
.A(n_3409),
.Y(n_3799)
);

INVxp67_ASAP7_75t_L g3800 ( 
.A(n_3427),
.Y(n_3800)
);

CKINVDCx20_ASAP7_75t_R g3801 ( 
.A(n_3498),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_3390),
.B(n_3068),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3302),
.B(n_3073),
.Y(n_3803)
);

INVx3_ASAP7_75t_L g3804 ( 
.A(n_3340),
.Y(n_3804)
);

BUFx8_ASAP7_75t_L g3805 ( 
.A(n_3279),
.Y(n_3805)
);

INVx2_ASAP7_75t_L g3806 ( 
.A(n_3433),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3439),
.Y(n_3807)
);

CKINVDCx20_ASAP7_75t_R g3808 ( 
.A(n_3498),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3441),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3302),
.B(n_3077),
.Y(n_3810)
);

BUFx2_ASAP7_75t_L g3811 ( 
.A(n_3224),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3409),
.Y(n_3812)
);

HB1xp67_ASAP7_75t_L g3813 ( 
.A(n_3415),
.Y(n_3813)
);

AOI22xp5_ASAP7_75t_L g3814 ( 
.A1(n_3247),
.A2(n_3060),
.B1(n_3122),
.B2(n_3078),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3415),
.Y(n_3815)
);

OR2x2_ASAP7_75t_L g3816 ( 
.A(n_3212),
.B(n_2766),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_3453),
.Y(n_3817)
);

AND2x4_ASAP7_75t_L g3818 ( 
.A(n_3481),
.B(n_3078),
.Y(n_3818)
);

AO22x1_ASAP7_75t_L g3819 ( 
.A1(n_3455),
.A2(n_3055),
.B1(n_3122),
.B2(n_3078),
.Y(n_3819)
);

AND2x4_ASAP7_75t_L g3820 ( 
.A(n_3481),
.B(n_3483),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3416),
.Y(n_3821)
);

AND2x2_ASAP7_75t_L g3822 ( 
.A(n_3212),
.B(n_3122),
.Y(n_3822)
);

INVx2_ASAP7_75t_L g3823 ( 
.A(n_3457),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_SL g3824 ( 
.A(n_3396),
.B(n_3130),
.Y(n_3824)
);

AOI22xp5_ASAP7_75t_SL g3825 ( 
.A1(n_3445),
.A2(n_3026),
.B1(n_745),
.B2(n_746),
.Y(n_3825)
);

INVx1_ASAP7_75t_SL g3826 ( 
.A(n_3219),
.Y(n_3826)
);

AND2x2_ASAP7_75t_L g3827 ( 
.A(n_3219),
.B(n_3174),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_SL g3828 ( 
.A(n_3396),
.B(n_3130),
.Y(n_3828)
);

O2A1O1Ixp33_ASAP7_75t_L g3829 ( 
.A1(n_3438),
.A2(n_3092),
.B(n_3082),
.C(n_3085),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3319),
.B(n_3416),
.Y(n_3830)
);

NAND2x1p5_ASAP7_75t_L g3831 ( 
.A(n_3343),
.B(n_2752),
.Y(n_3831)
);

AOI22xp33_ASAP7_75t_L g3832 ( 
.A1(n_3445),
.A2(n_3110),
.B1(n_3157),
.B2(n_3095),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3319),
.B(n_3079),
.Y(n_3833)
);

NAND2xp33_ASAP7_75t_L g3834 ( 
.A(n_3320),
.B(n_2901),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3354),
.Y(n_3835)
);

BUFx2_ASAP7_75t_L g3836 ( 
.A(n_3340),
.Y(n_3836)
);

BUFx3_ASAP7_75t_L g3837 ( 
.A(n_3495),
.Y(n_3837)
);

OAI21x1_ASAP7_75t_L g3838 ( 
.A1(n_3334),
.A2(n_3037),
.B(n_2732),
.Y(n_3838)
);

BUFx4f_ASAP7_75t_L g3839 ( 
.A(n_3246),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3373),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3386),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_3349),
.Y(n_3842)
);

BUFx4f_ASAP7_75t_L g3843 ( 
.A(n_3246),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3218),
.B(n_3404),
.Y(n_3844)
);

AND2x4_ASAP7_75t_L g3845 ( 
.A(n_3492),
.B(n_3134),
.Y(n_3845)
);

AND2x6_ASAP7_75t_SL g3846 ( 
.A(n_3512),
.B(n_3026),
.Y(n_3846)
);

NOR2xp33_ASAP7_75t_L g3847 ( 
.A(n_3404),
.B(n_3167),
.Y(n_3847)
);

AOI22xp33_ASAP7_75t_L g3848 ( 
.A1(n_3216),
.A2(n_3138),
.B1(n_3161),
.B2(n_3111),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3353),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3462),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_3386),
.B(n_3098),
.Y(n_3851)
);

BUFx3_ASAP7_75t_L g3852 ( 
.A(n_3512),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3394),
.Y(n_3853)
);

BUFx4f_ASAP7_75t_L g3854 ( 
.A(n_3412),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_3275),
.B(n_3293),
.Y(n_3855)
);

NOR2xp33_ASAP7_75t_L g3856 ( 
.A(n_3408),
.B(n_3168),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3464),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3703),
.Y(n_3858)
);

INVx5_ASAP7_75t_L g3859 ( 
.A(n_3566),
.Y(n_3859)
);

AND2x2_ASAP7_75t_L g3860 ( 
.A(n_3612),
.B(n_3218),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3584),
.B(n_3229),
.Y(n_3861)
);

AOI21xp5_ASAP7_75t_L g3862 ( 
.A1(n_3598),
.A2(n_3834),
.B(n_3285),
.Y(n_3862)
);

AOI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_3628),
.A2(n_3321),
.B(n_3316),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_SL g3864 ( 
.A(n_3826),
.B(n_3408),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3772),
.B(n_3336),
.Y(n_3865)
);

INVx3_ASAP7_75t_L g3866 ( 
.A(n_3839),
.Y(n_3866)
);

AOI21xp5_ASAP7_75t_L g3867 ( 
.A1(n_3628),
.A2(n_3321),
.B(n_3316),
.Y(n_3867)
);

O2A1O1Ixp33_ASAP7_75t_L g3868 ( 
.A1(n_3547),
.A2(n_3277),
.B(n_3442),
.C(n_3476),
.Y(n_3868)
);

AND2x4_ASAP7_75t_L g3869 ( 
.A(n_3562),
.B(n_3402),
.Y(n_3869)
);

AOI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_3590),
.A2(n_3326),
.B(n_3323),
.Y(n_3870)
);

AOI22xp5_ASAP7_75t_L g3871 ( 
.A1(n_3549),
.A2(n_3391),
.B1(n_3328),
.B2(n_3458),
.Y(n_3871)
);

BUFx6f_ASAP7_75t_L g3872 ( 
.A(n_3533),
.Y(n_3872)
);

AOI21xp5_ASAP7_75t_L g3873 ( 
.A1(n_3590),
.A2(n_3326),
.B(n_3323),
.Y(n_3873)
);

AOI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_3684),
.A2(n_3344),
.B(n_3280),
.Y(n_3874)
);

AND2x4_ASAP7_75t_L g3875 ( 
.A(n_3562),
.B(n_3418),
.Y(n_3875)
);

HB1xp67_ASAP7_75t_L g3876 ( 
.A(n_3625),
.Y(n_3876)
);

INVxp67_ASAP7_75t_SL g3877 ( 
.A(n_3625),
.Y(n_3877)
);

NOR2xp33_ASAP7_75t_L g3878 ( 
.A(n_3549),
.B(n_1600),
.Y(n_3878)
);

O2A1O1Ixp33_ASAP7_75t_SL g3879 ( 
.A1(n_3693),
.A2(n_3217),
.B(n_3187),
.C(n_3277),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3705),
.Y(n_3880)
);

INVx2_ASAP7_75t_L g3881 ( 
.A(n_3561),
.Y(n_3881)
);

AND2x4_ASAP7_75t_L g3882 ( 
.A(n_3550),
.B(n_3200),
.Y(n_3882)
);

NOR2xp33_ASAP7_75t_R g3883 ( 
.A(n_3676),
.B(n_3174),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3584),
.B(n_3229),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_3777),
.B(n_3236),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3780),
.B(n_3236),
.Y(n_3886)
);

O2A1O1Ixp33_ASAP7_75t_L g3887 ( 
.A1(n_3607),
.A2(n_3337),
.B(n_3365),
.C(n_3351),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3564),
.Y(n_3888)
);

OAI22x1_ASAP7_75t_L g3889 ( 
.A1(n_3601),
.A2(n_3511),
.B1(n_2405),
.B2(n_2909),
.Y(n_3889)
);

NAND2xp33_ASAP7_75t_SL g3890 ( 
.A(n_3533),
.B(n_2405),
.Y(n_3890)
);

A2O1A1Ixp33_ASAP7_75t_SL g3891 ( 
.A1(n_3620),
.A2(n_3259),
.B(n_3506),
.C(n_3454),
.Y(n_3891)
);

NOR2xp33_ASAP7_75t_L g3892 ( 
.A(n_3620),
.B(n_3677),
.Y(n_3892)
);

A2O1A1Ixp33_ASAP7_75t_L g3893 ( 
.A1(n_3632),
.A2(n_3346),
.B(n_3192),
.C(n_2947),
.Y(n_3893)
);

AOI21xp5_ASAP7_75t_L g3894 ( 
.A1(n_3684),
.A2(n_3344),
.B(n_3201),
.Y(n_3894)
);

AOI22x1_ASAP7_75t_L g3895 ( 
.A1(n_3835),
.A2(n_3117),
.B1(n_3121),
.B2(n_3113),
.Y(n_3895)
);

NOR2xp33_ASAP7_75t_L g3896 ( 
.A(n_3677),
.B(n_1600),
.Y(n_3896)
);

NOR2xp33_ASAP7_75t_L g3897 ( 
.A(n_3827),
.B(n_1601),
.Y(n_3897)
);

AO21x1_ASAP7_75t_L g3898 ( 
.A1(n_3650),
.A2(n_3365),
.B(n_3351),
.Y(n_3898)
);

BUFx2_ASAP7_75t_L g3899 ( 
.A(n_3558),
.Y(n_3899)
);

AND2x4_ASAP7_75t_L g3900 ( 
.A(n_3550),
.B(n_3205),
.Y(n_3900)
);

A2O1A1Ixp33_ASAP7_75t_L g3901 ( 
.A1(n_3632),
.A2(n_3233),
.B(n_3251),
.C(n_3502),
.Y(n_3901)
);

CKINVDCx5p33_ASAP7_75t_R g3902 ( 
.A(n_3596),
.Y(n_3902)
);

AOI21xp5_ASAP7_75t_L g3903 ( 
.A1(n_3545),
.A2(n_2746),
.B(n_3355),
.Y(n_3903)
);

NOR3xp33_ASAP7_75t_SL g3904 ( 
.A(n_3556),
.B(n_747),
.C(n_742),
.Y(n_3904)
);

NOR2xp33_ASAP7_75t_L g3905 ( 
.A(n_3642),
.B(n_1601),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3784),
.B(n_3194),
.Y(n_3906)
);

AOI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3545),
.A2(n_2746),
.B(n_3393),
.Y(n_3907)
);

BUFx6f_ASAP7_75t_L g3908 ( 
.A(n_3533),
.Y(n_3908)
);

AND2x4_ASAP7_75t_L g3909 ( 
.A(n_3540),
.B(n_3264),
.Y(n_3909)
);

NOR3xp33_ASAP7_75t_L g3910 ( 
.A(n_3773),
.B(n_3337),
.C(n_1508),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3789),
.B(n_3792),
.Y(n_3911)
);

INVxp67_ASAP7_75t_SL g3912 ( 
.A(n_3565),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3711),
.Y(n_3913)
);

OAI21xp5_ASAP7_75t_L g3914 ( 
.A1(n_3757),
.A2(n_3740),
.B(n_3829),
.Y(n_3914)
);

OR2x6_ASAP7_75t_L g3915 ( 
.A(n_3553),
.B(n_3217),
.Y(n_3915)
);

OAI22xp5_ASAP7_75t_L g3916 ( 
.A1(n_3650),
.A2(n_3332),
.B1(n_3251),
.B2(n_3450),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3740),
.A2(n_3366),
.B(n_3362),
.Y(n_3917)
);

A2O1A1Ixp33_ASAP7_75t_L g3918 ( 
.A1(n_3710),
.A2(n_3517),
.B(n_3504),
.C(n_3500),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_SL g3919 ( 
.A(n_3642),
.B(n_3332),
.Y(n_3919)
);

AO32x1_ASAP7_75t_L g3920 ( 
.A1(n_3842),
.A2(n_3170),
.A3(n_3129),
.B1(n_3140),
.B2(n_3128),
.Y(n_3920)
);

HB1xp67_ASAP7_75t_L g3921 ( 
.A(n_3565),
.Y(n_3921)
);

AOI22xp33_ASAP7_75t_L g3922 ( 
.A1(n_3747),
.A2(n_3471),
.B1(n_3472),
.B2(n_3503),
.Y(n_3922)
);

OAI22xp5_ASAP7_75t_L g3923 ( 
.A1(n_3710),
.A2(n_3454),
.B1(n_3463),
.B2(n_3450),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_SL g3924 ( 
.A(n_3800),
.B(n_3528),
.Y(n_3924)
);

INVxp67_ASAP7_75t_SL g3925 ( 
.A(n_3578),
.Y(n_3925)
);

BUFx6f_ASAP7_75t_L g3926 ( 
.A(n_3539),
.Y(n_3926)
);

INVx4_ASAP7_75t_L g3927 ( 
.A(n_3539),
.Y(n_3927)
);

AOI22xp33_ASAP7_75t_L g3928 ( 
.A1(n_3747),
.A2(n_3475),
.B1(n_3494),
.B2(n_3134),
.Y(n_3928)
);

AOI22xp5_ASAP7_75t_L g3929 ( 
.A1(n_3801),
.A2(n_3808),
.B1(n_3758),
.B2(n_3718),
.Y(n_3929)
);

INVx2_ASAP7_75t_L g3930 ( 
.A(n_3572),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3822),
.B(n_1457),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3715),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_SL g3933 ( 
.A(n_3800),
.B(n_2847),
.Y(n_3933)
);

O2A1O1Ixp5_ASAP7_75t_SL g3934 ( 
.A1(n_3757),
.A2(n_828),
.B(n_834),
.C(n_829),
.Y(n_3934)
);

AND2x2_ASAP7_75t_L g3935 ( 
.A(n_3672),
.B(n_1515),
.Y(n_3935)
);

XOR2x2_ASAP7_75t_L g3936 ( 
.A(n_3825),
.B(n_2445),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_L g3937 ( 
.A(n_3797),
.B(n_3726),
.Y(n_3937)
);

BUFx6f_ASAP7_75t_L g3938 ( 
.A(n_3539),
.Y(n_3938)
);

BUFx12f_ASAP7_75t_L g3939 ( 
.A(n_3555),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_SL g3940 ( 
.A(n_3734),
.B(n_2847),
.Y(n_3940)
);

O2A1O1Ixp33_ASAP7_75t_L g3941 ( 
.A1(n_3734),
.A2(n_1530),
.B(n_828),
.C(n_834),
.Y(n_3941)
);

OAI22xp5_ASAP7_75t_L g3942 ( 
.A1(n_3739),
.A2(n_3465),
.B1(n_3485),
.B2(n_3463),
.Y(n_3942)
);

BUFx8_ASAP7_75t_SL g3943 ( 
.A(n_3581),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_SL g3944 ( 
.A(n_3739),
.B(n_2847),
.Y(n_3944)
);

A2O1A1Ixp33_ASAP7_75t_L g3945 ( 
.A1(n_3631),
.A2(n_3016),
.B(n_2887),
.C(n_3181),
.Y(n_3945)
);

NAND2x1_ASAP7_75t_L g3946 ( 
.A(n_3553),
.B(n_2752),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3716),
.Y(n_3947)
);

AOI21x1_ASAP7_75t_L g3948 ( 
.A1(n_3730),
.A2(n_3419),
.B(n_3371),
.Y(n_3948)
);

AOI21xp5_ASAP7_75t_L g3949 ( 
.A1(n_3683),
.A2(n_3370),
.B(n_3369),
.Y(n_3949)
);

A2O1A1Ixp33_ASAP7_75t_L g3950 ( 
.A1(n_3631),
.A2(n_3016),
.B(n_2887),
.C(n_3235),
.Y(n_3950)
);

AOI21xp5_ASAP7_75t_L g3951 ( 
.A1(n_3692),
.A2(n_3370),
.B(n_3369),
.Y(n_3951)
);

AOI21xp5_ASAP7_75t_L g3952 ( 
.A1(n_3692),
.A2(n_3731),
.B(n_3730),
.Y(n_3952)
);

NOR2xp33_ASAP7_75t_SL g3953 ( 
.A(n_3805),
.B(n_3665),
.Y(n_3953)
);

AOI21x1_ASAP7_75t_L g3954 ( 
.A1(n_3731),
.A2(n_3425),
.B(n_3371),
.Y(n_3954)
);

NOR2xp33_ASAP7_75t_L g3955 ( 
.A(n_3735),
.B(n_1608),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3738),
.B(n_3144),
.Y(n_3956)
);

AOI21x1_ASAP7_75t_L g3957 ( 
.A1(n_3701),
.A2(n_3429),
.B(n_3425),
.Y(n_3957)
);

OAI22xp5_ASAP7_75t_L g3958 ( 
.A1(n_3812),
.A2(n_3465),
.B1(n_3488),
.B2(n_3485),
.Y(n_3958)
);

BUFx6f_ASAP7_75t_L g3959 ( 
.A(n_3660),
.Y(n_3959)
);

AOI21xp5_ASAP7_75t_L g3960 ( 
.A1(n_3770),
.A2(n_3276),
.B(n_2957),
.Y(n_3960)
);

AOI21xp5_ASAP7_75t_L g3961 ( 
.A1(n_3770),
.A2(n_3276),
.B(n_3005),
.Y(n_3961)
);

INVx6_ASAP7_75t_L g3962 ( 
.A(n_3805),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_SL g3963 ( 
.A(n_3756),
.B(n_2916),
.Y(n_3963)
);

A2O1A1Ixp33_ASAP7_75t_L g3964 ( 
.A1(n_3840),
.A2(n_3847),
.B(n_3856),
.C(n_3724),
.Y(n_3964)
);

NOR2xp33_ASAP7_75t_L g3965 ( 
.A(n_3791),
.B(n_1608),
.Y(n_3965)
);

INVx1_ASAP7_75t_SL g3966 ( 
.A(n_3691),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3741),
.B(n_3153),
.Y(n_3967)
);

O2A1O1Ixp33_ASAP7_75t_L g3968 ( 
.A1(n_3668),
.A2(n_829),
.B(n_838),
.C(n_837),
.Y(n_3968)
);

A2O1A1Ixp33_ASAP7_75t_SL g3969 ( 
.A1(n_3848),
.A2(n_3488),
.B(n_2872),
.C(n_3160),
.Y(n_3969)
);

AOI21xp5_ASAP7_75t_L g3970 ( 
.A1(n_3693),
.A2(n_3062),
.B(n_2899),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_3807),
.B(n_3809),
.Y(n_3971)
);

NAND2xp33_ASAP7_75t_L g3972 ( 
.A(n_3832),
.B(n_3320),
.Y(n_3972)
);

A2O1A1Ixp33_ASAP7_75t_L g3973 ( 
.A1(n_3847),
.A2(n_3016),
.B(n_3501),
.C(n_2928),
.Y(n_3973)
);

AOI22xp5_ASAP7_75t_L g3974 ( 
.A1(n_3626),
.A2(n_1611),
.B1(n_3300),
.B2(n_3292),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3534),
.Y(n_3975)
);

HB1xp67_ASAP7_75t_L g3976 ( 
.A(n_3578),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3663),
.B(n_3379),
.Y(n_3977)
);

NOR2xp33_ASAP7_75t_L g3978 ( 
.A(n_3837),
.B(n_1611),
.Y(n_3978)
);

NOR2xp33_ASAP7_75t_L g3979 ( 
.A(n_3552),
.B(n_2481),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3663),
.B(n_3379),
.Y(n_3980)
);

INVx1_ASAP7_75t_SL g3981 ( 
.A(n_3600),
.Y(n_3981)
);

NOR3xp33_ASAP7_75t_L g3982 ( 
.A(n_3720),
.B(n_1362),
.C(n_1359),
.Y(n_3982)
);

CKINVDCx20_ASAP7_75t_R g3983 ( 
.A(n_3568),
.Y(n_3983)
);

NAND2x1p5_ASAP7_75t_L g3984 ( 
.A(n_3755),
.B(n_2752),
.Y(n_3984)
);

O2A1O1Ixp33_ASAP7_75t_L g3985 ( 
.A1(n_3830),
.A2(n_837),
.B(n_840),
.C(n_838),
.Y(n_3985)
);

NOR2xp33_ASAP7_75t_L g3986 ( 
.A(n_3766),
.B(n_2582),
.Y(n_3986)
);

INVx4_ASAP7_75t_L g3987 ( 
.A(n_3786),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3802),
.A2(n_2901),
.B(n_3429),
.Y(n_3988)
);

NAND2x1p5_ASAP7_75t_L g3989 ( 
.A(n_3755),
.B(n_2755),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_3742),
.B(n_3166),
.Y(n_3990)
);

BUFx6f_ASAP7_75t_L g3991 ( 
.A(n_3660),
.Y(n_3991)
);

OAI22xp5_ASAP7_75t_L g3992 ( 
.A1(n_3815),
.A2(n_2974),
.B1(n_3097),
.B2(n_3057),
.Y(n_3992)
);

A2O1A1Ixp33_ASAP7_75t_L g3993 ( 
.A1(n_3856),
.A2(n_3519),
.B(n_3281),
.C(n_3152),
.Y(n_3993)
);

NAND3xp33_ASAP7_75t_SL g3994 ( 
.A(n_3714),
.B(n_751),
.C(n_749),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_SL g3995 ( 
.A(n_3756),
.B(n_2856),
.Y(n_3995)
);

INVx3_ASAP7_75t_L g3996 ( 
.A(n_3839),
.Y(n_3996)
);

AOI22xp33_ASAP7_75t_L g3997 ( 
.A1(n_3745),
.A2(n_3173),
.B1(n_3172),
.B2(n_3175),
.Y(n_3997)
);

BUFx10_ASAP7_75t_L g3998 ( 
.A(n_3846),
.Y(n_3998)
);

AND2x4_ASAP7_75t_L g3999 ( 
.A(n_3540),
.B(n_3591),
.Y(n_3999)
);

AOI21xp5_ASAP7_75t_L g4000 ( 
.A1(n_3802),
.A2(n_2901),
.B(n_3489),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_SL g4001 ( 
.A(n_3724),
.B(n_2856),
.Y(n_4001)
);

OAI22xp5_ASAP7_75t_L g4002 ( 
.A1(n_3821),
.A2(n_2934),
.B1(n_2916),
.B2(n_2856),
.Y(n_4002)
);

AND2x2_ASAP7_75t_L g4003 ( 
.A(n_3591),
.B(n_1426),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_L g4004 ( 
.A(n_3749),
.B(n_2767),
.Y(n_4004)
);

INVx3_ASAP7_75t_L g4005 ( 
.A(n_3843),
.Y(n_4005)
);

AOI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_3636),
.A2(n_3489),
.B(n_3357),
.Y(n_4006)
);

OR2x6_ASAP7_75t_L g4007 ( 
.A(n_3553),
.B(n_3054),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_SL g4008 ( 
.A(n_3639),
.B(n_2856),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3538),
.Y(n_4009)
);

AOI21xp5_ASAP7_75t_L g4010 ( 
.A1(n_3636),
.A2(n_3357),
.B(n_2762),
.Y(n_4010)
);

AOI21xp5_ASAP7_75t_L g4011 ( 
.A1(n_3701),
.A2(n_2762),
.B(n_2755),
.Y(n_4011)
);

OAI21x1_ASAP7_75t_L g4012 ( 
.A1(n_3838),
.A2(n_2148),
.B(n_3171),
.Y(n_4012)
);

AOI21xp5_ASAP7_75t_L g4013 ( 
.A1(n_3854),
.A2(n_2762),
.B(n_2755),
.Y(n_4013)
);

AOI21xp5_ASAP7_75t_L g4014 ( 
.A1(n_3854),
.A2(n_3776),
.B(n_3829),
.Y(n_4014)
);

O2A1O1Ixp33_ASAP7_75t_L g4015 ( 
.A1(n_3830),
.A2(n_840),
.B(n_848),
.C(n_843),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3776),
.A2(n_2907),
.B(n_2798),
.Y(n_4016)
);

O2A1O1Ixp33_ASAP7_75t_L g4017 ( 
.A1(n_3816),
.A2(n_843),
.B(n_849),
.C(n_848),
.Y(n_4017)
);

A2O1A1Ixp33_ASAP7_75t_L g4018 ( 
.A1(n_3848),
.A2(n_3107),
.B(n_2949),
.C(n_3304),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3723),
.B(n_1433),
.Y(n_4019)
);

BUFx3_ASAP7_75t_L g4020 ( 
.A(n_3529),
.Y(n_4020)
);

OAI22xp5_ASAP7_75t_L g4021 ( 
.A1(n_3855),
.A2(n_2916),
.B1(n_2907),
.B2(n_2914),
.Y(n_4021)
);

AOI21x1_ASAP7_75t_L g4022 ( 
.A1(n_3750),
.A2(n_2940),
.B(n_2819),
.Y(n_4022)
);

OAI21x1_ASAP7_75t_L g4023 ( 
.A1(n_3849),
.A2(n_3171),
.B(n_2417),
.Y(n_4023)
);

HB1xp67_ASAP7_75t_L g4024 ( 
.A(n_3605),
.Y(n_4024)
);

AOI21xp5_ASAP7_75t_L g4025 ( 
.A1(n_3546),
.A2(n_2914),
.B(n_2798),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_SL g4026 ( 
.A(n_3639),
.B(n_3717),
.Y(n_4026)
);

NAND3xp33_ASAP7_75t_SL g4027 ( 
.A(n_3832),
.B(n_756),
.C(n_753),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_3621),
.Y(n_4028)
);

OAI22xp5_ASAP7_75t_L g4029 ( 
.A1(n_3855),
.A2(n_2916),
.B1(n_2914),
.B2(n_2798),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_3687),
.B(n_2768),
.Y(n_4030)
);

INVx2_ASAP7_75t_SL g4031 ( 
.A(n_3593),
.Y(n_4031)
);

NOR2xp33_ASAP7_75t_L g4032 ( 
.A(n_3616),
.B(n_3272),
.Y(n_4032)
);

AOI22xp5_ASAP7_75t_L g4033 ( 
.A1(n_3785),
.A2(n_2760),
.B1(n_2831),
.B2(n_2757),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_3633),
.Y(n_4034)
);

NOR2xp33_ASAP7_75t_L g4035 ( 
.A(n_3624),
.B(n_3273),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_L g4036 ( 
.A(n_3760),
.B(n_3762),
.Y(n_4036)
);

AOI21xp5_ASAP7_75t_L g4037 ( 
.A1(n_3548),
.A2(n_2319),
.B(n_2315),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3557),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_3767),
.B(n_2770),
.Y(n_4039)
);

O2A1O1Ixp33_ASAP7_75t_L g4040 ( 
.A1(n_3570),
.A2(n_851),
.B(n_861),
.C(n_849),
.Y(n_4040)
);

O2A1O1Ixp33_ASAP7_75t_L g4041 ( 
.A1(n_3570),
.A2(n_861),
.B(n_863),
.C(n_851),
.Y(n_4041)
);

OAI22xp33_ASAP7_75t_SL g4042 ( 
.A1(n_3765),
.A2(n_872),
.B1(n_879),
.B2(n_863),
.Y(n_4042)
);

NAND2x1p5_ASAP7_75t_L g4043 ( 
.A(n_3755),
.B(n_3421),
.Y(n_4043)
);

O2A1O1Ixp33_ASAP7_75t_L g4044 ( 
.A1(n_3799),
.A2(n_877),
.B(n_879),
.C(n_872),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_3768),
.B(n_2773),
.Y(n_4045)
);

NAND2xp5_ASAP7_75t_L g4046 ( 
.A(n_3794),
.B(n_2776),
.Y(n_4046)
);

AND2x2_ASAP7_75t_L g4047 ( 
.A(n_3799),
.B(n_1434),
.Y(n_4047)
);

OAI221xp5_ASAP7_75t_L g4048 ( 
.A1(n_3645),
.A2(n_2906),
.B1(n_2841),
.B2(n_1365),
.C(n_1367),
.Y(n_4048)
);

AOI21xp5_ASAP7_75t_L g4049 ( 
.A1(n_3548),
.A2(n_3563),
.B(n_3554),
.Y(n_4049)
);

AOI21xp5_ASAP7_75t_L g4050 ( 
.A1(n_3554),
.A2(n_3089),
.B(n_3054),
.Y(n_4050)
);

AND2x4_ASAP7_75t_L g4051 ( 
.A(n_3656),
.B(n_3421),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3806),
.B(n_2778),
.Y(n_4052)
);

NOR2xp33_ASAP7_75t_R g4053 ( 
.A(n_3696),
.B(n_2872),
.Y(n_4053)
);

AOI21xp5_ASAP7_75t_L g4054 ( 
.A1(n_3563),
.A2(n_3089),
.B(n_3107),
.Y(n_4054)
);

INVxp67_ASAP7_75t_L g4055 ( 
.A(n_3661),
.Y(n_4055)
);

AOI21x1_ASAP7_75t_L g4056 ( 
.A1(n_3824),
.A2(n_2532),
.B(n_2733),
.Y(n_4056)
);

BUFx6f_ASAP7_75t_L g4057 ( 
.A(n_3577),
.Y(n_4057)
);

INVx2_ASAP7_75t_SL g4058 ( 
.A(n_3627),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3759),
.B(n_2780),
.Y(n_4059)
);

INVx3_ASAP7_75t_L g4060 ( 
.A(n_3843),
.Y(n_4060)
);

AOI21xp5_ASAP7_75t_L g4061 ( 
.A1(n_3537),
.A2(n_3089),
.B(n_2969),
.Y(n_4061)
);

INVxp67_ASAP7_75t_SL g4062 ( 
.A(n_3813),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3813),
.B(n_2781),
.Y(n_4063)
);

AOI21xp5_ASAP7_75t_L g4064 ( 
.A1(n_3537),
.A2(n_3089),
.B(n_2969),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3850),
.B(n_2786),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_SL g4066 ( 
.A(n_3717),
.B(n_3320),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_SL g4067 ( 
.A(n_3761),
.B(n_3320),
.Y(n_4067)
);

OAI21x1_ASAP7_75t_L g4068 ( 
.A1(n_3831),
.A2(n_2417),
.B(n_2416),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3560),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3687),
.B(n_3765),
.Y(n_4070)
);

OAI22xp5_ASAP7_75t_L g4071 ( 
.A1(n_3645),
.A2(n_3412),
.B1(n_3459),
.B2(n_3434),
.Y(n_4071)
);

A2O1A1Ixp33_ASAP7_75t_SL g4072 ( 
.A1(n_3614),
.A2(n_2791),
.B(n_2792),
.C(n_2789),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_SL g4073 ( 
.A(n_3814),
.B(n_3024),
.Y(n_4073)
);

OR2x6_ASAP7_75t_L g4074 ( 
.A(n_3579),
.B(n_3434),
.Y(n_4074)
);

BUFx6f_ASAP7_75t_L g4075 ( 
.A(n_3577),
.Y(n_4075)
);

AOI22xp33_ASAP7_75t_L g4076 ( 
.A1(n_3782),
.A2(n_3771),
.B1(n_3852),
.B2(n_3785),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_SL g4077 ( 
.A(n_3820),
.B(n_3024),
.Y(n_4077)
);

O2A1O1Ixp5_ASAP7_75t_L g4078 ( 
.A1(n_3819),
.A2(n_3151),
.B(n_3108),
.C(n_2800),
.Y(n_4078)
);

INVx3_ASAP7_75t_L g4079 ( 
.A(n_3542),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3567),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_SL g4081 ( 
.A(n_3820),
.B(n_3024),
.Y(n_4081)
);

AOI22xp5_ASAP7_75t_L g4082 ( 
.A1(n_3771),
.A2(n_3070),
.B1(n_3175),
.B2(n_3177),
.Y(n_4082)
);

A2O1A1Ixp33_ASAP7_75t_L g4083 ( 
.A1(n_3713),
.A2(n_2935),
.B(n_2834),
.C(n_3175),
.Y(n_4083)
);

OAI21xp5_ASAP7_75t_L g4084 ( 
.A1(n_3544),
.A2(n_2804),
.B(n_2793),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_SL g4085 ( 
.A(n_3788),
.B(n_3779),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3857),
.B(n_3779),
.Y(n_4086)
);

A2O1A1Ixp33_ASAP7_75t_L g4087 ( 
.A1(n_3853),
.A2(n_2810),
.B(n_2821),
.C(n_2805),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3635),
.Y(n_4088)
);

AOI22xp5_ASAP7_75t_L g4089 ( 
.A1(n_3798),
.A2(n_3070),
.B1(n_2825),
.B2(n_2769),
.Y(n_4089)
);

OAI22x1_ASAP7_75t_L g4090 ( 
.A1(n_3754),
.A2(n_884),
.B1(n_888),
.B2(n_877),
.Y(n_4090)
);

AOI22xp33_ASAP7_75t_L g4091 ( 
.A1(n_3844),
.A2(n_2849),
.B1(n_2873),
.B2(n_2829),
.Y(n_4091)
);

INVx2_ASAP7_75t_L g4092 ( 
.A(n_3638),
.Y(n_4092)
);

AOI22xp5_ASAP7_75t_L g4093 ( 
.A1(n_3798),
.A2(n_3070),
.B1(n_2825),
.B2(n_2769),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_SL g4094 ( 
.A(n_3752),
.B(n_3031),
.Y(n_4094)
);

INVx3_ASAP7_75t_L g4095 ( 
.A(n_3542),
.Y(n_4095)
);

AOI22xp33_ASAP7_75t_L g4096 ( 
.A1(n_3818),
.A2(n_2863),
.B1(n_2894),
.B2(n_2839),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3817),
.B(n_2824),
.Y(n_4097)
);

CKINVDCx20_ASAP7_75t_R g4098 ( 
.A(n_3680),
.Y(n_4098)
);

BUFx6f_ASAP7_75t_L g4099 ( 
.A(n_3577),
.Y(n_4099)
);

AOI21xp5_ASAP7_75t_L g4100 ( 
.A1(n_3544),
.A2(n_3665),
.B(n_3613),
.Y(n_4100)
);

AOI21xp5_ASAP7_75t_L g4101 ( 
.A1(n_3599),
.A2(n_2969),
.B(n_2967),
.Y(n_4101)
);

A2O1A1Ixp33_ASAP7_75t_L g4102 ( 
.A1(n_3737),
.A2(n_2827),
.B(n_2828),
.C(n_2826),
.Y(n_4102)
);

O2A1O1Ixp33_ASAP7_75t_L g4103 ( 
.A1(n_3790),
.A2(n_3824),
.B(n_3828),
.C(n_3775),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3574),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_L g4105 ( 
.A(n_3823),
.B(n_2833),
.Y(n_4105)
);

HB1xp67_ASAP7_75t_L g4106 ( 
.A(n_3686),
.Y(n_4106)
);

AOI21xp5_ASAP7_75t_L g4107 ( 
.A1(n_3599),
.A2(n_2987),
.B(n_2967),
.Y(n_4107)
);

O2A1O1Ixp5_ASAP7_75t_L g4108 ( 
.A1(n_3828),
.A2(n_3841),
.B(n_3810),
.C(n_3833),
.Y(n_4108)
);

INVx3_ASAP7_75t_L g4109 ( 
.A(n_3542),
.Y(n_4109)
);

OAI22xp5_ASAP7_75t_L g4110 ( 
.A1(n_3796),
.A2(n_3459),
.B1(n_2388),
.B2(n_2390),
.Y(n_4110)
);

AOI21xp5_ASAP7_75t_L g4111 ( 
.A1(n_3613),
.A2(n_2987),
.B(n_2967),
.Y(n_4111)
);

OAI21xp5_ASAP7_75t_L g4112 ( 
.A1(n_3803),
.A2(n_2842),
.B(n_2836),
.Y(n_4112)
);

NOR2xp33_ASAP7_75t_L g4113 ( 
.A(n_3604),
.B(n_767),
.Y(n_4113)
);

NOR2xp33_ASAP7_75t_R g4114 ( 
.A(n_3604),
.B(n_2920),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_3582),
.Y(n_4115)
);

O2A1O1Ixp33_ASAP7_75t_L g4116 ( 
.A1(n_3614),
.A2(n_888),
.B(n_893),
.C(n_884),
.Y(n_4116)
);

OAI22xp5_ASAP7_75t_L g4117 ( 
.A1(n_3796),
.A2(n_2388),
.B1(n_2390),
.B2(n_2382),
.Y(n_4117)
);

INVx2_ASAP7_75t_L g4118 ( 
.A(n_3655),
.Y(n_4118)
);

OR2x6_ASAP7_75t_L g4119 ( 
.A(n_3579),
.B(n_3070),
.Y(n_4119)
);

BUFx6f_ASAP7_75t_L g4120 ( 
.A(n_3586),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_3619),
.B(n_2843),
.Y(n_4121)
);

HB1xp67_ASAP7_75t_L g4122 ( 
.A(n_3722),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_3619),
.B(n_2846),
.Y(n_4123)
);

CKINVDCx20_ASAP7_75t_R g4124 ( 
.A(n_3551),
.Y(n_4124)
);

O2A1O1Ixp33_ASAP7_75t_L g4125 ( 
.A1(n_3609),
.A2(n_899),
.B(n_900),
.C(n_893),
.Y(n_4125)
);

NOR2xp33_ASAP7_75t_L g4126 ( 
.A(n_3752),
.B(n_769),
.Y(n_4126)
);

AOI21xp5_ASAP7_75t_L g4127 ( 
.A1(n_3573),
.A2(n_2994),
.B(n_2987),
.Y(n_4127)
);

NOR2xp33_ASAP7_75t_L g4128 ( 
.A(n_3764),
.B(n_773),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_SL g4129 ( 
.A(n_3764),
.B(n_3818),
.Y(n_4129)
);

AOI21x1_ASAP7_75t_L g4130 ( 
.A1(n_3803),
.A2(n_2612),
.B(n_2607),
.Y(n_4130)
);

NOR2xp33_ASAP7_75t_L g4131 ( 
.A(n_3603),
.B(n_780),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_3597),
.B(n_3774),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_3597),
.B(n_2848),
.Y(n_4133)
);

INVx2_ASAP7_75t_L g4134 ( 
.A(n_3689),
.Y(n_4134)
);

AOI21xp5_ASAP7_75t_L g4135 ( 
.A1(n_3576),
.A2(n_2994),
.B(n_2505),
.Y(n_4135)
);

INVx2_ASAP7_75t_L g4136 ( 
.A(n_3694),
.Y(n_4136)
);

HB1xp67_ASAP7_75t_L g4137 ( 
.A(n_3811),
.Y(n_4137)
);

AOI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_3576),
.A2(n_3571),
.B(n_3729),
.Y(n_4138)
);

OAI22xp5_ASAP7_75t_L g4139 ( 
.A1(n_3702),
.A2(n_2388),
.B1(n_2390),
.B2(n_2382),
.Y(n_4139)
);

AOI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_3729),
.A2(n_2542),
.B(n_2440),
.Y(n_4140)
);

NAND2x1p5_ASAP7_75t_L g4141 ( 
.A(n_3755),
.B(n_3031),
.Y(n_4141)
);

NOR2xp67_ASAP7_75t_SL g4142 ( 
.A(n_3786),
.B(n_3031),
.Y(n_4142)
);

NOR2xp33_ASAP7_75t_L g4143 ( 
.A(n_3603),
.B(n_783),
.Y(n_4143)
);

NOR2xp33_ASAP7_75t_L g4144 ( 
.A(n_3748),
.B(n_784),
.Y(n_4144)
);

AOI21xp5_ASAP7_75t_L g4145 ( 
.A1(n_3643),
.A2(n_2542),
.B(n_2440),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_3721),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_SL g4147 ( 
.A(n_3737),
.B(n_3031),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_3585),
.Y(n_4148)
);

A2O1A1Ixp33_ASAP7_75t_L g4149 ( 
.A1(n_3708),
.A2(n_2858),
.B(n_2866),
.C(n_2850),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_3587),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_3588),
.Y(n_4151)
);

AO32x2_ASAP7_75t_L g4152 ( 
.A1(n_3535),
.A2(n_2794),
.A3(n_1895),
.B1(n_1111),
.B2(n_2267),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_3708),
.B(n_2871),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3709),
.B(n_2877),
.Y(n_4154)
);

OA22x2_ASAP7_75t_L g4155 ( 
.A1(n_3845),
.A2(n_900),
.B1(n_911),
.B2(n_899),
.Y(n_4155)
);

BUFx6f_ASAP7_75t_L g4156 ( 
.A(n_3586),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3594),
.Y(n_4157)
);

AOI22xp5_ASAP7_75t_L g4158 ( 
.A1(n_3704),
.A2(n_2995),
.B1(n_3033),
.B2(n_2992),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3595),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_3664),
.B(n_1435),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3602),
.Y(n_4161)
);

O2A1O1Ixp33_ASAP7_75t_L g4162 ( 
.A1(n_3810),
.A2(n_917),
.B(n_920),
.C(n_911),
.Y(n_4162)
);

NOR2xp33_ASAP7_75t_L g4163 ( 
.A(n_3653),
.B(n_785),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_SL g4164 ( 
.A(n_3667),
.B(n_3058),
.Y(n_4164)
);

INVx5_ASAP7_75t_L g4165 ( 
.A(n_3566),
.Y(n_4165)
);

BUFx6f_ASAP7_75t_L g4166 ( 
.A(n_3586),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_3733),
.B(n_2886),
.Y(n_4167)
);

OR2x2_ASAP7_75t_SL g4168 ( 
.A(n_3541),
.B(n_917),
.Y(n_4168)
);

NOR2xp33_ASAP7_75t_R g4169 ( 
.A(n_3611),
.B(n_2920),
.Y(n_4169)
);

BUFx3_ASAP7_75t_L g4170 ( 
.A(n_3712),
.Y(n_4170)
);

AOI21xp5_ASAP7_75t_L g4171 ( 
.A1(n_3658),
.A2(n_3674),
.B(n_3659),
.Y(n_4171)
);

AOI22xp5_ASAP7_75t_L g4172 ( 
.A1(n_3704),
.A2(n_2995),
.B1(n_3033),
.B2(n_2992),
.Y(n_4172)
);

NOR2xp33_ASAP7_75t_L g4173 ( 
.A(n_3664),
.B(n_786),
.Y(n_4173)
);

INVx3_ASAP7_75t_L g4174 ( 
.A(n_3579),
.Y(n_4174)
);

BUFx12f_ASAP7_75t_L g4175 ( 
.A(n_3611),
.Y(n_4175)
);

CKINVDCx11_ASAP7_75t_R g4176 ( 
.A(n_3793),
.Y(n_4176)
);

AOI21xp5_ASAP7_75t_L g4177 ( 
.A1(n_3658),
.A2(n_2572),
.B(n_2542),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_SL g4178 ( 
.A(n_3702),
.B(n_3063),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_3606),
.Y(n_4179)
);

INVx2_ASAP7_75t_L g4180 ( 
.A(n_3725),
.Y(n_4180)
);

OR2x6_ASAP7_75t_L g4181 ( 
.A(n_3580),
.B(n_3058),
.Y(n_4181)
);

BUFx6f_ASAP7_75t_L g4182 ( 
.A(n_3651),
.Y(n_4182)
);

OAI22x1_ASAP7_75t_L g4183 ( 
.A1(n_3608),
.A2(n_923),
.B1(n_925),
.B2(n_920),
.Y(n_4183)
);

AOI22xp5_ASAP7_75t_L g4184 ( 
.A1(n_3536),
.A2(n_3678),
.B1(n_3690),
.B2(n_3674),
.Y(n_4184)
);

OAI22xp5_ASAP7_75t_L g4185 ( 
.A1(n_3781),
.A2(n_2396),
.B1(n_2374),
.B2(n_2376),
.Y(n_4185)
);

AO21x1_ASAP7_75t_L g4186 ( 
.A1(n_3833),
.A2(n_2905),
.B(n_2897),
.Y(n_4186)
);

INVx2_ASAP7_75t_L g4187 ( 
.A(n_3530),
.Y(n_4187)
);

AOI21xp5_ASAP7_75t_L g4188 ( 
.A1(n_3678),
.A2(n_2572),
.B(n_2542),
.Y(n_4188)
);

BUFx6f_ASAP7_75t_L g4189 ( 
.A(n_3651),
.Y(n_4189)
);

AOI21xp5_ASAP7_75t_L g4190 ( 
.A1(n_3690),
.A2(n_2572),
.B(n_2542),
.Y(n_4190)
);

NOR2xp33_ASAP7_75t_L g4191 ( 
.A(n_3769),
.B(n_788),
.Y(n_4191)
);

NAND3xp33_ASAP7_75t_L g4192 ( 
.A(n_3675),
.B(n_794),
.C(n_791),
.Y(n_4192)
);

AND2x2_ASAP7_75t_L g4193 ( 
.A(n_3532),
.B(n_1436),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_SL g4194 ( 
.A(n_3781),
.B(n_3795),
.Y(n_4194)
);

AND2x2_ASAP7_75t_L g4195 ( 
.A(n_3543),
.B(n_1437),
.Y(n_4195)
);

A2O1A1Ixp33_ASAP7_75t_L g4196 ( 
.A1(n_3732),
.A2(n_2913),
.B(n_2918),
.C(n_2908),
.Y(n_4196)
);

AOI21x1_ASAP7_75t_L g4197 ( 
.A1(n_3851),
.A2(n_2927),
.B(n_2922),
.Y(n_4197)
);

BUFx5_ASAP7_75t_L g4198 ( 
.A(n_3975),
.Y(n_4198)
);

AOI22xp5_ASAP7_75t_L g4199 ( 
.A1(n_3878),
.A2(n_3649),
.B1(n_3623),
.B2(n_3732),
.Y(n_4199)
);

AOI22xp5_ASAP7_75t_L g4200 ( 
.A1(n_3994),
.A2(n_3649),
.B1(n_3746),
.B2(n_3744),
.Y(n_4200)
);

AOI21xp5_ASAP7_75t_L g4201 ( 
.A1(n_3862),
.A2(n_3851),
.B(n_3795),
.Y(n_4201)
);

BUFx6f_ASAP7_75t_L g4202 ( 
.A(n_4176),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4009),
.Y(n_4203)
);

OR2x6_ASAP7_75t_SL g4204 ( 
.A(n_3902),
.B(n_799),
.Y(n_4204)
);

NAND2x1_ASAP7_75t_L g4205 ( 
.A(n_4142),
.B(n_3575),
.Y(n_4205)
);

AOI22xp5_ASAP7_75t_L g4206 ( 
.A1(n_3892),
.A2(n_3778),
.B1(n_3751),
.B2(n_803),
.Y(n_4206)
);

BUFx6f_ASAP7_75t_L g4207 ( 
.A(n_3959),
.Y(n_4207)
);

OR2x2_ASAP7_75t_L g4208 ( 
.A(n_3877),
.B(n_3876),
.Y(n_4208)
);

AOI21xp5_ASAP7_75t_L g4209 ( 
.A1(n_4171),
.A2(n_3778),
.B(n_2794),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_4038),
.Y(n_4210)
);

OAI22xp5_ASAP7_75t_L g4211 ( 
.A1(n_4070),
.A2(n_3699),
.B1(n_3675),
.B2(n_3617),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_3881),
.Y(n_4212)
);

INVx2_ASAP7_75t_L g4213 ( 
.A(n_3888),
.Y(n_4213)
);

NAND2x1_ASAP7_75t_SL g4214 ( 
.A(n_3866),
.B(n_3996),
.Y(n_4214)
);

BUFx6f_ASAP7_75t_L g4215 ( 
.A(n_3959),
.Y(n_4215)
);

BUFx3_ASAP7_75t_L g4216 ( 
.A(n_4020),
.Y(n_4216)
);

OAI22xp33_ASAP7_75t_L g4217 ( 
.A1(n_3871),
.A2(n_3622),
.B1(n_3629),
.B2(n_3610),
.Y(n_4217)
);

NAND3xp33_ASAP7_75t_L g4218 ( 
.A(n_3910),
.B(n_804),
.C(n_802),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_3930),
.Y(n_4219)
);

BUFx3_ASAP7_75t_L g4220 ( 
.A(n_4170),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_4069),
.Y(n_4221)
);

NOR2x1_ASAP7_75t_R g4222 ( 
.A(n_4175),
.B(n_3786),
.Y(n_4222)
);

INVx3_ASAP7_75t_L g4223 ( 
.A(n_3996),
.Y(n_4223)
);

AND2x4_ASAP7_75t_L g4224 ( 
.A(n_4079),
.B(n_3836),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_4070),
.B(n_3634),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4080),
.Y(n_4226)
);

CKINVDCx20_ASAP7_75t_R g4227 ( 
.A(n_4098),
.Y(n_4227)
);

BUFx6f_ASAP7_75t_L g4228 ( 
.A(n_3959),
.Y(n_4228)
);

AOI22xp33_ASAP7_75t_L g4229 ( 
.A1(n_4027),
.A2(n_925),
.B1(n_927),
.B2(n_923),
.Y(n_4229)
);

INVx4_ASAP7_75t_L g4230 ( 
.A(n_3991),
.Y(n_4230)
);

BUFx6f_ASAP7_75t_L g4231 ( 
.A(n_3991),
.Y(n_4231)
);

AO21x2_ASAP7_75t_L g4232 ( 
.A1(n_4000),
.A2(n_3640),
.B(n_3637),
.Y(n_4232)
);

INVx3_ASAP7_75t_L g4233 ( 
.A(n_4005),
.Y(n_4233)
);

INVx3_ASAP7_75t_L g4234 ( 
.A(n_4005),
.Y(n_4234)
);

O2A1O1Ixp33_ASAP7_75t_SL g4235 ( 
.A1(n_4072),
.A2(n_932),
.B(n_934),
.C(n_927),
.Y(n_4235)
);

INVx2_ASAP7_75t_SL g4236 ( 
.A(n_3962),
.Y(n_4236)
);

BUFx6f_ASAP7_75t_L g4237 ( 
.A(n_3872),
.Y(n_4237)
);

INVx3_ASAP7_75t_L g4238 ( 
.A(n_4060),
.Y(n_4238)
);

BUFx6f_ASAP7_75t_L g4239 ( 
.A(n_3872),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4104),
.Y(n_4240)
);

BUFx6f_ASAP7_75t_L g4241 ( 
.A(n_3872),
.Y(n_4241)
);

AOI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_3972),
.A2(n_3699),
.B(n_2462),
.Y(n_4242)
);

INVx5_ASAP7_75t_L g4243 ( 
.A(n_4119),
.Y(n_4243)
);

BUFx4f_ASAP7_75t_SL g4244 ( 
.A(n_3939),
.Y(n_4244)
);

AOI22xp5_ASAP7_75t_L g4245 ( 
.A1(n_3929),
.A2(n_812),
.B1(n_814),
.B2(n_810),
.Y(n_4245)
);

INVx1_ASAP7_75t_SL g4246 ( 
.A(n_3981),
.Y(n_4246)
);

INVx2_ASAP7_75t_SL g4247 ( 
.A(n_3962),
.Y(n_4247)
);

AOI21xp5_ASAP7_75t_L g4248 ( 
.A1(n_4101),
.A2(n_2462),
.B(n_2456),
.Y(n_4248)
);

AND2x4_ASAP7_75t_L g4249 ( 
.A(n_4079),
.B(n_3580),
.Y(n_4249)
);

O2A1O1Ixp33_ASAP7_75t_L g4250 ( 
.A1(n_3887),
.A2(n_1014),
.B(n_1022),
.C(n_935),
.Y(n_4250)
);

OR2x6_ASAP7_75t_L g4251 ( 
.A(n_4014),
.B(n_3580),
.Y(n_4251)
);

OR2x6_ASAP7_75t_L g4252 ( 
.A(n_4007),
.B(n_3583),
.Y(n_4252)
);

CKINVDCx11_ASAP7_75t_R g4253 ( 
.A(n_3983),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_4085),
.B(n_4132),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4115),
.Y(n_4255)
);

OAI22xp5_ASAP7_75t_L g4256 ( 
.A1(n_3916),
.A2(n_3644),
.B1(n_3646),
.B2(n_3641),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_4049),
.B(n_3647),
.Y(n_4257)
);

INVx4_ASAP7_75t_L g4258 ( 
.A(n_3908),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4148),
.Y(n_4259)
);

AND2x2_ASAP7_75t_L g4260 ( 
.A(n_3999),
.B(n_3648),
.Y(n_4260)
);

OAI21xp33_ASAP7_75t_L g4261 ( 
.A1(n_3865),
.A2(n_4184),
.B(n_3964),
.Y(n_4261)
);

INVxp67_ASAP7_75t_SL g4262 ( 
.A(n_4186),
.Y(n_4262)
);

OAI221xp5_ASAP7_75t_L g4263 ( 
.A1(n_3974),
.A2(n_3941),
.B1(n_4015),
.B2(n_3985),
.C(n_3982),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_SL g4264 ( 
.A(n_4026),
.B(n_3786),
.Y(n_4264)
);

OAI22xp5_ASAP7_75t_L g4265 ( 
.A1(n_4168),
.A2(n_3670),
.B1(n_3671),
.B2(n_3662),
.Y(n_4265)
);

CKINVDCx5p33_ASAP7_75t_R g4266 ( 
.A(n_3943),
.Y(n_4266)
);

NOR2xp67_ASAP7_75t_SL g4267 ( 
.A(n_3859),
.B(n_3575),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4150),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_4086),
.B(n_3679),
.Y(n_4269)
);

BUFx2_ASAP7_75t_L g4270 ( 
.A(n_3899),
.Y(n_4270)
);

OR2x6_ASAP7_75t_L g4271 ( 
.A(n_4007),
.B(n_3915),
.Y(n_4271)
);

INVxp67_ASAP7_75t_SL g4272 ( 
.A(n_4062),
.Y(n_4272)
);

O2A1O1Ixp33_ASAP7_75t_SL g4273 ( 
.A1(n_3891),
.A2(n_943),
.B(n_944),
.C(n_938),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4151),
.Y(n_4274)
);

INVx3_ASAP7_75t_L g4275 ( 
.A(n_4060),
.Y(n_4275)
);

INVx2_ASAP7_75t_L g4276 ( 
.A(n_4028),
.Y(n_4276)
);

AND2x4_ASAP7_75t_L g4277 ( 
.A(n_4095),
.B(n_4109),
.Y(n_4277)
);

NOR2x1_ASAP7_75t_L g4278 ( 
.A(n_3864),
.B(n_3618),
.Y(n_4278)
);

INVx2_ASAP7_75t_L g4279 ( 
.A(n_4034),
.Y(n_4279)
);

CKINVDCx20_ASAP7_75t_R g4280 ( 
.A(n_4124),
.Y(n_4280)
);

BUFx2_ASAP7_75t_L g4281 ( 
.A(n_4024),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4157),
.Y(n_4282)
);

NOR2xp33_ASAP7_75t_L g4283 ( 
.A(n_3860),
.B(n_3681),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4159),
.Y(n_4284)
);

AOI22xp33_ASAP7_75t_L g4285 ( 
.A1(n_3898),
.A2(n_943),
.B1(n_944),
.B2(n_938),
.Y(n_4285)
);

AND2x4_ASAP7_75t_L g4286 ( 
.A(n_4095),
.B(n_3583),
.Y(n_4286)
);

OR2x2_ASAP7_75t_L g4287 ( 
.A(n_3921),
.B(n_3682),
.Y(n_4287)
);

AND2x2_ASAP7_75t_L g4288 ( 
.A(n_3931),
.B(n_3685),
.Y(n_4288)
);

AO22x2_ASAP7_75t_L g4289 ( 
.A1(n_3952),
.A2(n_3695),
.B1(n_3698),
.B2(n_3688),
.Y(n_4289)
);

INVx3_ASAP7_75t_L g4290 ( 
.A(n_4057),
.Y(n_4290)
);

INVx3_ASAP7_75t_L g4291 ( 
.A(n_4057),
.Y(n_4291)
);

A2O1A1Ixp33_ASAP7_75t_L g4292 ( 
.A1(n_3868),
.A2(n_953),
.B(n_958),
.C(n_946),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4161),
.Y(n_4293)
);

OR2x6_ASAP7_75t_L g4294 ( 
.A(n_4007),
.B(n_3583),
.Y(n_4294)
);

BUFx6f_ASAP7_75t_L g4295 ( 
.A(n_3926),
.Y(n_4295)
);

AND2x4_ASAP7_75t_L g4296 ( 
.A(n_4109),
.B(n_3589),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4179),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4106),
.Y(n_4298)
);

BUFx12f_ASAP7_75t_L g4299 ( 
.A(n_3926),
.Y(n_4299)
);

INVx1_ASAP7_75t_SL g4300 ( 
.A(n_3981),
.Y(n_4300)
);

AND2x2_ASAP7_75t_L g4301 ( 
.A(n_4019),
.B(n_3700),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4122),
.Y(n_4302)
);

INVx3_ASAP7_75t_L g4303 ( 
.A(n_4075),
.Y(n_4303)
);

INVx3_ASAP7_75t_L g4304 ( 
.A(n_4075),
.Y(n_4304)
);

BUFx4f_ASAP7_75t_L g4305 ( 
.A(n_3926),
.Y(n_4305)
);

INVx2_ASAP7_75t_SL g4306 ( 
.A(n_4058),
.Y(n_4306)
);

INVx2_ASAP7_75t_L g4307 ( 
.A(n_4088),
.Y(n_4307)
);

INVx4_ASAP7_75t_L g4308 ( 
.A(n_3938),
.Y(n_4308)
);

CKINVDCx5p33_ASAP7_75t_R g4309 ( 
.A(n_3883),
.Y(n_4309)
);

AOI21xp33_ASAP7_75t_L g4310 ( 
.A1(n_4162),
.A2(n_2941),
.B(n_2938),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4194),
.B(n_3531),
.Y(n_4311)
);

INVxp67_ASAP7_75t_L g4312 ( 
.A(n_3976),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_4138),
.B(n_3531),
.Y(n_4313)
);

AOI21xp5_ASAP7_75t_L g4314 ( 
.A1(n_4107),
.A2(n_2462),
.B(n_2456),
.Y(n_4314)
);

BUFx4f_ASAP7_75t_L g4315 ( 
.A(n_3938),
.Y(n_4315)
);

INVx5_ASAP7_75t_L g4316 ( 
.A(n_4119),
.Y(n_4316)
);

NAND2x1_ASAP7_75t_L g4317 ( 
.A(n_4074),
.B(n_3618),
.Y(n_4317)
);

AOI22xp5_ASAP7_75t_L g4318 ( 
.A1(n_3896),
.A2(n_819),
.B1(n_820),
.B2(n_816),
.Y(n_4318)
);

OAI221xp5_ASAP7_75t_L g4319 ( 
.A1(n_4192),
.A2(n_958),
.B1(n_967),
.B2(n_953),
.C(n_946),
.Y(n_4319)
);

INVx3_ASAP7_75t_L g4320 ( 
.A(n_4075),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_4092),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_3858),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_L g4323 ( 
.A(n_4100),
.B(n_3569),
.Y(n_4323)
);

INVx2_ASAP7_75t_L g4324 ( 
.A(n_4118),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_3977),
.B(n_3569),
.Y(n_4325)
);

NAND2x1_ASAP7_75t_SL g4326 ( 
.A(n_3905),
.B(n_4137),
.Y(n_4326)
);

INVx5_ASAP7_75t_SL g4327 ( 
.A(n_4181),
.Y(n_4327)
);

INVx2_ASAP7_75t_SL g4328 ( 
.A(n_4031),
.Y(n_4328)
);

OR2x2_ASAP7_75t_L g4329 ( 
.A(n_3912),
.B(n_3630),
.Y(n_4329)
);

INVx3_ASAP7_75t_L g4330 ( 
.A(n_4099),
.Y(n_4330)
);

AOI22xp5_ASAP7_75t_L g4331 ( 
.A1(n_4144),
.A2(n_825),
.B1(n_830),
.B2(n_823),
.Y(n_4331)
);

OAI22xp5_ASAP7_75t_L g4332 ( 
.A1(n_3861),
.A2(n_3589),
.B1(n_3592),
.B2(n_3559),
.Y(n_4332)
);

NAND2x1p5_ASAP7_75t_L g4333 ( 
.A(n_4174),
.B(n_3743),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_3880),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_3977),
.B(n_3980),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_3913),
.Y(n_4336)
);

INVx4_ASAP7_75t_L g4337 ( 
.A(n_3859),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_3932),
.Y(n_4338)
);

AND2x4_ASAP7_75t_L g4339 ( 
.A(n_4119),
.B(n_3589),
.Y(n_4339)
);

BUFx6f_ASAP7_75t_L g4340 ( 
.A(n_4099),
.Y(n_4340)
);

AOI21xp5_ASAP7_75t_SL g4341 ( 
.A1(n_3973),
.A2(n_3592),
.B(n_3615),
.Y(n_4341)
);

AOI22xp5_ASAP7_75t_L g4342 ( 
.A1(n_3897),
.A2(n_3889),
.B1(n_3955),
.B2(n_4113),
.Y(n_4342)
);

INVx4_ASAP7_75t_L g4343 ( 
.A(n_3859),
.Y(n_4343)
);

BUFx8_ASAP7_75t_L g4344 ( 
.A(n_3935),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_3980),
.B(n_3630),
.Y(n_4345)
);

INVx3_ASAP7_75t_L g4346 ( 
.A(n_4099),
.Y(n_4346)
);

CKINVDCx8_ASAP7_75t_R g4347 ( 
.A(n_4120),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_4160),
.B(n_3651),
.Y(n_4348)
);

INVx1_ASAP7_75t_SL g4349 ( 
.A(n_3966),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_L g4350 ( 
.A(n_3911),
.B(n_3652),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_4134),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_L g4352 ( 
.A(n_4036),
.B(n_3652),
.Y(n_4352)
);

OR2x6_ASAP7_75t_L g4353 ( 
.A(n_3915),
.B(n_3592),
.Y(n_4353)
);

INVxp67_ASAP7_75t_L g4354 ( 
.A(n_3925),
.Y(n_4354)
);

AND2x4_ASAP7_75t_L g4355 ( 
.A(n_3915),
.B(n_3793),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_3947),
.Y(n_4356)
);

INVx3_ASAP7_75t_L g4357 ( 
.A(n_4120),
.Y(n_4357)
);

INVx3_ASAP7_75t_L g4358 ( 
.A(n_4120),
.Y(n_4358)
);

INVx2_ASAP7_75t_L g4359 ( 
.A(n_4136),
.Y(n_4359)
);

BUFx3_ASAP7_75t_L g4360 ( 
.A(n_4003),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_3885),
.B(n_3654),
.Y(n_4361)
);

AND2x4_ASAP7_75t_L g4362 ( 
.A(n_4051),
.B(n_4074),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4146),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4180),
.Y(n_4364)
);

CKINVDCx8_ASAP7_75t_R g4365 ( 
.A(n_4156),
.Y(n_4365)
);

OAI21x1_ASAP7_75t_SL g4366 ( 
.A1(n_4103),
.A2(n_3787),
.B(n_2945),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_4187),
.Y(n_4367)
);

NAND2x1p5_ASAP7_75t_L g4368 ( 
.A(n_3859),
.B(n_3559),
.Y(n_4368)
);

INVx2_ASAP7_75t_SL g4369 ( 
.A(n_4156),
.Y(n_4369)
);

AND3x2_ASAP7_75t_L g4370 ( 
.A(n_3953),
.B(n_968),
.C(n_967),
.Y(n_4370)
);

CKINVDCx5p33_ASAP7_75t_R g4371 ( 
.A(n_4053),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_L g4372 ( 
.A(n_3886),
.B(n_3654),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_3937),
.B(n_3657),
.Y(n_4373)
);

INVx2_ASAP7_75t_SL g4374 ( 
.A(n_4156),
.Y(n_4374)
);

BUFx3_ASAP7_75t_L g4375 ( 
.A(n_3927),
.Y(n_4375)
);

NOR2xp33_ASAP7_75t_L g4376 ( 
.A(n_3919),
.B(n_3657),
.Y(n_4376)
);

AOI22xp33_ASAP7_75t_L g4377 ( 
.A1(n_4042),
.A2(n_969),
.B1(n_977),
.B2(n_968),
.Y(n_4377)
);

HB1xp67_ASAP7_75t_L g4378 ( 
.A(n_3914),
.Y(n_4378)
);

OR2x6_ASAP7_75t_L g4379 ( 
.A(n_4050),
.B(n_3615),
.Y(n_4379)
);

BUFx2_ASAP7_75t_L g4380 ( 
.A(n_4114),
.Y(n_4380)
);

AOI21xp5_ASAP7_75t_L g4381 ( 
.A1(n_4111),
.A2(n_2467),
.B(n_2456),
.Y(n_4381)
);

NOR2xp33_ASAP7_75t_L g4382 ( 
.A(n_3924),
.B(n_3719),
.Y(n_4382)
);

INVx2_ASAP7_75t_SL g4383 ( 
.A(n_4166),
.Y(n_4383)
);

BUFx3_ASAP7_75t_L g4384 ( 
.A(n_3927),
.Y(n_4384)
);

INVx2_ASAP7_75t_L g4385 ( 
.A(n_4193),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_4195),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4167),
.Y(n_4387)
);

INVx2_ASAP7_75t_L g4388 ( 
.A(n_3971),
.Y(n_4388)
);

OR2x6_ASAP7_75t_L g4389 ( 
.A(n_4074),
.B(n_3719),
.Y(n_4389)
);

NOR2xp33_ASAP7_75t_L g4390 ( 
.A(n_4055),
.B(n_3953),
.Y(n_4390)
);

OAI21xp5_ASAP7_75t_L g4391 ( 
.A1(n_3893),
.A2(n_2948),
.B(n_2943),
.Y(n_4391)
);

OR2x2_ASAP7_75t_L g4392 ( 
.A(n_3861),
.B(n_3727),
.Y(n_4392)
);

OA21x2_ASAP7_75t_L g4393 ( 
.A1(n_3914),
.A2(n_2376),
.B(n_2374),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4063),
.Y(n_4394)
);

A2O1A1Ixp33_ASAP7_75t_L g4395 ( 
.A1(n_3901),
.A2(n_977),
.B(n_979),
.C(n_969),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_L g4396 ( 
.A(n_3884),
.B(n_3727),
.Y(n_4396)
);

INVx2_ASAP7_75t_L g4397 ( 
.A(n_4059),
.Y(n_4397)
);

AO21x2_ASAP7_75t_L g4398 ( 
.A1(n_3903),
.A2(n_2442),
.B(n_3108),
.Y(n_4398)
);

NAND2xp33_ASAP7_75t_L g4399 ( 
.A(n_4169),
.B(n_3793),
.Y(n_4399)
);

INVx2_ASAP7_75t_SL g4400 ( 
.A(n_4166),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4108),
.Y(n_4401)
);

HAxp5_ASAP7_75t_L g4402 ( 
.A(n_3936),
.B(n_831),
.CON(n_4402),
.SN(n_4402)
);

NOR2xp33_ASAP7_75t_L g4403 ( 
.A(n_3906),
.B(n_3753),
.Y(n_4403)
);

BUFx2_ASAP7_75t_L g4404 ( 
.A(n_4182),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4197),
.Y(n_4405)
);

AND2x4_ASAP7_75t_L g4406 ( 
.A(n_4051),
.B(n_3666),
.Y(n_4406)
);

NOR2xp67_ASAP7_75t_SL g4407 ( 
.A(n_4165),
.B(n_3559),
.Y(n_4407)
);

INVx2_ASAP7_75t_L g4408 ( 
.A(n_4046),
.Y(n_4408)
);

NOR2xp33_ASAP7_75t_L g4409 ( 
.A(n_3940),
.B(n_3753),
.Y(n_4409)
);

AOI22xp33_ASAP7_75t_SL g4410 ( 
.A1(n_3884),
.A2(n_980),
.B1(n_988),
.B2(n_979),
.Y(n_4410)
);

OAI221xp5_ASAP7_75t_L g4411 ( 
.A1(n_4017),
.A2(n_4044),
.B1(n_3904),
.B2(n_4033),
.C(n_3922),
.Y(n_4411)
);

CKINVDCx8_ASAP7_75t_R g4412 ( 
.A(n_4182),
.Y(n_4412)
);

BUFx4_ASAP7_75t_SL g4413 ( 
.A(n_4181),
.Y(n_4413)
);

INVx2_ASAP7_75t_SL g4414 ( 
.A(n_4182),
.Y(n_4414)
);

AND2x4_ASAP7_75t_L g4415 ( 
.A(n_4077),
.B(n_3666),
.Y(n_4415)
);

INVx2_ASAP7_75t_L g4416 ( 
.A(n_4052),
.Y(n_4416)
);

NAND2xp5_ASAP7_75t_L g4417 ( 
.A(n_4030),
.B(n_3728),
.Y(n_4417)
);

BUFx12f_ASAP7_75t_L g4418 ( 
.A(n_3998),
.Y(n_4418)
);

INVx2_ASAP7_75t_L g4419 ( 
.A(n_3990),
.Y(n_4419)
);

CKINVDCx11_ASAP7_75t_R g4420 ( 
.A(n_4189),
.Y(n_4420)
);

BUFx6f_ASAP7_75t_L g4421 ( 
.A(n_4189),
.Y(n_4421)
);

NAND2xp33_ASAP7_75t_L g4422 ( 
.A(n_3890),
.B(n_2923),
.Y(n_4422)
);

OAI22xp5_ASAP7_75t_L g4423 ( 
.A1(n_3923),
.A2(n_3942),
.B1(n_4155),
.B2(n_4076),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4065),
.Y(n_4424)
);

AOI22xp33_ASAP7_75t_SL g4425 ( 
.A1(n_4155),
.A2(n_988),
.B1(n_989),
.B2(n_980),
.Y(n_4425)
);

AND2x2_ASAP7_75t_L g4426 ( 
.A(n_4047),
.B(n_3666),
.Y(n_4426)
);

INVx6_ASAP7_75t_L g4427 ( 
.A(n_4165),
.Y(n_4427)
);

OAI21xp33_ASAP7_75t_L g4428 ( 
.A1(n_4191),
.A2(n_836),
.B(n_835),
.Y(n_4428)
);

INVx2_ASAP7_75t_L g4429 ( 
.A(n_3882),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_L g4430 ( 
.A(n_4030),
.B(n_3728),
.Y(n_4430)
);

INVx1_ASAP7_75t_SL g4431 ( 
.A(n_3944),
.Y(n_4431)
);

O2A1O1Ixp33_ASAP7_75t_L g4432 ( 
.A1(n_3969),
.A2(n_1006),
.B(n_1032),
.C(n_995),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_3882),
.Y(n_4433)
);

INVx3_ASAP7_75t_L g4434 ( 
.A(n_3900),
.Y(n_4434)
);

NOR2xp33_ASAP7_75t_L g4435 ( 
.A(n_4032),
.B(n_3763),
.Y(n_4435)
);

OAI21xp5_ASAP7_75t_L g4436 ( 
.A1(n_4018),
.A2(n_3151),
.B(n_2576),
.Y(n_4436)
);

BUFx3_ASAP7_75t_L g4437 ( 
.A(n_3965),
.Y(n_4437)
);

AOI21xp5_ASAP7_75t_L g4438 ( 
.A1(n_3874),
.A2(n_2471),
.B(n_2467),
.Y(n_4438)
);

INVx2_ASAP7_75t_L g4439 ( 
.A(n_3900),
.Y(n_4439)
);

BUFx6f_ASAP7_75t_L g4440 ( 
.A(n_3869),
.Y(n_4440)
);

AND2x4_ASAP7_75t_L g4441 ( 
.A(n_4081),
.B(n_3669),
.Y(n_4441)
);

BUFx2_ASAP7_75t_L g4442 ( 
.A(n_3909),
.Y(n_4442)
);

BUFx3_ASAP7_75t_L g4443 ( 
.A(n_3978),
.Y(n_4443)
);

NOR2xp33_ASAP7_75t_L g4444 ( 
.A(n_4035),
.B(n_3763),
.Y(n_4444)
);

INVx3_ASAP7_75t_L g4445 ( 
.A(n_3869),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4008),
.Y(n_4446)
);

BUFx2_ASAP7_75t_L g4447 ( 
.A(n_3909),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_3933),
.Y(n_4448)
);

O2A1O1Ixp33_ASAP7_75t_L g4449 ( 
.A1(n_3993),
.A2(n_1006),
.B(n_1032),
.C(n_995),
.Y(n_4449)
);

INVx2_ASAP7_75t_L g4450 ( 
.A(n_4097),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_4105),
.Y(n_4451)
);

HB1xp67_ASAP7_75t_L g4452 ( 
.A(n_3948),
.Y(n_4452)
);

BUFx3_ASAP7_75t_L g4453 ( 
.A(n_3986),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_4121),
.B(n_3783),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_L g4455 ( 
.A(n_4121),
.B(n_3804),
.Y(n_4455)
);

BUFx6f_ASAP7_75t_L g4456 ( 
.A(n_3875),
.Y(n_4456)
);

NOR2xp33_ASAP7_75t_SL g4457 ( 
.A(n_3987),
.B(n_3559),
.Y(n_4457)
);

AND2x4_ASAP7_75t_L g4458 ( 
.A(n_4181),
.B(n_3669),
.Y(n_4458)
);

INVx2_ASAP7_75t_L g4459 ( 
.A(n_3956),
.Y(n_4459)
);

BUFx6f_ASAP7_75t_L g4460 ( 
.A(n_3875),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_L g4461 ( 
.A(n_4123),
.B(n_3804),
.Y(n_4461)
);

NOR2xp33_ASAP7_75t_L g4462 ( 
.A(n_4129),
.B(n_3787),
.Y(n_4462)
);

INVx2_ASAP7_75t_L g4463 ( 
.A(n_3967),
.Y(n_4463)
);

INVx2_ASAP7_75t_SL g4464 ( 
.A(n_3963),
.Y(n_4464)
);

INVx2_ASAP7_75t_SL g4465 ( 
.A(n_3995),
.Y(n_4465)
);

INVx2_ASAP7_75t_L g4466 ( 
.A(n_4004),
.Y(n_4466)
);

INVx5_ASAP7_75t_L g4467 ( 
.A(n_3987),
.Y(n_4467)
);

NOR2x1_ASAP7_75t_L g4468 ( 
.A(n_4164),
.B(n_3736),
.Y(n_4468)
);

AOI21xp5_ASAP7_75t_L g4469 ( 
.A1(n_3894),
.A2(n_2471),
.B(n_2467),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4039),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4045),
.Y(n_4471)
);

AND2x2_ASAP7_75t_L g4472 ( 
.A(n_4126),
.B(n_3673),
.Y(n_4472)
);

CKINVDCx20_ASAP7_75t_R g4473 ( 
.A(n_4128),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_3954),
.Y(n_4474)
);

BUFx10_ASAP7_75t_L g4475 ( 
.A(n_4163),
.Y(n_4475)
);

AOI21xp5_ASAP7_75t_L g4476 ( 
.A1(n_3970),
.A2(n_2471),
.B(n_2683),
.Y(n_4476)
);

BUFx10_ASAP7_75t_L g4477 ( 
.A(n_3979),
.Y(n_4477)
);

AOI21x1_ASAP7_75t_L g4478 ( 
.A1(n_4056),
.A2(n_2376),
.B(n_2396),
.Y(n_4478)
);

BUFx2_ASAP7_75t_L g4479 ( 
.A(n_4141),
.Y(n_4479)
);

NOR2x1p5_ASAP7_75t_L g4480 ( 
.A(n_3946),
.B(n_3673),
.Y(n_4480)
);

OR2x6_ASAP7_75t_L g4481 ( 
.A(n_3870),
.B(n_3673),
.Y(n_4481)
);

INVx2_ASAP7_75t_L g4482 ( 
.A(n_4023),
.Y(n_4482)
);

BUFx3_ASAP7_75t_L g4483 ( 
.A(n_4173),
.Y(n_4483)
);

BUFx8_ASAP7_75t_L g4484 ( 
.A(n_4152),
.Y(n_4484)
);

NOR2xp33_ASAP7_75t_L g4485 ( 
.A(n_4001),
.B(n_3706),
.Y(n_4485)
);

BUFx6f_ASAP7_75t_L g4486 ( 
.A(n_4165),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4112),
.Y(n_4487)
);

INVx2_ASAP7_75t_L g4488 ( 
.A(n_3895),
.Y(n_4488)
);

OAI21x1_ASAP7_75t_L g4489 ( 
.A1(n_3907),
.A2(n_2417),
.B(n_2416),
.Y(n_4489)
);

CKINVDCx5p33_ASAP7_75t_R g4490 ( 
.A(n_4131),
.Y(n_4490)
);

AOI22xp33_ASAP7_75t_L g4491 ( 
.A1(n_4183),
.A2(n_993),
.B1(n_1000),
.B2(n_989),
.Y(n_4491)
);

INVx2_ASAP7_75t_L g4492 ( 
.A(n_4022),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4112),
.Y(n_4493)
);

BUFx3_ASAP7_75t_L g4494 ( 
.A(n_4143),
.Y(n_4494)
);

BUFx8_ASAP7_75t_SL g4495 ( 
.A(n_4133),
.Y(n_4495)
);

NOR2xp33_ASAP7_75t_L g4496 ( 
.A(n_4094),
.B(n_3706),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_3957),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_4123),
.B(n_3697),
.Y(n_4498)
);

AND2x4_ASAP7_75t_L g4499 ( 
.A(n_4147),
.B(n_3707),
.Y(n_4499)
);

INVxp67_ASAP7_75t_SL g4500 ( 
.A(n_4006),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4178),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_SL g4502 ( 
.A(n_4082),
.B(n_3743),
.Y(n_4502)
);

AND2x4_ASAP7_75t_L g4503 ( 
.A(n_4066),
.B(n_3707),
.Y(n_4503)
);

INVx3_ASAP7_75t_L g4504 ( 
.A(n_4043),
.Y(n_4504)
);

INVx3_ASAP7_75t_SL g4505 ( 
.A(n_4165),
.Y(n_4505)
);

BUFx2_ASAP7_75t_SL g4506 ( 
.A(n_4013),
.Y(n_4506)
);

BUFx2_ASAP7_75t_L g4507 ( 
.A(n_3984),
.Y(n_4507)
);

OR2x6_ASAP7_75t_SL g4508 ( 
.A(n_4110),
.B(n_841),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4152),
.B(n_3736),
.Y(n_4509)
);

INVx1_ASAP7_75t_SL g4510 ( 
.A(n_4073),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4084),
.Y(n_4511)
);

AOI21xp5_ASAP7_75t_L g4512 ( 
.A1(n_4127),
.A2(n_2684),
.B(n_2683),
.Y(n_4512)
);

OAI22xp5_ASAP7_75t_L g4513 ( 
.A1(n_3923),
.A2(n_3942),
.B1(n_4048),
.B2(n_4110),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_L g4514 ( 
.A(n_4153),
.B(n_3697),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4084),
.Y(n_4515)
);

AND2x2_ASAP7_75t_L g4516 ( 
.A(n_4152),
.B(n_3736),
.Y(n_4516)
);

INVx3_ASAP7_75t_L g4517 ( 
.A(n_3984),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_4090),
.B(n_1438),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_3968),
.Y(n_4519)
);

AND2x4_ASAP7_75t_L g4520 ( 
.A(n_4089),
.B(n_3697),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_4154),
.B(n_3697),
.Y(n_4521)
);

INVx5_ASAP7_75t_L g4522 ( 
.A(n_4078),
.Y(n_4522)
);

NAND2x1p5_ASAP7_75t_L g4523 ( 
.A(n_4067),
.B(n_3743),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_3879),
.Y(n_4524)
);

AOI22xp33_ASAP7_75t_L g4525 ( 
.A1(n_3992),
.A2(n_1000),
.B1(n_1011),
.B2(n_993),
.Y(n_4525)
);

AND2x4_ASAP7_75t_L g4526 ( 
.A(n_4093),
.B(n_3058),
.Y(n_4526)
);

OAI22xp5_ASAP7_75t_L g4527 ( 
.A1(n_4117),
.A2(n_1013),
.B1(n_1014),
.B2(n_1011),
.Y(n_4527)
);

AOI22xp33_ASAP7_75t_L g4528 ( 
.A1(n_3992),
.A2(n_1020),
.B1(n_1022),
.B2(n_1013),
.Y(n_4528)
);

INVx4_ASAP7_75t_L g4529 ( 
.A(n_3989),
.Y(n_4529)
);

BUFx2_ASAP7_75t_L g4530 ( 
.A(n_4158),
.Y(n_4530)
);

INVxp67_ASAP7_75t_SL g4531 ( 
.A(n_3863),
.Y(n_4531)
);

BUFx3_ASAP7_75t_L g4532 ( 
.A(n_4068),
.Y(n_4532)
);

AOI22xp33_ASAP7_75t_SL g4533 ( 
.A1(n_4117),
.A2(n_1025),
.B1(n_1026),
.B2(n_1020),
.Y(n_4533)
);

INVx4_ASAP7_75t_L g4534 ( 
.A(n_3997),
.Y(n_4534)
);

INVx3_ASAP7_75t_L g4535 ( 
.A(n_4012),
.Y(n_4535)
);

NOR2xp33_ASAP7_75t_L g4536 ( 
.A(n_3918),
.B(n_3063),
.Y(n_4536)
);

INVx3_ASAP7_75t_L g4537 ( 
.A(n_4130),
.Y(n_4537)
);

AND3x1_ASAP7_75t_SL g4538 ( 
.A(n_4040),
.B(n_1026),
.C(n_1025),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_3917),
.B(n_2396),
.Y(n_4539)
);

AOI22xp33_ASAP7_75t_L g4540 ( 
.A1(n_3928),
.A2(n_1030),
.B1(n_1033),
.B2(n_1027),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_3873),
.B(n_3063),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_SL g4542 ( 
.A(n_3960),
.B(n_3063),
.Y(n_4542)
);

AOI22xp5_ASAP7_75t_L g4543 ( 
.A1(n_4071),
.A2(n_845),
.B1(n_846),
.B2(n_842),
.Y(n_4543)
);

AND2x2_ASAP7_75t_L g4544 ( 
.A(n_4096),
.B(n_1440),
.Y(n_4544)
);

BUFx3_ASAP7_75t_L g4545 ( 
.A(n_4172),
.Y(n_4545)
);

INVx3_ASAP7_75t_L g4546 ( 
.A(n_4021),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_4139),
.Y(n_4547)
);

AOI22xp5_ASAP7_75t_L g4548 ( 
.A1(n_4261),
.A2(n_4071),
.B1(n_3958),
.B2(n_4091),
.Y(n_4548)
);

INVx2_ASAP7_75t_L g4549 ( 
.A(n_4203),
.Y(n_4549)
);

INVxp67_ASAP7_75t_L g4550 ( 
.A(n_4281),
.Y(n_4550)
);

OAI22xp5_ASAP7_75t_L g4551 ( 
.A1(n_4508),
.A2(n_3950),
.B1(n_3945),
.B2(n_4102),
.Y(n_4551)
);

A2O1A1Ixp33_ASAP7_75t_L g4552 ( 
.A1(n_4449),
.A2(n_4041),
.B(n_4116),
.C(n_4125),
.Y(n_4552)
);

CKINVDCx5p33_ASAP7_75t_R g4553 ( 
.A(n_4253),
.Y(n_4553)
);

INVx4_ASAP7_75t_L g4554 ( 
.A(n_4486),
.Y(n_4554)
);

O2A1O1Ixp33_ASAP7_75t_SL g4555 ( 
.A1(n_4395),
.A2(n_4292),
.B(n_4265),
.C(n_4264),
.Y(n_4555)
);

AOI22xp5_ASAP7_75t_L g4556 ( 
.A1(n_4263),
.A2(n_3958),
.B1(n_857),
.B2(n_858),
.Y(n_4556)
);

A2O1A1Ixp33_ASAP7_75t_L g4557 ( 
.A1(n_4449),
.A2(n_3867),
.B(n_4083),
.C(n_3961),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4210),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4221),
.Y(n_4559)
);

O2A1O1Ixp33_ASAP7_75t_SL g4560 ( 
.A1(n_4265),
.A2(n_1030),
.B(n_1033),
.C(n_1027),
.Y(n_4560)
);

INVx3_ASAP7_75t_L g4561 ( 
.A(n_4277),
.Y(n_4561)
);

A2O1A1Ixp33_ASAP7_75t_L g4562 ( 
.A1(n_4250),
.A2(n_3951),
.B(n_3949),
.C(n_4054),
.Y(n_4562)
);

A2O1A1Ixp33_ASAP7_75t_L g4563 ( 
.A1(n_4250),
.A2(n_4011),
.B(n_4010),
.C(n_3988),
.Y(n_4563)
);

INVx2_ASAP7_75t_L g4564 ( 
.A(n_4226),
.Y(n_4564)
);

AND2x4_ASAP7_75t_L g4565 ( 
.A(n_4243),
.B(n_4016),
.Y(n_4565)
);

OAI21xp5_ASAP7_75t_L g4566 ( 
.A1(n_4218),
.A2(n_3934),
.B(n_4087),
.Y(n_4566)
);

AOI22xp5_ASAP7_75t_L g4567 ( 
.A1(n_4263),
.A2(n_4411),
.B1(n_4342),
.B2(n_4513),
.Y(n_4567)
);

AND2x4_ASAP7_75t_L g4568 ( 
.A(n_4243),
.B(n_4025),
.Y(n_4568)
);

A2O1A1Ixp33_ASAP7_75t_L g4569 ( 
.A1(n_4411),
.A2(n_1045),
.B(n_1049),
.C(n_1038),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4240),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_SL g4571 ( 
.A(n_4200),
.B(n_4149),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4255),
.Y(n_4572)
);

AO31x2_ASAP7_75t_L g4573 ( 
.A1(n_4405),
.A2(n_4185),
.A3(n_4196),
.B(n_4029),
.Y(n_4573)
);

AOI21xp33_ASAP7_75t_L g4574 ( 
.A1(n_4217),
.A2(n_4029),
.B(n_4021),
.Y(n_4574)
);

AOI22xp33_ASAP7_75t_L g4575 ( 
.A1(n_4484),
.A2(n_1059),
.B1(n_1060),
.B2(n_1054),
.Y(n_4575)
);

NAND2xp5_ASAP7_75t_L g4576 ( 
.A(n_4388),
.B(n_4394),
.Y(n_4576)
);

A2O1A1Ixp33_ASAP7_75t_L g4577 ( 
.A1(n_4206),
.A2(n_1059),
.B(n_1060),
.C(n_1054),
.Y(n_4577)
);

BUFx3_ASAP7_75t_L g4578 ( 
.A(n_4216),
.Y(n_4578)
);

AO31x2_ASAP7_75t_L g4579 ( 
.A1(n_4476),
.A2(n_4248),
.A3(n_4381),
.B(n_4314),
.Y(n_4579)
);

OAI21xp5_ASAP7_75t_L g4580 ( 
.A1(n_4229),
.A2(n_4002),
.B(n_4061),
.Y(n_4580)
);

AOI21x1_ASAP7_75t_SL g4581 ( 
.A1(n_4509),
.A2(n_4516),
.B(n_4518),
.Y(n_4581)
);

A2O1A1Ixp33_ASAP7_75t_L g4582 ( 
.A1(n_4513),
.A2(n_1064),
.B(n_1065),
.C(n_1061),
.Y(n_4582)
);

OA21x2_ASAP7_75t_L g4583 ( 
.A1(n_4262),
.A2(n_4037),
.B(n_4140),
.Y(n_4583)
);

AO32x2_ASAP7_75t_L g4584 ( 
.A1(n_4423),
.A2(n_4185),
.A3(n_3920),
.B1(n_6),
.B2(n_4),
.Y(n_4584)
);

OA21x2_ASAP7_75t_L g4585 ( 
.A1(n_4262),
.A2(n_4177),
.B(n_4145),
.Y(n_4585)
);

AOI22xp33_ASAP7_75t_L g4586 ( 
.A1(n_4484),
.A2(n_1089),
.B1(n_1090),
.B2(n_1082),
.Y(n_4586)
);

AOI221xp5_ASAP7_75t_L g4587 ( 
.A1(n_4319),
.A2(n_860),
.B1(n_864),
.B2(n_859),
.C(n_856),
.Y(n_4587)
);

INVx2_ASAP7_75t_SL g4588 ( 
.A(n_4220),
.Y(n_4588)
);

AO21x2_ASAP7_75t_L g4589 ( 
.A1(n_4512),
.A2(n_4064),
.B(n_4188),
.Y(n_4589)
);

O2A1O1Ixp33_ASAP7_75t_L g4590 ( 
.A1(n_4273),
.A2(n_1089),
.B(n_1090),
.C(n_1082),
.Y(n_4590)
);

AO31x2_ASAP7_75t_L g4591 ( 
.A1(n_4476),
.A2(n_4190),
.A3(n_3920),
.B(n_4135),
.Y(n_4591)
);

AO31x2_ASAP7_75t_L g4592 ( 
.A1(n_4248),
.A2(n_4314),
.A3(n_4381),
.B(n_4492),
.Y(n_4592)
);

AO31x2_ASAP7_75t_L g4593 ( 
.A1(n_4488),
.A2(n_3920),
.A3(n_2684),
.B(n_2683),
.Y(n_4593)
);

AO31x2_ASAP7_75t_L g4594 ( 
.A1(n_4512),
.A2(n_2684),
.A3(n_1093),
.B(n_1094),
.Y(n_4594)
);

AOI21xp5_ASAP7_75t_L g4595 ( 
.A1(n_4531),
.A2(n_3104),
.B(n_3045),
.Y(n_4595)
);

O2A1O1Ixp33_ASAP7_75t_L g4596 ( 
.A1(n_4319),
.A2(n_1093),
.B(n_1094),
.C(n_1091),
.Y(n_4596)
);

INVx2_ASAP7_75t_L g4597 ( 
.A(n_4259),
.Y(n_4597)
);

AOI21xp5_ASAP7_75t_L g4598 ( 
.A1(n_4242),
.A2(n_3104),
.B(n_3045),
.Y(n_4598)
);

INVxp67_ASAP7_75t_SL g4599 ( 
.A(n_4272),
.Y(n_4599)
);

A2O1A1Ixp33_ASAP7_75t_L g4600 ( 
.A1(n_4432),
.A2(n_1102),
.B(n_1105),
.C(n_1091),
.Y(n_4600)
);

OAI22xp33_ASAP7_75t_L g4601 ( 
.A1(n_4423),
.A2(n_1105),
.B1(n_1108),
.B2(n_1102),
.Y(n_4601)
);

INVx6_ASAP7_75t_L g4602 ( 
.A(n_4202),
.Y(n_4602)
);

OAI21xp5_ASAP7_75t_L g4603 ( 
.A1(n_4318),
.A2(n_1110),
.B(n_1108),
.Y(n_4603)
);

INVx2_ASAP7_75t_L g4604 ( 
.A(n_4268),
.Y(n_4604)
);

A2O1A1Ixp33_ASAP7_75t_L g4605 ( 
.A1(n_4432),
.A2(n_1116),
.B(n_1117),
.C(n_1110),
.Y(n_4605)
);

AO31x2_ASAP7_75t_L g4606 ( 
.A1(n_4497),
.A2(n_1117),
.A3(n_1120),
.B(n_1116),
.Y(n_4606)
);

AOI22xp33_ASAP7_75t_SL g4607 ( 
.A1(n_4378),
.A2(n_867),
.B1(n_868),
.B2(n_865),
.Y(n_4607)
);

AOI211xp5_ASAP7_75t_L g4608 ( 
.A1(n_4428),
.A2(n_892),
.B(n_903),
.C(n_878),
.Y(n_4608)
);

NAND3xp33_ASAP7_75t_L g4609 ( 
.A(n_4543),
.B(n_1442),
.C(n_1441),
.Y(n_4609)
);

O2A1O1Ixp33_ASAP7_75t_SL g4610 ( 
.A1(n_4527),
.A2(n_1448),
.B(n_1450),
.C(n_1445),
.Y(n_4610)
);

AOI21xp5_ASAP7_75t_L g4611 ( 
.A1(n_4242),
.A2(n_2923),
.B(n_2920),
.Y(n_4611)
);

HB1xp67_ASAP7_75t_L g4612 ( 
.A(n_4354),
.Y(n_4612)
);

OAI21xp5_ASAP7_75t_L g4613 ( 
.A1(n_4285),
.A2(n_1453),
.B(n_1452),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4274),
.Y(n_4614)
);

OR2x6_ASAP7_75t_L g4615 ( 
.A(n_4341),
.B(n_3067),
.Y(n_4615)
);

AOI21xp5_ASAP7_75t_L g4616 ( 
.A1(n_4209),
.A2(n_2932),
.B(n_2923),
.Y(n_4616)
);

NOR2xp33_ASAP7_75t_L g4617 ( 
.A(n_4494),
.B(n_869),
.Y(n_4617)
);

NAND2xp5_ASAP7_75t_L g4618 ( 
.A(n_4387),
.B(n_871),
.Y(n_4618)
);

INVx2_ASAP7_75t_L g4619 ( 
.A(n_4282),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_L g4620 ( 
.A(n_4254),
.B(n_873),
.Y(n_4620)
);

BUFx2_ASAP7_75t_L g4621 ( 
.A(n_4326),
.Y(n_4621)
);

OAI22xp5_ASAP7_75t_SL g4622 ( 
.A1(n_4473),
.A2(n_876),
.B1(n_882),
.B2(n_874),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4284),
.Y(n_4623)
);

AO31x2_ASAP7_75t_L g4624 ( 
.A1(n_4474),
.A2(n_2318),
.A3(n_2320),
.B(n_2312),
.Y(n_4624)
);

AOI21xp5_ASAP7_75t_L g4625 ( 
.A1(n_4209),
.A2(n_2932),
.B(n_2923),
.Y(n_4625)
);

INVx1_ASAP7_75t_SL g4626 ( 
.A(n_4349),
.Y(n_4626)
);

AO31x2_ASAP7_75t_L g4627 ( 
.A1(n_4524),
.A2(n_2318),
.A3(n_2320),
.B(n_2312),
.Y(n_4627)
);

AOI21xp5_ASAP7_75t_L g4628 ( 
.A1(n_4201),
.A2(n_2972),
.B(n_2932),
.Y(n_4628)
);

OAI21xp5_ASAP7_75t_L g4629 ( 
.A1(n_4525),
.A2(n_1460),
.B(n_1454),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4293),
.Y(n_4630)
);

CKINVDCx5p33_ASAP7_75t_R g4631 ( 
.A(n_4227),
.Y(n_4631)
);

AND2x4_ASAP7_75t_L g4632 ( 
.A(n_4243),
.B(n_3067),
.Y(n_4632)
);

INVxp33_ASAP7_75t_SL g4633 ( 
.A(n_4266),
.Y(n_4633)
);

AOI21xp5_ASAP7_75t_L g4634 ( 
.A1(n_4201),
.A2(n_2972),
.B(n_2932),
.Y(n_4634)
);

AO31x2_ASAP7_75t_L g4635 ( 
.A1(n_4401),
.A2(n_2329),
.A3(n_2330),
.B(n_2321),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4297),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4254),
.B(n_883),
.Y(n_4637)
);

AND2x2_ASAP7_75t_L g4638 ( 
.A(n_4442),
.B(n_1461),
.Y(n_4638)
);

BUFx12f_ASAP7_75t_L g4639 ( 
.A(n_4202),
.Y(n_4639)
);

O2A1O1Ixp33_ASAP7_75t_SL g4640 ( 
.A1(n_4527),
.A2(n_1464),
.B(n_1465),
.C(n_1462),
.Y(n_4640)
);

NOR2xp33_ASAP7_75t_L g4641 ( 
.A(n_4483),
.B(n_889),
.Y(n_4641)
);

OAI221xp5_ASAP7_75t_L g4642 ( 
.A1(n_4245),
.A2(n_895),
.B1(n_896),
.B2(n_894),
.C(n_891),
.Y(n_4642)
);

CKINVDCx20_ASAP7_75t_R g4643 ( 
.A(n_4280),
.Y(n_4643)
);

AO31x2_ASAP7_75t_L g4644 ( 
.A1(n_4332),
.A2(n_2329),
.A3(n_2330),
.B(n_2321),
.Y(n_4644)
);

CKINVDCx5p33_ASAP7_75t_R g4645 ( 
.A(n_4309),
.Y(n_4645)
);

OAI21x1_ASAP7_75t_L g4646 ( 
.A1(n_4438),
.A2(n_4469),
.B(n_4478),
.Y(n_4646)
);

CKINVDCx20_ASAP7_75t_R g4647 ( 
.A(n_4244),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4272),
.Y(n_4648)
);

O2A1O1Ixp33_ASAP7_75t_SL g4649 ( 
.A1(n_4217),
.A2(n_1469),
.B(n_1471),
.C(n_1467),
.Y(n_4649)
);

O2A1O1Ixp33_ASAP7_75t_L g4650 ( 
.A1(n_4235),
.A2(n_1479),
.B(n_1483),
.C(n_1477),
.Y(n_4650)
);

O2A1O1Ixp33_ASAP7_75t_SL g4651 ( 
.A1(n_4502),
.A2(n_4317),
.B(n_4498),
.C(n_4514),
.Y(n_4651)
);

NOR2xp33_ASAP7_75t_SL g4652 ( 
.A(n_4490),
.B(n_4371),
.Y(n_4652)
);

AOI221x1_ASAP7_75t_L g4653 ( 
.A1(n_4390),
.A2(n_1488),
.B1(n_1491),
.B2(n_1487),
.C(n_1485),
.Y(n_4653)
);

INVxp67_ASAP7_75t_SL g4654 ( 
.A(n_4257),
.Y(n_4654)
);

AOI21xp5_ASAP7_75t_L g4655 ( 
.A1(n_4500),
.A2(n_2975),
.B(n_2972),
.Y(n_4655)
);

BUFx10_ASAP7_75t_L g4656 ( 
.A(n_4202),
.Y(n_4656)
);

OAI21xp5_ASAP7_75t_L g4657 ( 
.A1(n_4528),
.A2(n_1501),
.B(n_1498),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4322),
.Y(n_4658)
);

OAI22xp5_ASAP7_75t_SL g4659 ( 
.A1(n_4437),
.A2(n_905),
.B1(n_906),
.B2(n_904),
.Y(n_4659)
);

OR2x2_ASAP7_75t_L g4660 ( 
.A(n_4208),
.B(n_1363),
.Y(n_4660)
);

AO31x2_ASAP7_75t_L g4661 ( 
.A1(n_4332),
.A2(n_2334),
.A3(n_2335),
.B(n_2331),
.Y(n_4661)
);

O2A1O1Ixp33_ASAP7_75t_L g4662 ( 
.A1(n_4402),
.A2(n_1369),
.B(n_1372),
.C(n_1368),
.Y(n_4662)
);

A2O1A1Ixp33_ASAP7_75t_L g4663 ( 
.A1(n_4378),
.A2(n_908),
.B(n_913),
.C(n_907),
.Y(n_4663)
);

O2A1O1Ixp33_ASAP7_75t_L g4664 ( 
.A1(n_4519),
.A2(n_1378),
.B(n_1380),
.C(n_1376),
.Y(n_4664)
);

AOI21x1_ASAP7_75t_L g4665 ( 
.A1(n_4407),
.A2(n_4267),
.B(n_4541),
.Y(n_4665)
);

NAND2x1p5_ASAP7_75t_L g4666 ( 
.A(n_4278),
.B(n_3067),
.Y(n_4666)
);

OAI22xp5_ASAP7_75t_L g4667 ( 
.A1(n_4533),
.A2(n_915),
.B1(n_916),
.B2(n_914),
.Y(n_4667)
);

AOI221x1_ASAP7_75t_L g4668 ( 
.A1(n_4390),
.A2(n_1533),
.B1(n_1537),
.B2(n_1532),
.C(n_1531),
.Y(n_4668)
);

OAI22x1_ASAP7_75t_L g4669 ( 
.A1(n_4199),
.A2(n_952),
.B1(n_973),
.B2(n_931),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_4335),
.B(n_918),
.Y(n_4670)
);

AOI22xp5_ASAP7_75t_L g4671 ( 
.A1(n_4534),
.A2(n_4538),
.B1(n_4462),
.B2(n_4418),
.Y(n_4671)
);

AND2x2_ASAP7_75t_SL g4672 ( 
.A(n_4339),
.B(n_2972),
.Y(n_4672)
);

AND2x2_ASAP7_75t_L g4673 ( 
.A(n_4447),
.B(n_1381),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_4349),
.B(n_926),
.Y(n_4674)
);

AOI21xp5_ASAP7_75t_L g4675 ( 
.A1(n_4500),
.A2(n_3001),
.B(n_2975),
.Y(n_4675)
);

OAI21x1_ASAP7_75t_SL g4676 ( 
.A1(n_4366),
.A2(n_1391),
.B(n_1389),
.Y(n_4676)
);

INVx4_ASAP7_75t_SL g4677 ( 
.A(n_4443),
.Y(n_4677)
);

BUFx6f_ASAP7_75t_L g4678 ( 
.A(n_4420),
.Y(n_4678)
);

AO32x2_ASAP7_75t_L g4679 ( 
.A1(n_4256),
.A2(n_8),
.A3(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_4679)
);

AOI22xp5_ASAP7_75t_L g4680 ( 
.A1(n_4534),
.A2(n_949),
.B1(n_950),
.B2(n_947),
.Y(n_4680)
);

OAI21x1_ASAP7_75t_L g4681 ( 
.A1(n_4469),
.A2(n_2416),
.B(n_2400),
.Y(n_4681)
);

OAI21x1_ASAP7_75t_L g4682 ( 
.A1(n_4489),
.A2(n_2400),
.B(n_2367),
.Y(n_4682)
);

AOI22xp33_ASAP7_75t_L g4683 ( 
.A1(n_4545),
.A2(n_1395),
.B1(n_1393),
.B2(n_957),
.Y(n_4683)
);

CKINVDCx20_ASAP7_75t_R g4684 ( 
.A(n_4495),
.Y(n_4684)
);

NOR2xp33_ASAP7_75t_L g4685 ( 
.A(n_4360),
.B(n_951),
.Y(n_4685)
);

AOI21xp5_ASAP7_75t_L g4686 ( 
.A1(n_4257),
.A2(n_3001),
.B(n_2975),
.Y(n_4686)
);

AOI22xp33_ASAP7_75t_L g4687 ( 
.A1(n_4530),
.A2(n_961),
.B1(n_965),
.B2(n_960),
.Y(n_4687)
);

O2A1O1Ixp33_ASAP7_75t_SL g4688 ( 
.A1(n_4514),
.A2(n_1532),
.B(n_1533),
.C(n_1531),
.Y(n_4688)
);

OAI221xp5_ASAP7_75t_L g4689 ( 
.A1(n_4410),
.A2(n_971),
.B1(n_974),
.B2(n_970),
.C(n_966),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4334),
.Y(n_4690)
);

AO32x2_ASAP7_75t_L g4691 ( 
.A1(n_4256),
.A2(n_8),
.A3(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_L g4692 ( 
.A(n_4419),
.B(n_975),
.Y(n_4692)
);

O2A1O1Ixp33_ASAP7_75t_L g4693 ( 
.A1(n_4422),
.A2(n_1539),
.B(n_1541),
.C(n_1537),
.Y(n_4693)
);

NAND3xp33_ASAP7_75t_L g4694 ( 
.A(n_4376),
.B(n_4377),
.C(n_4491),
.Y(n_4694)
);

OR2x2_ASAP7_75t_L g4695 ( 
.A(n_4298),
.B(n_1539),
.Y(n_4695)
);

O2A1O1Ixp33_ASAP7_75t_SL g4696 ( 
.A1(n_4521),
.A2(n_1544),
.B(n_1545),
.C(n_1541),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4336),
.Y(n_4697)
);

AO31x2_ASAP7_75t_L g4698 ( 
.A1(n_4482),
.A2(n_2334),
.A3(n_2335),
.B(n_2331),
.Y(n_4698)
);

NOR2x1_ASAP7_75t_L g4699 ( 
.A(n_4506),
.B(n_1544),
.Y(n_4699)
);

AOI22xp33_ASAP7_75t_SL g4700 ( 
.A1(n_4546),
.A2(n_983),
.B1(n_986),
.B2(n_982),
.Y(n_4700)
);

O2A1O1Ixp33_ASAP7_75t_L g4701 ( 
.A1(n_4377),
.A2(n_1546),
.B(n_1547),
.C(n_1545),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4338),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4356),
.Y(n_4703)
);

OAI21x1_ASAP7_75t_L g4704 ( 
.A1(n_4537),
.A2(n_2400),
.B(n_2367),
.Y(n_4704)
);

AOI21xp5_ASAP7_75t_L g4705 ( 
.A1(n_4313),
.A2(n_3001),
.B(n_2975),
.Y(n_4705)
);

O2A1O1Ixp33_ASAP7_75t_SL g4706 ( 
.A1(n_4521),
.A2(n_1547),
.B(n_1548),
.C(n_1546),
.Y(n_4706)
);

OAI22xp5_ASAP7_75t_L g4707 ( 
.A1(n_4425),
.A2(n_999),
.B1(n_1001),
.B2(n_996),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_4459),
.B(n_1002),
.Y(n_4708)
);

OAI21x1_ASAP7_75t_L g4709 ( 
.A1(n_4537),
.A2(n_2413),
.B(n_2367),
.Y(n_4709)
);

AOI21xp5_ASAP7_75t_L g4710 ( 
.A1(n_4313),
.A2(n_3002),
.B(n_3001),
.Y(n_4710)
);

A2O1A1Ixp33_ASAP7_75t_L g4711 ( 
.A1(n_4425),
.A2(n_1005),
.B(n_1007),
.C(n_1003),
.Y(n_4711)
);

INVx4_ASAP7_75t_SL g4712 ( 
.A(n_4207),
.Y(n_4712)
);

AOI21xp5_ASAP7_75t_L g4713 ( 
.A1(n_4457),
.A2(n_3015),
.B(n_3002),
.Y(n_4713)
);

A2O1A1Ixp33_ASAP7_75t_L g4714 ( 
.A1(n_4536),
.A2(n_1009),
.B(n_1012),
.C(n_1008),
.Y(n_4714)
);

INVx4_ASAP7_75t_L g4715 ( 
.A(n_4486),
.Y(n_4715)
);

OAI21xp5_ASAP7_75t_L g4716 ( 
.A1(n_4331),
.A2(n_4540),
.B(n_4544),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4302),
.Y(n_4717)
);

HB1xp67_ASAP7_75t_L g4718 ( 
.A(n_4246),
.Y(n_4718)
);

AO31x2_ASAP7_75t_L g4719 ( 
.A1(n_4536),
.A2(n_2342),
.A3(n_2340),
.B(n_1549),
.Y(n_4719)
);

NAND2xp5_ASAP7_75t_L g4720 ( 
.A(n_4463),
.B(n_1018),
.Y(n_4720)
);

INVx2_ASAP7_75t_L g4721 ( 
.A(n_4363),
.Y(n_4721)
);

AOI22xp5_ASAP7_75t_L g4722 ( 
.A1(n_4538),
.A2(n_1023),
.B1(n_1024),
.B2(n_1019),
.Y(n_4722)
);

O2A1O1Ixp33_ASAP7_75t_SL g4723 ( 
.A1(n_4205),
.A2(n_1549),
.B(n_1550),
.C(n_1548),
.Y(n_4723)
);

OAI21xp5_ASAP7_75t_L g4724 ( 
.A1(n_4540),
.A2(n_1036),
.B(n_1034),
.Y(n_4724)
);

AOI21xp5_ASAP7_75t_L g4725 ( 
.A1(n_4457),
.A2(n_3015),
.B(n_3002),
.Y(n_4725)
);

INVx1_ASAP7_75t_L g4726 ( 
.A(n_4312),
.Y(n_4726)
);

INVx4_ASAP7_75t_L g4727 ( 
.A(n_4486),
.Y(n_4727)
);

O2A1O1Ixp33_ASAP7_75t_SL g4728 ( 
.A1(n_4236),
.A2(n_1551),
.B(n_1553),
.C(n_1550),
.Y(n_4728)
);

CKINVDCx5p33_ASAP7_75t_R g4729 ( 
.A(n_4344),
.Y(n_4729)
);

NOR2xp33_ASAP7_75t_SL g4730 ( 
.A(n_4230),
.B(n_3067),
.Y(n_4730)
);

O2A1O1Ixp33_ASAP7_75t_SL g4731 ( 
.A1(n_4247),
.A2(n_1553),
.B(n_1554),
.C(n_1551),
.Y(n_4731)
);

AOI21xp5_ASAP7_75t_L g4732 ( 
.A1(n_4542),
.A2(n_3015),
.B(n_3002),
.Y(n_4732)
);

A2O1A1Ixp33_ASAP7_75t_L g4733 ( 
.A1(n_4283),
.A2(n_1040),
.B(n_1041),
.C(n_1037),
.Y(n_4733)
);

OAI21x1_ASAP7_75t_L g4734 ( 
.A1(n_4535),
.A2(n_2414),
.B(n_2413),
.Y(n_4734)
);

INVx1_ASAP7_75t_L g4735 ( 
.A(n_4287),
.Y(n_4735)
);

CKINVDCx11_ASAP7_75t_R g4736 ( 
.A(n_4204),
.Y(n_4736)
);

INVx4_ASAP7_75t_L g4737 ( 
.A(n_4380),
.Y(n_4737)
);

A2O1A1Ixp33_ASAP7_75t_L g4738 ( 
.A1(n_4283),
.A2(n_1046),
.B(n_1047),
.C(n_1042),
.Y(n_4738)
);

AOI21xp5_ASAP7_75t_L g4739 ( 
.A1(n_4251),
.A2(n_3015),
.B(n_3094),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4466),
.B(n_1048),
.Y(n_4740)
);

AO31x2_ASAP7_75t_L g4741 ( 
.A1(n_4539),
.A2(n_4541),
.A3(n_4493),
.B(n_4487),
.Y(n_4741)
);

OAI21x1_ASAP7_75t_L g4742 ( 
.A1(n_4535),
.A2(n_2414),
.B(n_2413),
.Y(n_4742)
);

O2A1O1Ixp33_ASAP7_75t_L g4743 ( 
.A1(n_4211),
.A2(n_1558),
.B(n_1559),
.C(n_1554),
.Y(n_4743)
);

O2A1O1Ixp33_ASAP7_75t_SL g4744 ( 
.A1(n_4246),
.A2(n_1559),
.B(n_1561),
.C(n_1558),
.Y(n_4744)
);

O2A1O1Ixp33_ASAP7_75t_L g4745 ( 
.A1(n_4211),
.A2(n_1561),
.B(n_1860),
.C(n_1857),
.Y(n_4745)
);

O2A1O1Ixp33_ASAP7_75t_L g4746 ( 
.A1(n_4385),
.A2(n_1860),
.B(n_1867),
.C(n_1857),
.Y(n_4746)
);

AOI21xp5_ASAP7_75t_L g4747 ( 
.A1(n_4251),
.A2(n_3164),
.B(n_3094),
.Y(n_4747)
);

AOI21xp5_ASAP7_75t_L g4748 ( 
.A1(n_4539),
.A2(n_3164),
.B(n_3094),
.Y(n_4748)
);

OAI22xp33_ASAP7_75t_L g4749 ( 
.A1(n_4271),
.A2(n_1101),
.B1(n_1127),
.B2(n_1081),
.Y(n_4749)
);

OAI21xp5_ASAP7_75t_L g4750 ( 
.A1(n_4323),
.A2(n_1070),
.B(n_1066),
.Y(n_4750)
);

AOI22xp33_ASAP7_75t_L g4751 ( 
.A1(n_4271),
.A2(n_1072),
.B1(n_1073),
.B2(n_1071),
.Y(n_4751)
);

AOI21xp5_ASAP7_75t_L g4752 ( 
.A1(n_4323),
.A2(n_3164),
.B(n_3094),
.Y(n_4752)
);

BUFx12f_ASAP7_75t_L g4753 ( 
.A(n_4477),
.Y(n_4753)
);

AOI221xp5_ASAP7_75t_L g4754 ( 
.A1(n_4386),
.A2(n_1086),
.B1(n_1088),
.B2(n_1078),
.C(n_1075),
.Y(n_4754)
);

O2A1O1Ixp33_ASAP7_75t_L g4755 ( 
.A1(n_4300),
.A2(n_1867),
.B(n_2294),
.C(n_2291),
.Y(n_4755)
);

OAI22xp33_ASAP7_75t_L g4756 ( 
.A1(n_4271),
.A2(n_1113),
.B1(n_1092),
.B2(n_1095),
.Y(n_4756)
);

CKINVDCx5p33_ASAP7_75t_R g4757 ( 
.A(n_4475),
.Y(n_4757)
);

AO31x2_ASAP7_75t_L g4758 ( 
.A1(n_4511),
.A2(n_2342),
.A3(n_2340),
.B(n_1909),
.Y(n_4758)
);

AOI21xp33_ASAP7_75t_L g4759 ( 
.A1(n_4510),
.A2(n_3164),
.B(n_1098),
.Y(n_4759)
);

BUFx3_ASAP7_75t_L g4760 ( 
.A(n_4270),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4470),
.B(n_1104),
.Y(n_4761)
);

OAI21x1_ASAP7_75t_L g4762 ( 
.A1(n_4391),
.A2(n_2414),
.B(n_2449),
.Y(n_4762)
);

NOR2xp33_ASAP7_75t_L g4763 ( 
.A(n_4472),
.B(n_1107),
.Y(n_4763)
);

INVx1_ASAP7_75t_SL g4764 ( 
.A(n_4300),
.Y(n_4764)
);

AOI21xp5_ASAP7_75t_L g4765 ( 
.A1(n_4436),
.A2(n_2414),
.B(n_2572),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_L g4766 ( 
.A(n_4471),
.B(n_1114),
.Y(n_4766)
);

AOI21xp5_ASAP7_75t_L g4767 ( 
.A1(n_4436),
.A2(n_4391),
.B(n_4289),
.Y(n_4767)
);

A2O1A1Ixp33_ASAP7_75t_L g4768 ( 
.A1(n_4382),
.A2(n_1125),
.B(n_1126),
.C(n_1118),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4289),
.Y(n_4769)
);

NAND2xp5_ASAP7_75t_L g4770 ( 
.A(n_4424),
.B(n_1135),
.Y(n_4770)
);

OAI22xp5_ASAP7_75t_L g4771 ( 
.A1(n_4510),
.A2(n_1136),
.B1(n_2642),
.B2(n_2639),
.Y(n_4771)
);

INVx2_ASAP7_75t_L g4772 ( 
.A(n_4364),
.Y(n_4772)
);

BUFx6f_ASAP7_75t_L g4773 ( 
.A(n_4207),
.Y(n_4773)
);

AND2x4_ASAP7_75t_L g4774 ( 
.A(n_4243),
.B(n_2756),
.Y(n_4774)
);

OAI21xp5_ASAP7_75t_L g4775 ( 
.A1(n_4523),
.A2(n_1915),
.B(n_1908),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4198),
.Y(n_4776)
);

AO31x2_ASAP7_75t_L g4777 ( 
.A1(n_4515),
.A2(n_1924),
.A3(n_1936),
.B(n_1908),
.Y(n_4777)
);

A2O1A1Ixp33_ASAP7_75t_L g4778 ( 
.A1(n_4382),
.A2(n_1203),
.B(n_1220),
.C(n_1219),
.Y(n_4778)
);

AOI22xp5_ASAP7_75t_SL g4779 ( 
.A1(n_4339),
.A2(n_10),
.B1(n_5),
.B2(n_9),
.Y(n_4779)
);

NAND2x1p5_ASAP7_75t_L g4780 ( 
.A(n_4529),
.B(n_2639),
.Y(n_4780)
);

OAI22xp5_ASAP7_75t_L g4781 ( 
.A1(n_4435),
.A2(n_2642),
.B1(n_2665),
.B2(n_2338),
.Y(n_4781)
);

AO32x2_ASAP7_75t_L g4782 ( 
.A1(n_4464),
.A2(n_13),
.A3(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_4782)
);

AOI21xp5_ASAP7_75t_L g4783 ( 
.A1(n_4393),
.A2(n_2735),
.B(n_2572),
.Y(n_4783)
);

OR2x6_ASAP7_75t_L g4784 ( 
.A(n_4353),
.B(n_4252),
.Y(n_4784)
);

OAI21x1_ASAP7_75t_L g4785 ( 
.A1(n_4393),
.A2(n_1936),
.B(n_1924),
.Y(n_4785)
);

AOI22xp33_ASAP7_75t_L g4786 ( 
.A1(n_4445),
.A2(n_2995),
.B1(n_3033),
.B2(n_2992),
.Y(n_4786)
);

OAI21xp5_ASAP7_75t_L g4787 ( 
.A1(n_4523),
.A2(n_1939),
.B(n_1937),
.Y(n_4787)
);

NAND2xp5_ASAP7_75t_L g4788 ( 
.A(n_4397),
.B(n_58),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4198),
.Y(n_4789)
);

AOI21xp5_ASAP7_75t_L g4790 ( 
.A1(n_4379),
.A2(n_2735),
.B(n_2081),
.Y(n_4790)
);

OR2x2_ASAP7_75t_L g4791 ( 
.A(n_4325),
.B(n_1219),
.Y(n_4791)
);

AOI221xp5_ASAP7_75t_SL g4792 ( 
.A1(n_4431),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.C(n_15),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4198),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4408),
.B(n_59),
.Y(n_4794)
);

OAI221xp5_ASAP7_75t_L g4795 ( 
.A1(n_4435),
.A2(n_1225),
.B1(n_1224),
.B2(n_1222),
.C(n_2475),
.Y(n_4795)
);

OAI21xp5_ASAP7_75t_L g4796 ( 
.A1(n_4288),
.A2(n_1944),
.B(n_1941),
.Y(n_4796)
);

INVx3_ASAP7_75t_L g4797 ( 
.A(n_4277),
.Y(n_4797)
);

AO21x1_ASAP7_75t_L g4798 ( 
.A1(n_4448),
.A2(n_15),
.B(n_16),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4198),
.Y(n_4799)
);

OAI21x1_ASAP7_75t_L g4800 ( 
.A1(n_4311),
.A2(n_1944),
.B(n_1941),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_L g4801 ( 
.A(n_4416),
.B(n_59),
.Y(n_4801)
);

INVx1_ASAP7_75t_L g4802 ( 
.A(n_4198),
.Y(n_4802)
);

AOI21xp5_ASAP7_75t_L g4803 ( 
.A1(n_4379),
.A2(n_2735),
.B(n_2665),
.Y(n_4803)
);

CKINVDCx11_ASAP7_75t_R g4804 ( 
.A(n_4475),
.Y(n_4804)
);

OAI22xp33_ASAP7_75t_L g4805 ( 
.A1(n_4353),
.A2(n_2665),
.B1(n_2642),
.B2(n_2338),
.Y(n_4805)
);

A2O1A1Ixp33_ASAP7_75t_L g4806 ( 
.A1(n_4214),
.A2(n_1222),
.B(n_61),
.C(n_63),
.Y(n_4806)
);

NOR2xp33_ASAP7_75t_L g4807 ( 
.A(n_4453),
.B(n_60),
.Y(n_4807)
);

INVx3_ASAP7_75t_L g4808 ( 
.A(n_4224),
.Y(n_4808)
);

O2A1O1Ixp33_ASAP7_75t_L g4809 ( 
.A1(n_4223),
.A2(n_4233),
.B(n_4238),
.C(n_4234),
.Y(n_4809)
);

AOI21xp5_ASAP7_75t_L g4810 ( 
.A1(n_4232),
.A2(n_2735),
.B(n_2665),
.Y(n_4810)
);

INVx3_ASAP7_75t_L g4811 ( 
.A(n_4224),
.Y(n_4811)
);

OAI21x1_ASAP7_75t_L g4812 ( 
.A1(n_4311),
.A2(n_1954),
.B(n_1946),
.Y(n_4812)
);

OR2x2_ASAP7_75t_L g4813 ( 
.A(n_4325),
.B(n_1853),
.Y(n_4813)
);

NAND2xp5_ASAP7_75t_L g4814 ( 
.A(n_4450),
.B(n_60),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4501),
.Y(n_4815)
);

AO31x2_ASAP7_75t_L g4816 ( 
.A1(n_4547),
.A2(n_1960),
.A3(n_1963),
.B(n_1956),
.Y(n_4816)
);

AOI21xp33_ASAP7_75t_L g4817 ( 
.A1(n_4345),
.A2(n_1963),
.B(n_1960),
.Y(n_4817)
);

OAI21xp33_ASAP7_75t_L g4818 ( 
.A1(n_4403),
.A2(n_1864),
.B(n_1853),
.Y(n_4818)
);

AND2x2_ASAP7_75t_L g4819 ( 
.A(n_4426),
.B(n_64),
.Y(n_4819)
);

AOI22xp5_ASAP7_75t_L g4820 ( 
.A1(n_4353),
.A2(n_2995),
.B1(n_3033),
.B2(n_2992),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4446),
.Y(n_4821)
);

HB1xp67_ASAP7_75t_L g4822 ( 
.A(n_4329),
.Y(n_4822)
);

OAI22xp33_ASAP7_75t_L g4823 ( 
.A1(n_4252),
.A2(n_2642),
.B1(n_2338),
.B2(n_19),
.Y(n_4823)
);

NOR2xp67_ASAP7_75t_SL g4824 ( 
.A(n_4316),
.B(n_2642),
.Y(n_4824)
);

AND2x4_ASAP7_75t_L g4825 ( 
.A(n_4316),
.B(n_2756),
.Y(n_4825)
);

NAND2x1p5_ASAP7_75t_L g4826 ( 
.A(n_4529),
.B(n_4504),
.Y(n_4826)
);

O2A1O1Ixp33_ASAP7_75t_SL g4827 ( 
.A1(n_4465),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_4827)
);

OAI21xp5_ASAP7_75t_L g4828 ( 
.A1(n_4444),
.A2(n_1969),
.B(n_1968),
.Y(n_4828)
);

CKINVDCx6p67_ASAP7_75t_R g4829 ( 
.A(n_4299),
.Y(n_4829)
);

OAI22x1_ASAP7_75t_L g4830 ( 
.A1(n_4431),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_4830)
);

NAND2xp5_ASAP7_75t_SL g4831 ( 
.A(n_4249),
.B(n_1873),
.Y(n_4831)
);

INVx2_ASAP7_75t_L g4832 ( 
.A(n_4212),
.Y(n_4832)
);

A2O1A1Ixp33_ASAP7_75t_L g4833 ( 
.A1(n_4444),
.A2(n_4403),
.B(n_4520),
.C(n_4409),
.Y(n_4833)
);

O2A1O1Ixp33_ASAP7_75t_SL g4834 ( 
.A1(n_4225),
.A2(n_21),
.B(n_17),
.C(n_20),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_SL g4835 ( 
.A(n_4249),
.B(n_1873),
.Y(n_4835)
);

AO31x2_ASAP7_75t_L g4836 ( 
.A1(n_4337),
.A2(n_1969),
.A3(n_1978),
.B(n_1968),
.Y(n_4836)
);

CKINVDCx8_ASAP7_75t_R g4837 ( 
.A(n_4207),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_4452),
.Y(n_4838)
);

CKINVDCx16_ASAP7_75t_R g4839 ( 
.A(n_4477),
.Y(n_4839)
);

BUFx3_ASAP7_75t_L g4840 ( 
.A(n_4306),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_4451),
.B(n_65),
.Y(n_4841)
);

AOI21xp5_ASAP7_75t_L g4842 ( 
.A1(n_4481),
.A2(n_2815),
.B(n_2756),
.Y(n_4842)
);

A2O1A1Ixp33_ASAP7_75t_L g4843 ( 
.A1(n_4409),
.A2(n_68),
.B(n_69),
.C(n_65),
.Y(n_4843)
);

A2O1A1Ixp33_ASAP7_75t_L g4844 ( 
.A1(n_4301),
.A2(n_71),
.B(n_72),
.C(n_70),
.Y(n_4844)
);

AO31x2_ASAP7_75t_L g4845 ( 
.A1(n_4337),
.A2(n_1980),
.A3(n_1990),
.B(n_1978),
.Y(n_4845)
);

O2A1O1Ixp33_ASAP7_75t_SL g4846 ( 
.A1(n_4225),
.A2(n_23),
.B(n_20),
.C(n_22),
.Y(n_4846)
);

A2O1A1Ixp33_ASAP7_75t_L g4847 ( 
.A1(n_4305),
.A2(n_73),
.B(n_74),
.C(n_71),
.Y(n_4847)
);

NOR2xp33_ASAP7_75t_L g4848 ( 
.A(n_4348),
.B(n_73),
.Y(n_4848)
);

AOI21xp5_ASAP7_75t_L g4849 ( 
.A1(n_4481),
.A2(n_3061),
.B(n_2815),
.Y(n_4849)
);

NOR2xp33_ASAP7_75t_L g4850 ( 
.A(n_4260),
.B(n_74),
.Y(n_4850)
);

AOI22xp33_ASAP7_75t_L g4851 ( 
.A1(n_4445),
.A2(n_2995),
.B1(n_3033),
.B2(n_2992),
.Y(n_4851)
);

OAI21xp5_ASAP7_75t_L g4852 ( 
.A1(n_4310),
.A2(n_4468),
.B(n_4455),
.Y(n_4852)
);

O2A1O1Ixp5_ASAP7_75t_SL g4853 ( 
.A1(n_4223),
.A2(n_1863),
.B(n_1892),
.C(n_1852),
.Y(n_4853)
);

CKINVDCx5p33_ASAP7_75t_R g4854 ( 
.A(n_4328),
.Y(n_4854)
);

AOI21xp5_ASAP7_75t_L g4855 ( 
.A1(n_4481),
.A2(n_3101),
.B(n_3061),
.Y(n_4855)
);

INVx2_ASAP7_75t_L g4856 ( 
.A(n_4213),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4219),
.Y(n_4857)
);

AND2x4_ASAP7_75t_L g4858 ( 
.A(n_4252),
.B(n_3061),
.Y(n_4858)
);

OAI21x1_ASAP7_75t_L g4859 ( 
.A1(n_4454),
.A2(n_1990),
.B(n_1980),
.Y(n_4859)
);

AOI22xp33_ASAP7_75t_L g4860 ( 
.A1(n_4434),
.A2(n_2995),
.B1(n_3033),
.B2(n_2992),
.Y(n_4860)
);

AOI22xp5_ASAP7_75t_L g4861 ( 
.A1(n_4286),
.A2(n_3101),
.B1(n_2870),
.B2(n_2915),
.Y(n_4861)
);

AOI21xp5_ASAP7_75t_L g4862 ( 
.A1(n_4269),
.A2(n_3101),
.B(n_2302),
.Y(n_4862)
);

OAI22xp5_ASAP7_75t_L g4863 ( 
.A1(n_4233),
.A2(n_2007),
.B1(n_2020),
.B2(n_1995),
.Y(n_4863)
);

A2O1A1Ixp33_ASAP7_75t_L g4864 ( 
.A1(n_4305),
.A2(n_76),
.B(n_79),
.C(n_75),
.Y(n_4864)
);

OAI21xp5_ASAP7_75t_L g4865 ( 
.A1(n_4310),
.A2(n_2007),
.B(n_1995),
.Y(n_4865)
);

A2O1A1Ixp33_ASAP7_75t_L g4866 ( 
.A1(n_4315),
.A2(n_80),
.B(n_81),
.C(n_75),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4350),
.B(n_80),
.Y(n_4867)
);

OAI21x1_ASAP7_75t_L g4868 ( 
.A1(n_4454),
.A2(n_2026),
.B(n_2024),
.Y(n_4868)
);

OAI21x1_ASAP7_75t_L g4869 ( 
.A1(n_4455),
.A2(n_2028),
.B(n_2026),
.Y(n_4869)
);

AOI22xp33_ASAP7_75t_L g4870 ( 
.A1(n_4567),
.A2(n_4440),
.B1(n_4460),
.B2(n_4456),
.Y(n_4870)
);

AND2x4_ASAP7_75t_L g4871 ( 
.A(n_4784),
.B(n_4294),
.Y(n_4871)
);

INVx2_ASAP7_75t_L g4872 ( 
.A(n_4821),
.Y(n_4872)
);

AND2x2_ASAP7_75t_L g4873 ( 
.A(n_4822),
.B(n_4434),
.Y(n_4873)
);

INVxp67_ASAP7_75t_L g4874 ( 
.A(n_4718),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4558),
.Y(n_4875)
);

BUFx6f_ASAP7_75t_L g4876 ( 
.A(n_4804),
.Y(n_4876)
);

CKINVDCx6p67_ASAP7_75t_R g4877 ( 
.A(n_4639),
.Y(n_4877)
);

AOI22xp33_ASAP7_75t_L g4878 ( 
.A1(n_4571),
.A2(n_4456),
.B1(n_4460),
.B2(n_4440),
.Y(n_4878)
);

INVx1_ASAP7_75t_SL g4879 ( 
.A(n_4626),
.Y(n_4879)
);

INVx8_ASAP7_75t_L g4880 ( 
.A(n_4678),
.Y(n_4880)
);

AND2x2_ASAP7_75t_L g4881 ( 
.A(n_4735),
.B(n_4808),
.Y(n_4881)
);

CKINVDCx20_ASAP7_75t_R g4882 ( 
.A(n_4643),
.Y(n_4882)
);

OAI221xp5_ASAP7_75t_L g4883 ( 
.A1(n_4569),
.A2(n_4269),
.B1(n_4230),
.B2(n_4238),
.C(n_4234),
.Y(n_4883)
);

OAI221xp5_ASAP7_75t_L g4884 ( 
.A1(n_4556),
.A2(n_4607),
.B1(n_4716),
.B2(n_4750),
.C(n_4577),
.Y(n_4884)
);

INVx1_ASAP7_75t_SL g4885 ( 
.A(n_4764),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4559),
.Y(n_4886)
);

AOI22xp33_ASAP7_75t_L g4887 ( 
.A1(n_4601),
.A2(n_4526),
.B1(n_4294),
.B2(n_4433),
.Y(n_4887)
);

AOI22xp33_ASAP7_75t_L g4888 ( 
.A1(n_4551),
.A2(n_4526),
.B1(n_4294),
.B2(n_4439),
.Y(n_4888)
);

OAI22xp33_ASAP7_75t_L g4889 ( 
.A1(n_4548),
.A2(n_4389),
.B1(n_4392),
.B2(n_4522),
.Y(n_4889)
);

AND2x2_ASAP7_75t_L g4890 ( 
.A(n_4811),
.B(n_4362),
.Y(n_4890)
);

AOI22xp33_ASAP7_75t_SL g4891 ( 
.A1(n_4779),
.A2(n_4522),
.B1(n_4327),
.B2(n_4362),
.Y(n_4891)
);

O2A1O1Ixp33_ASAP7_75t_L g4892 ( 
.A1(n_4843),
.A2(n_4275),
.B(n_4396),
.C(n_4399),
.Y(n_4892)
);

AOI22xp33_ASAP7_75t_L g4893 ( 
.A1(n_4694),
.A2(n_4429),
.B1(n_4286),
.B2(n_4296),
.Y(n_4893)
);

OR2x6_ASAP7_75t_L g4894 ( 
.A(n_4784),
.B(n_4389),
.Y(n_4894)
);

BUFx2_ASAP7_75t_L g4895 ( 
.A(n_4561),
.Y(n_4895)
);

NOR2xp33_ASAP7_75t_L g4896 ( 
.A(n_4839),
.B(n_4757),
.Y(n_4896)
);

OAI22xp5_ASAP7_75t_L g4897 ( 
.A1(n_4575),
.A2(n_4327),
.B1(n_4396),
.B2(n_4461),
.Y(n_4897)
);

BUFx12f_ASAP7_75t_L g4898 ( 
.A(n_4553),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4654),
.B(n_4522),
.Y(n_4899)
);

AO21x2_ASAP7_75t_L g4900 ( 
.A1(n_4810),
.A2(n_4767),
.B(n_4752),
.Y(n_4900)
);

AOI22xp33_ASAP7_75t_L g4901 ( 
.A1(n_4642),
.A2(n_4355),
.B1(n_4370),
.B2(n_4503),
.Y(n_4901)
);

BUFx12f_ASAP7_75t_L g4902 ( 
.A(n_4656),
.Y(n_4902)
);

AOI22xp33_ASAP7_75t_L g4903 ( 
.A1(n_4669),
.A2(n_4370),
.B1(n_4503),
.B2(n_4275),
.Y(n_4903)
);

AOI22xp33_ASAP7_75t_L g4904 ( 
.A1(n_4580),
.A2(n_4372),
.B1(n_4361),
.B2(n_4507),
.Y(n_4904)
);

NOR2xp67_ASAP7_75t_L g4905 ( 
.A(n_4753),
.B(n_4717),
.Y(n_4905)
);

AOI22xp5_ASAP7_75t_L g4906 ( 
.A1(n_4671),
.A2(n_4504),
.B1(n_4406),
.B2(n_4228),
.Y(n_4906)
);

AOI22xp33_ASAP7_75t_L g4907 ( 
.A1(n_4586),
.A2(n_4798),
.B1(n_4621),
.B2(n_4700),
.Y(n_4907)
);

INVx2_ASAP7_75t_L g4908 ( 
.A(n_4549),
.Y(n_4908)
);

OAI22xp5_ASAP7_75t_L g4909 ( 
.A1(n_4844),
.A2(n_4327),
.B1(n_4461),
.B2(n_4352),
.Y(n_4909)
);

AOI21xp5_ASAP7_75t_L g4910 ( 
.A1(n_4557),
.A2(n_4368),
.B(n_4398),
.Y(n_4910)
);

OAI22xp33_ASAP7_75t_L g4911 ( 
.A1(n_4653),
.A2(n_4350),
.B1(n_4373),
.B2(n_4352),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_L g4912 ( 
.A(n_4612),
.B(n_4417),
.Y(n_4912)
);

OAI22xp33_ASAP7_75t_L g4913 ( 
.A1(n_4615),
.A2(n_4820),
.B1(n_4830),
.B2(n_4861),
.Y(n_4913)
);

AOI22xp33_ASAP7_75t_L g4914 ( 
.A1(n_4759),
.A2(n_4441),
.B1(n_4415),
.B2(n_4517),
.Y(n_4914)
);

AND2x4_ASAP7_75t_L g4915 ( 
.A(n_4561),
.B(n_4532),
.Y(n_4915)
);

AND2x2_ASAP7_75t_L g4916 ( 
.A(n_4760),
.B(n_4404),
.Y(n_4916)
);

OAI22xp5_ASAP7_75t_L g4917 ( 
.A1(n_4847),
.A2(n_4373),
.B1(n_4430),
.B2(n_4417),
.Y(n_4917)
);

AND2x4_ASAP7_75t_L g4918 ( 
.A(n_4797),
.B(n_4815),
.Y(n_4918)
);

AND2x2_ASAP7_75t_L g4919 ( 
.A(n_4550),
.B(n_4479),
.Y(n_4919)
);

AND2x6_ASAP7_75t_L g4920 ( 
.A(n_4858),
.B(n_4458),
.Y(n_4920)
);

INVx2_ASAP7_75t_L g4921 ( 
.A(n_4564),
.Y(n_4921)
);

NAND3xp33_ASAP7_75t_L g4922 ( 
.A(n_4582),
.B(n_4496),
.C(n_4430),
.Y(n_4922)
);

AOI21xp5_ASAP7_75t_L g4923 ( 
.A1(n_4562),
.A2(n_4368),
.B(n_4398),
.Y(n_4923)
);

AOI22xp33_ASAP7_75t_L g4924 ( 
.A1(n_4823),
.A2(n_4499),
.B1(n_4228),
.B2(n_4231),
.Y(n_4924)
);

OR2x2_ASAP7_75t_L g4925 ( 
.A(n_4838),
.B(n_4276),
.Y(n_4925)
);

INVx2_ASAP7_75t_L g4926 ( 
.A(n_4597),
.Y(n_4926)
);

AO21x2_ASAP7_75t_L g4927 ( 
.A1(n_4748),
.A2(n_4625),
.B(n_4616),
.Y(n_4927)
);

AOI22xp33_ASAP7_75t_L g4928 ( 
.A1(n_4763),
.A2(n_4231),
.B1(n_4215),
.B2(n_4375),
.Y(n_4928)
);

BUFx10_ASAP7_75t_L g4929 ( 
.A(n_4678),
.Y(n_4929)
);

INVxp67_ASAP7_75t_L g4930 ( 
.A(n_4660),
.Y(n_4930)
);

O2A1O1Ixp33_ASAP7_75t_L g4931 ( 
.A1(n_4864),
.A2(n_4485),
.B(n_4333),
.C(n_4279),
.Y(n_4931)
);

NAND2x1p5_ASAP7_75t_L g4932 ( 
.A(n_4824),
.B(n_4467),
.Y(n_4932)
);

AOI22xp5_ASAP7_75t_L g4933 ( 
.A1(n_4552),
.A2(n_4406),
.B1(n_4215),
.B2(n_4458),
.Y(n_4933)
);

BUFx6f_ASAP7_75t_L g4934 ( 
.A(n_4678),
.Y(n_4934)
);

AOI22xp33_ASAP7_75t_L g4935 ( 
.A1(n_4603),
.A2(n_4384),
.B1(n_4321),
.B2(n_4324),
.Y(n_4935)
);

OAI22xp5_ASAP7_75t_L g4936 ( 
.A1(n_4866),
.A2(n_4365),
.B1(n_4412),
.B2(n_4347),
.Y(n_4936)
);

OAI22xp33_ASAP7_75t_SL g4937 ( 
.A1(n_4782),
.A2(n_4427),
.B1(n_4307),
.B2(n_4351),
.Y(n_4937)
);

OAI22xp5_ASAP7_75t_L g4938 ( 
.A1(n_4600),
.A2(n_4485),
.B1(n_4315),
.B2(n_4427),
.Y(n_4938)
);

NOR2xp67_ASAP7_75t_SL g4939 ( 
.A(n_4729),
.B(n_4467),
.Y(n_4939)
);

CKINVDCx20_ASAP7_75t_R g4940 ( 
.A(n_4647),
.Y(n_4940)
);

AOI22xp33_ASAP7_75t_L g4941 ( 
.A1(n_4736),
.A2(n_4756),
.B1(n_4749),
.B2(n_4587),
.Y(n_4941)
);

OR2x2_ASAP7_75t_L g4942 ( 
.A(n_4769),
.B(n_4359),
.Y(n_4942)
);

INVx1_ASAP7_75t_L g4943 ( 
.A(n_4570),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4599),
.B(n_4367),
.Y(n_4944)
);

OAI21xp5_ASAP7_75t_L g4945 ( 
.A1(n_4605),
.A2(n_4343),
.B(n_4467),
.Y(n_4945)
);

AOI22xp33_ASAP7_75t_SL g4946 ( 
.A1(n_4676),
.A2(n_4427),
.B1(n_4467),
.B2(n_4343),
.Y(n_4946)
);

NAND2x1p5_ASAP7_75t_L g4947 ( 
.A(n_4565),
.B(n_4480),
.Y(n_4947)
);

INVx3_ASAP7_75t_L g4948 ( 
.A(n_4737),
.Y(n_4948)
);

INVx4_ASAP7_75t_L g4949 ( 
.A(n_4677),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4572),
.Y(n_4950)
);

INVx2_ASAP7_75t_SL g4951 ( 
.A(n_4602),
.Y(n_4951)
);

INVx3_ASAP7_75t_SL g4952 ( 
.A(n_4631),
.Y(n_4952)
);

OAI222xp33_ASAP7_75t_L g4953 ( 
.A1(n_4867),
.A2(n_4258),
.B1(n_4308),
.B2(n_4374),
.C1(n_4383),
.C2(n_4369),
.Y(n_4953)
);

AND2x4_ASAP7_75t_L g4954 ( 
.A(n_4726),
.B(n_4290),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4614),
.Y(n_4955)
);

AOI22xp33_ASAP7_75t_L g4956 ( 
.A1(n_4848),
.A2(n_4239),
.B1(n_4241),
.B2(n_4237),
.Y(n_4956)
);

CKINVDCx11_ASAP7_75t_R g4957 ( 
.A(n_4684),
.Y(n_4957)
);

AND2x4_ASAP7_75t_L g4958 ( 
.A(n_4648),
.B(n_4291),
.Y(n_4958)
);

OAI22xp5_ASAP7_75t_L g4959 ( 
.A1(n_4806),
.A2(n_4505),
.B1(n_4413),
.B2(n_4303),
.Y(n_4959)
);

INVx2_ASAP7_75t_L g4960 ( 
.A(n_4604),
.Y(n_4960)
);

AOI21xp5_ASAP7_75t_L g4961 ( 
.A1(n_4563),
.A2(n_4222),
.B(n_4413),
.Y(n_4961)
);

OR2x2_ASAP7_75t_L g4962 ( 
.A(n_4741),
.B(n_4505),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4623),
.Y(n_4963)
);

INVx6_ASAP7_75t_L g4964 ( 
.A(n_4677),
.Y(n_4964)
);

HB1xp67_ASAP7_75t_L g4965 ( 
.A(n_4619),
.Y(n_4965)
);

NAND2xp5_ASAP7_75t_L g4966 ( 
.A(n_4576),
.B(n_4303),
.Y(n_4966)
);

INVx4_ASAP7_75t_L g4967 ( 
.A(n_4737),
.Y(n_4967)
);

AOI22xp33_ASAP7_75t_L g4968 ( 
.A1(n_4807),
.A2(n_4239),
.B1(n_4241),
.B2(n_4237),
.Y(n_4968)
);

OAI22xp5_ASAP7_75t_L g4969 ( 
.A1(n_4733),
.A2(n_4320),
.B1(n_4330),
.B2(n_4304),
.Y(n_4969)
);

NOR2x1_ASAP7_75t_SL g4970 ( 
.A(n_4615),
.B(n_4237),
.Y(n_4970)
);

OAI22xp5_ASAP7_75t_L g4971 ( 
.A1(n_4738),
.A2(n_4751),
.B1(n_4680),
.B2(n_4833),
.Y(n_4971)
);

O2A1O1Ixp33_ASAP7_75t_L g4972 ( 
.A1(n_4663),
.A2(n_4320),
.B(n_4330),
.C(n_4304),
.Y(n_4972)
);

AOI21xp5_ASAP7_75t_L g4973 ( 
.A1(n_4765),
.A2(n_4414),
.B(n_4400),
.Y(n_4973)
);

INVx2_ASAP7_75t_L g4974 ( 
.A(n_4630),
.Y(n_4974)
);

AOI22xp33_ASAP7_75t_L g4975 ( 
.A1(n_4687),
.A2(n_4295),
.B1(n_4241),
.B2(n_4346),
.Y(n_4975)
);

AOI22xp33_ASAP7_75t_L g4976 ( 
.A1(n_4574),
.A2(n_4295),
.B1(n_4358),
.B2(n_4357),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4721),
.B(n_4340),
.Y(n_4977)
);

AOI22xp5_ASAP7_75t_L g4978 ( 
.A1(n_4555),
.A2(n_4295),
.B1(n_4421),
.B2(n_4340),
.Y(n_4978)
);

A2O1A1Ixp33_ASAP7_75t_L g4979 ( 
.A1(n_4596),
.A2(n_4792),
.B(n_4714),
.C(n_4590),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4636),
.Y(n_4980)
);

INVx3_ASAP7_75t_L g4981 ( 
.A(n_4826),
.Y(n_4981)
);

INVx2_ASAP7_75t_L g4982 ( 
.A(n_4658),
.Y(n_4982)
);

INVx2_ASAP7_75t_SL g4983 ( 
.A(n_4602),
.Y(n_4983)
);

AOI221xp5_ASAP7_75t_L g4984 ( 
.A1(n_4827),
.A2(n_4846),
.B1(n_4834),
.B2(n_4689),
.C(n_4667),
.Y(n_4984)
);

AOI22xp33_ASAP7_75t_L g4985 ( 
.A1(n_4566),
.A2(n_4421),
.B1(n_4340),
.B2(n_2870),
.Y(n_4985)
);

INVx2_ASAP7_75t_L g4986 ( 
.A(n_4690),
.Y(n_4986)
);

NAND2x1_ASAP7_75t_L g4987 ( 
.A(n_4776),
.B(n_2852),
.Y(n_4987)
);

OR2x2_ASAP7_75t_L g4988 ( 
.A(n_4741),
.B(n_83),
.Y(n_4988)
);

INVx1_ASAP7_75t_SL g4989 ( 
.A(n_4695),
.Y(n_4989)
);

AOI22xp5_ASAP7_75t_L g4990 ( 
.A1(n_4850),
.A2(n_2870),
.B1(n_2915),
.B2(n_2852),
.Y(n_4990)
);

OAI22xp33_ASAP7_75t_L g4991 ( 
.A1(n_4588),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4697),
.Y(n_4992)
);

NOR2xp67_ASAP7_75t_SL g4993 ( 
.A(n_4837),
.B(n_1864),
.Y(n_4993)
);

INVx6_ASAP7_75t_L g4994 ( 
.A(n_4578),
.Y(n_4994)
);

NAND2xp5_ASAP7_75t_L g4995 ( 
.A(n_4772),
.B(n_84),
.Y(n_4995)
);

INVx1_ASAP7_75t_SL g4996 ( 
.A(n_4673),
.Y(n_4996)
);

INVx2_ASAP7_75t_L g4997 ( 
.A(n_4702),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4703),
.Y(n_4998)
);

INVx2_ASAP7_75t_L g4999 ( 
.A(n_4857),
.Y(n_4999)
);

OAI221xp5_ASAP7_75t_L g5000 ( 
.A1(n_4608),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.C(n_26),
.Y(n_5000)
);

AOI22xp33_ASAP7_75t_L g5001 ( 
.A1(n_4724),
.A2(n_2870),
.B1(n_2915),
.B2(n_2852),
.Y(n_5001)
);

AOI22xp33_ASAP7_75t_L g5002 ( 
.A1(n_4617),
.A2(n_2870),
.B1(n_2915),
.B2(n_2852),
.Y(n_5002)
);

AOI22xp33_ASAP7_75t_SL g5003 ( 
.A1(n_4672),
.A2(n_2870),
.B1(n_2915),
.B2(n_2852),
.Y(n_5003)
);

AOI22xp33_ASAP7_75t_L g5004 ( 
.A1(n_4641),
.A2(n_2915),
.B1(n_1876),
.B2(n_1885),
.Y(n_5004)
);

OAI21xp5_ASAP7_75t_L g5005 ( 
.A1(n_4649),
.A2(n_2032),
.B(n_2028),
.Y(n_5005)
);

AOI22xp33_ASAP7_75t_L g5006 ( 
.A1(n_4638),
.A2(n_1876),
.B1(n_1885),
.B2(n_1868),
.Y(n_5006)
);

OR2x6_ASAP7_75t_L g5007 ( 
.A(n_4747),
.B(n_2271),
.Y(n_5007)
);

CKINVDCx11_ASAP7_75t_R g5008 ( 
.A(n_4829),
.Y(n_5008)
);

OAI22xp5_ASAP7_75t_L g5009 ( 
.A1(n_4722),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_5009)
);

INVx2_ASAP7_75t_SL g5010 ( 
.A(n_4840),
.Y(n_5010)
);

AND2x4_ASAP7_75t_L g5011 ( 
.A(n_4568),
.B(n_86),
.Y(n_5011)
);

OAI21x1_ASAP7_75t_L g5012 ( 
.A1(n_4646),
.A2(n_2054),
.B(n_2032),
.Y(n_5012)
);

INVx2_ASAP7_75t_L g5013 ( 
.A(n_4832),
.Y(n_5013)
);

AND2x4_ASAP7_75t_L g5014 ( 
.A(n_4568),
.B(n_87),
.Y(n_5014)
);

INVx2_ASAP7_75t_L g5015 ( 
.A(n_4856),
.Y(n_5015)
);

OAI21xp5_ASAP7_75t_L g5016 ( 
.A1(n_4778),
.A2(n_2055),
.B(n_2054),
.Y(n_5016)
);

AND2x4_ASAP7_75t_L g5017 ( 
.A(n_4789),
.B(n_87),
.Y(n_5017)
);

OR2x6_ASAP7_75t_L g5018 ( 
.A(n_4739),
.B(n_2293),
.Y(n_5018)
);

AND2x4_ASAP7_75t_L g5019 ( 
.A(n_4793),
.B(n_88),
.Y(n_5019)
);

AOI22xp33_ASAP7_75t_L g5020 ( 
.A1(n_4685),
.A2(n_1887),
.B1(n_1888),
.B2(n_1868),
.Y(n_5020)
);

HB1xp67_ASAP7_75t_L g5021 ( 
.A(n_4741),
.Y(n_5021)
);

AOI22xp33_ASAP7_75t_L g5022 ( 
.A1(n_4609),
.A2(n_4699),
.B1(n_4818),
.B2(n_4852),
.Y(n_5022)
);

AOI22xp33_ASAP7_75t_L g5023 ( 
.A1(n_4858),
.A2(n_1888),
.B1(n_1896),
.B2(n_1887),
.Y(n_5023)
);

OAI22xp5_ASAP7_75t_L g5024 ( 
.A1(n_4683),
.A2(n_28),
.B1(n_25),
.B2(n_27),
.Y(n_5024)
);

INVx2_ASAP7_75t_L g5025 ( 
.A(n_4799),
.Y(n_5025)
);

NAND2x1p5_ASAP7_75t_L g5026 ( 
.A(n_4665),
.B(n_4713),
.Y(n_5026)
);

O2A1O1Ixp33_ASAP7_75t_L g5027 ( 
.A1(n_4560),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_5027)
);

INVx2_ASAP7_75t_L g5028 ( 
.A(n_4802),
.Y(n_5028)
);

OAI21xp5_ASAP7_75t_L g5029 ( 
.A1(n_4743),
.A2(n_2061),
.B(n_2060),
.Y(n_5029)
);

AND2x6_ASAP7_75t_L g5030 ( 
.A(n_4774),
.B(n_1896),
.Y(n_5030)
);

OR2x2_ASAP7_75t_L g5031 ( 
.A(n_4813),
.B(n_89),
.Y(n_5031)
);

AOI22xp33_ASAP7_75t_SL g5032 ( 
.A1(n_4622),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_5032)
);

AOI22xp33_ASAP7_75t_L g5033 ( 
.A1(n_4819),
.A2(n_2079),
.B1(n_2082),
.B2(n_2061),
.Y(n_5033)
);

BUFx3_ASAP7_75t_L g5034 ( 
.A(n_4854),
.Y(n_5034)
);

INVx3_ASAP7_75t_L g5035 ( 
.A(n_4554),
.Y(n_5035)
);

BUFx12f_ASAP7_75t_L g5036 ( 
.A(n_4645),
.Y(n_5036)
);

BUFx6f_ASAP7_75t_L g5037 ( 
.A(n_4773),
.Y(n_5037)
);

OR2x2_ASAP7_75t_L g5038 ( 
.A(n_4606),
.B(n_90),
.Y(n_5038)
);

INVxp67_ASAP7_75t_SL g5039 ( 
.A(n_4809),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_4670),
.B(n_4620),
.Y(n_5040)
);

OR2x2_ASAP7_75t_L g5041 ( 
.A(n_4606),
.B(n_90),
.Y(n_5041)
);

O2A1O1Ixp33_ASAP7_75t_SL g5042 ( 
.A1(n_4768),
.A2(n_92),
.B(n_94),
.C(n_91),
.Y(n_5042)
);

INVx2_ASAP7_75t_L g5043 ( 
.A(n_4644),
.Y(n_5043)
);

AOI22xp33_ASAP7_75t_SL g5044 ( 
.A1(n_4613),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_5044)
);

INVx8_ASAP7_75t_L g5045 ( 
.A(n_4773),
.Y(n_5045)
);

AOI22xp5_ASAP7_75t_L g5046 ( 
.A1(n_4651),
.A2(n_2082),
.B1(n_2090),
.B2(n_2079),
.Y(n_5046)
);

NOR2xp33_ASAP7_75t_L g5047 ( 
.A(n_4637),
.B(n_94),
.Y(n_5047)
);

AOI22xp33_ASAP7_75t_L g5048 ( 
.A1(n_4659),
.A2(n_2096),
.B1(n_2106),
.B2(n_2090),
.Y(n_5048)
);

NAND2xp5_ASAP7_75t_L g5049 ( 
.A(n_4791),
.B(n_95),
.Y(n_5049)
);

CKINVDCx5p33_ASAP7_75t_R g5050 ( 
.A(n_4633),
.Y(n_5050)
);

NAND2xp5_ASAP7_75t_L g5051 ( 
.A(n_4788),
.B(n_97),
.Y(n_5051)
);

CKINVDCx20_ASAP7_75t_R g5052 ( 
.A(n_4712),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4606),
.Y(n_5053)
);

OAI22xp33_ASAP7_75t_L g5054 ( 
.A1(n_4794),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_5054)
);

OAI22xp5_ASAP7_75t_L g5055 ( 
.A1(n_4711),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_5055)
);

AOI221xp5_ASAP7_75t_L g5056 ( 
.A1(n_4707),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.C(n_39),
.Y(n_5056)
);

OA21x2_ASAP7_75t_L g5057 ( 
.A1(n_4686),
.A2(n_2106),
.B(n_2096),
.Y(n_5057)
);

NAND2x1p5_ASAP7_75t_L g5058 ( 
.A(n_4725),
.B(n_2108),
.Y(n_5058)
);

OR2x2_ASAP7_75t_L g5059 ( 
.A(n_4644),
.B(n_97),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_SL g5060 ( 
.A(n_4652),
.B(n_1842),
.Y(n_5060)
);

OAI22xp5_ASAP7_75t_L g5061 ( 
.A1(n_4801),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_5061)
);

AOI22xp33_ASAP7_75t_L g5062 ( 
.A1(n_4771),
.A2(n_2126),
.B1(n_2131),
.B2(n_2120),
.Y(n_5062)
);

CKINVDCx5p33_ASAP7_75t_R g5063 ( 
.A(n_4674),
.Y(n_5063)
);

AO32x2_ASAP7_75t_L g5064 ( 
.A1(n_4554),
.A2(n_42),
.A3(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_5064)
);

AOI22xp33_ASAP7_75t_SL g5065 ( 
.A1(n_4629),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_5065)
);

OAI22xp5_ASAP7_75t_L g5066 ( 
.A1(n_4814),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_5066)
);

AOI21xp33_ASAP7_75t_L g5067 ( 
.A1(n_4745),
.A2(n_43),
.B(n_44),
.Y(n_5067)
);

AOI22xp33_ASAP7_75t_L g5068 ( 
.A1(n_4754),
.A2(n_2131),
.B1(n_2135),
.B2(n_2126),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_L g5069 ( 
.A(n_4705),
.B(n_44),
.Y(n_5069)
);

AND2x2_ASAP7_75t_L g5070 ( 
.A(n_4715),
.B(n_98),
.Y(n_5070)
);

OAI22xp5_ASAP7_75t_L g5071 ( 
.A1(n_4841),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_4710),
.B(n_46),
.Y(n_5072)
);

INVx2_ASAP7_75t_L g5073 ( 
.A(n_4661),
.Y(n_5073)
);

AND2x4_ASAP7_75t_L g5074 ( 
.A(n_4715),
.B(n_100),
.Y(n_5074)
);

AND2x2_ASAP7_75t_L g5075 ( 
.A(n_4727),
.B(n_101),
.Y(n_5075)
);

AND2x2_ASAP7_75t_L g5076 ( 
.A(n_4727),
.B(n_102),
.Y(n_5076)
);

OAI22xp5_ASAP7_75t_L g5077 ( 
.A1(n_4618),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_5077)
);

OAI22xp33_ASAP7_75t_L g5078 ( 
.A1(n_4668),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_5078)
);

OAI221xp5_ASAP7_75t_L g5079 ( 
.A1(n_4770),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.C(n_53),
.Y(n_5079)
);

AOI22xp33_ASAP7_75t_L g5080 ( 
.A1(n_4831),
.A2(n_2138),
.B1(n_2139),
.B2(n_2136),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_4816),
.Y(n_5081)
);

AND2x2_ASAP7_75t_L g5082 ( 
.A(n_4666),
.B(n_102),
.Y(n_5082)
);

INVx2_ASAP7_75t_L g5083 ( 
.A(n_4661),
.Y(n_5083)
);

OAI22xp5_ASAP7_75t_L g5084 ( 
.A1(n_4679),
.A2(n_51),
.B1(n_54),
.B2(n_113),
.Y(n_5084)
);

OAI22xp5_ASAP7_75t_L g5085 ( 
.A1(n_4679),
.A2(n_51),
.B1(n_54),
.B2(n_113),
.Y(n_5085)
);

OAI22xp5_ASAP7_75t_L g5086 ( 
.A1(n_4679),
.A2(n_117),
.B1(n_127),
.B2(n_104),
.Y(n_5086)
);

AOI22xp33_ASAP7_75t_L g5087 ( 
.A1(n_4835),
.A2(n_2146),
.B1(n_2150),
.B2(n_2139),
.Y(n_5087)
);

BUFx2_ASAP7_75t_L g5088 ( 
.A(n_4712),
.Y(n_5088)
);

OAI22xp5_ASAP7_75t_L g5089 ( 
.A1(n_4691),
.A2(n_117),
.B1(n_127),
.B2(n_104),
.Y(n_5089)
);

OAI22xp5_ASAP7_75t_L g5090 ( 
.A1(n_4691),
.A2(n_119),
.B1(n_130),
.B2(n_106),
.Y(n_5090)
);

OAI22xp33_ASAP7_75t_L g5091 ( 
.A1(n_4730),
.A2(n_2164),
.B1(n_2165),
.B2(n_2160),
.Y(n_5091)
);

CKINVDCx5p33_ASAP7_75t_R g5092 ( 
.A(n_4692),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4816),
.Y(n_5093)
);

OAI22xp5_ASAP7_75t_L g5094 ( 
.A1(n_4691),
.A2(n_120),
.B1(n_131),
.B2(n_107),
.Y(n_5094)
);

INVx6_ASAP7_75t_L g5095 ( 
.A(n_4774),
.Y(n_5095)
);

AOI21xp5_ASAP7_75t_L g5096 ( 
.A1(n_4628),
.A2(n_4634),
.B(n_4595),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_4816),
.Y(n_5097)
);

AOI221xp5_ASAP7_75t_L g5098 ( 
.A1(n_4662),
.A2(n_110),
.B1(n_107),
.B2(n_108),
.C(n_112),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_4777),
.Y(n_5099)
);

INVx2_ASAP7_75t_L g5100 ( 
.A(n_4859),
.Y(n_5100)
);

BUFx2_ASAP7_75t_L g5101 ( 
.A(n_4632),
.Y(n_5101)
);

A2O1A1Ixp33_ASAP7_75t_L g5102 ( 
.A1(n_4650),
.A2(n_118),
.B(n_115),
.C(n_116),
.Y(n_5102)
);

OAI222xp33_ASAP7_75t_L g5103 ( 
.A1(n_4782),
.A2(n_119),
.B1(n_123),
.B2(n_116),
.C1(n_118),
.C2(n_121),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_4777),
.Y(n_5104)
);

INVx2_ASAP7_75t_SL g5105 ( 
.A(n_4825),
.Y(n_5105)
);

AOI221xp5_ASAP7_75t_L g5106 ( 
.A1(n_4664),
.A2(n_126),
.B1(n_123),
.B2(n_124),
.C(n_128),
.Y(n_5106)
);

AOI22xp33_ASAP7_75t_L g5107 ( 
.A1(n_4761),
.A2(n_2185),
.B1(n_2196),
.B2(n_2183),
.Y(n_5107)
);

OAI22xp5_ASAP7_75t_L g5108 ( 
.A1(n_4766),
.A2(n_136),
.B1(n_145),
.B2(n_124),
.Y(n_5108)
);

AOI22xp33_ASAP7_75t_L g5109 ( 
.A1(n_4657),
.A2(n_2196),
.B1(n_2208),
.B2(n_2203),
.Y(n_5109)
);

AOI31xp67_ASAP7_75t_L g5110 ( 
.A1(n_4708),
.A2(n_2208),
.A3(n_2219),
.B(n_2203),
.Y(n_5110)
);

OAI221xp5_ASAP7_75t_L g5111 ( 
.A1(n_4720),
.A2(n_130),
.B1(n_126),
.B2(n_129),
.C(n_131),
.Y(n_5111)
);

OAI222xp33_ASAP7_75t_L g5112 ( 
.A1(n_4782),
.A2(n_134),
.B1(n_138),
.B2(n_132),
.C1(n_133),
.C2(n_137),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_4758),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_4758),
.Y(n_5114)
);

AND2x4_ASAP7_75t_L g5115 ( 
.A(n_4868),
.B(n_138),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_4758),
.Y(n_5116)
);

AOI22xp33_ASAP7_75t_L g5117 ( 
.A1(n_4740),
.A2(n_2219),
.B1(n_2234),
.B2(n_2224),
.Y(n_5117)
);

INVx2_ASAP7_75t_SL g5118 ( 
.A(n_4780),
.Y(n_5118)
);

HB1xp67_ASAP7_75t_L g5119 ( 
.A(n_4719),
.Y(n_5119)
);

NOR2xp33_ASAP7_75t_L g5120 ( 
.A(n_4796),
.B(n_139),
.Y(n_5120)
);

INVx2_ASAP7_75t_L g5121 ( 
.A(n_4869),
.Y(n_5121)
);

BUFx2_ASAP7_75t_L g5122 ( 
.A(n_4836),
.Y(n_5122)
);

AOI222xp33_ASAP7_75t_L g5123 ( 
.A1(n_4795),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.C1(n_140),
.C2(n_143),
.Y(n_5123)
);

INVx1_ASAP7_75t_L g5124 ( 
.A(n_4635),
.Y(n_5124)
);

NAND2xp5_ASAP7_75t_L g5125 ( 
.A(n_4583),
.B(n_139),
.Y(n_5125)
);

INVx1_ASAP7_75t_SL g5126 ( 
.A(n_4585),
.Y(n_5126)
);

BUFx4f_ASAP7_75t_SL g5127 ( 
.A(n_4581),
.Y(n_5127)
);

AOI22xp33_ASAP7_75t_L g5128 ( 
.A1(n_4828),
.A2(n_2241),
.B1(n_2247),
.B2(n_2246),
.Y(n_5128)
);

OR2x6_ASAP7_75t_L g5129 ( 
.A(n_4803),
.B(n_2269),
.Y(n_5129)
);

AND2x2_ASAP7_75t_L g5130 ( 
.A(n_4573),
.B(n_142),
.Y(n_5130)
);

NAND2xp5_ASAP7_75t_L g5131 ( 
.A(n_4583),
.B(n_143),
.Y(n_5131)
);

INVx2_ASAP7_75t_L g5132 ( 
.A(n_4800),
.Y(n_5132)
);

AOI22xp33_ASAP7_75t_L g5133 ( 
.A1(n_4817),
.A2(n_2241),
.B1(n_2247),
.B2(n_2246),
.Y(n_5133)
);

OAI22xp5_ASAP7_75t_L g5134 ( 
.A1(n_4786),
.A2(n_155),
.B1(n_166),
.B2(n_146),
.Y(n_5134)
);

CKINVDCx5p33_ASAP7_75t_R g5135 ( 
.A(n_4957),
.Y(n_5135)
);

INVx3_ASAP7_75t_L g5136 ( 
.A(n_4967),
.Y(n_5136)
);

OAI21xp5_ASAP7_75t_L g5137 ( 
.A1(n_4884),
.A2(n_4862),
.B(n_4849),
.Y(n_5137)
);

INVx2_ASAP7_75t_L g5138 ( 
.A(n_5025),
.Y(n_5138)
);

OAI21xp5_ASAP7_75t_L g5139 ( 
.A1(n_4971),
.A2(n_4855),
.B(n_4842),
.Y(n_5139)
);

INVx2_ASAP7_75t_L g5140 ( 
.A(n_5028),
.Y(n_5140)
);

OAI21x1_ASAP7_75t_L g5141 ( 
.A1(n_5096),
.A2(n_4812),
.B(n_4785),
.Y(n_5141)
);

NAND4xp25_ASAP7_75t_L g5142 ( 
.A(n_5032),
.B(n_4610),
.C(n_4640),
.D(n_4693),
.Y(n_5142)
);

HB1xp67_ASAP7_75t_L g5143 ( 
.A(n_5021),
.Y(n_5143)
);

INVx2_ASAP7_75t_SL g5144 ( 
.A(n_4948),
.Y(n_5144)
);

AOI22xp33_ASAP7_75t_SL g5145 ( 
.A1(n_5127),
.A2(n_4584),
.B1(n_4781),
.B2(n_4775),
.Y(n_5145)
);

INVx2_ASAP7_75t_L g5146 ( 
.A(n_4872),
.Y(n_5146)
);

AND2x2_ASAP7_75t_L g5147 ( 
.A(n_4881),
.B(n_4589),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_4875),
.Y(n_5148)
);

AOI21x1_ASAP7_75t_L g5149 ( 
.A1(n_5125),
.A2(n_4732),
.B(n_4675),
.Y(n_5149)
);

INVx3_ASAP7_75t_L g5150 ( 
.A(n_4967),
.Y(n_5150)
);

INVx1_ASAP7_75t_SL g5151 ( 
.A(n_4952),
.Y(n_5151)
);

AND2x2_ASAP7_75t_L g5152 ( 
.A(n_4873),
.B(n_4589),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_4886),
.Y(n_5153)
);

INVx2_ASAP7_75t_L g5154 ( 
.A(n_4974),
.Y(n_5154)
);

INVx2_ASAP7_75t_L g5155 ( 
.A(n_4982),
.Y(n_5155)
);

BUFx6f_ASAP7_75t_L g5156 ( 
.A(n_4876),
.Y(n_5156)
);

INVx2_ASAP7_75t_L g5157 ( 
.A(n_4986),
.Y(n_5157)
);

HB1xp67_ASAP7_75t_L g5158 ( 
.A(n_4899),
.Y(n_5158)
);

BUFx2_ASAP7_75t_L g5159 ( 
.A(n_4948),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_4943),
.Y(n_5160)
);

INVx2_ASAP7_75t_L g5161 ( 
.A(n_4997),
.Y(n_5161)
);

HB1xp67_ASAP7_75t_L g5162 ( 
.A(n_4899),
.Y(n_5162)
);

AND2x4_ASAP7_75t_L g5163 ( 
.A(n_4894),
.B(n_4871),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_4950),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_4955),
.Y(n_5165)
);

OAI21x1_ASAP7_75t_L g5166 ( 
.A1(n_4923),
.A2(n_4681),
.B(n_4762),
.Y(n_5166)
);

INVx1_ASAP7_75t_L g5167 ( 
.A(n_4963),
.Y(n_5167)
);

OAI21x1_ASAP7_75t_L g5168 ( 
.A1(n_5012),
.A2(n_4742),
.B(n_4734),
.Y(n_5168)
);

INVx1_ASAP7_75t_L g5169 ( 
.A(n_4980),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_4992),
.Y(n_5170)
);

INVx2_ASAP7_75t_L g5171 ( 
.A(n_4998),
.Y(n_5171)
);

OAI21x1_ASAP7_75t_L g5172 ( 
.A1(n_4910),
.A2(n_4655),
.B(n_4682),
.Y(n_5172)
);

INVx3_ASAP7_75t_L g5173 ( 
.A(n_4918),
.Y(n_5173)
);

AND2x2_ASAP7_75t_L g5174 ( 
.A(n_4895),
.B(n_4592),
.Y(n_5174)
);

OAI22xp5_ASAP7_75t_SL g5175 ( 
.A1(n_5052),
.A2(n_4584),
.B1(n_4860),
.B2(n_4851),
.Y(n_5175)
);

AND2x2_ASAP7_75t_L g5176 ( 
.A(n_4890),
.B(n_4592),
.Y(n_5176)
);

HB1xp67_ASAP7_75t_L g5177 ( 
.A(n_4965),
.Y(n_5177)
);

INVxp67_ASAP7_75t_L g5178 ( 
.A(n_5039),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_4999),
.Y(n_5179)
);

INVx2_ASAP7_75t_L g5180 ( 
.A(n_4942),
.Y(n_5180)
);

INVx2_ASAP7_75t_L g5181 ( 
.A(n_4908),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_4921),
.Y(n_5182)
);

OA21x2_ASAP7_75t_L g5183 ( 
.A1(n_5131),
.A2(n_4783),
.B(n_4790),
.Y(n_5183)
);

BUFx3_ASAP7_75t_L g5184 ( 
.A(n_4876),
.Y(n_5184)
);

AOI21x1_ASAP7_75t_L g5185 ( 
.A1(n_5069),
.A2(n_4611),
.B(n_4598),
.Y(n_5185)
);

INVx2_ASAP7_75t_L g5186 ( 
.A(n_4926),
.Y(n_5186)
);

OAI22xp5_ASAP7_75t_L g5187 ( 
.A1(n_4907),
.A2(n_4805),
.B1(n_4787),
.B2(n_4863),
.Y(n_5187)
);

INVx1_ASAP7_75t_L g5188 ( 
.A(n_4960),
.Y(n_5188)
);

OAI21xp5_ASAP7_75t_L g5189 ( 
.A1(n_4971),
.A2(n_4696),
.B(n_4688),
.Y(n_5189)
);

OR2x2_ASAP7_75t_L g5190 ( 
.A(n_4912),
.B(n_4592),
.Y(n_5190)
);

INVx2_ASAP7_75t_SL g5191 ( 
.A(n_4964),
.Y(n_5191)
);

INVx2_ASAP7_75t_SL g5192 ( 
.A(n_4964),
.Y(n_5192)
);

OAI22xp5_ASAP7_75t_L g5193 ( 
.A1(n_4891),
.A2(n_4746),
.B1(n_4755),
.B2(n_4584),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_5013),
.Y(n_5194)
);

OAI21x1_ASAP7_75t_L g5195 ( 
.A1(n_4973),
.A2(n_4709),
.B(n_4704),
.Y(n_5195)
);

BUFx4f_ASAP7_75t_SL g5196 ( 
.A(n_4898),
.Y(n_5196)
);

BUFx2_ASAP7_75t_L g5197 ( 
.A(n_5035),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_5015),
.Y(n_5198)
);

INVx3_ASAP7_75t_L g5199 ( 
.A(n_4949),
.Y(n_5199)
);

AND2x2_ASAP7_75t_L g5200 ( 
.A(n_4874),
.B(n_4579),
.Y(n_5200)
);

AND2x4_ASAP7_75t_L g5201 ( 
.A(n_4894),
.B(n_4871),
.Y(n_5201)
);

HB1xp67_ASAP7_75t_L g5202 ( 
.A(n_4989),
.Y(n_5202)
);

AOI22xp5_ASAP7_75t_L g5203 ( 
.A1(n_4959),
.A2(n_4706),
.B1(n_4744),
.B2(n_4731),
.Y(n_5203)
);

INVx2_ASAP7_75t_L g5204 ( 
.A(n_4925),
.Y(n_5204)
);

BUFx6f_ASAP7_75t_L g5205 ( 
.A(n_4876),
.Y(n_5205)
);

AND2x4_ASAP7_75t_L g5206 ( 
.A(n_4894),
.B(n_4836),
.Y(n_5206)
);

HB1xp67_ASAP7_75t_L g5207 ( 
.A(n_5053),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_4944),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_4944),
.Y(n_5209)
);

INVx2_ASAP7_75t_L g5210 ( 
.A(n_4988),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_4958),
.Y(n_5211)
);

INVx2_ASAP7_75t_L g5212 ( 
.A(n_4962),
.Y(n_5212)
);

INVx2_ASAP7_75t_L g5213 ( 
.A(n_4958),
.Y(n_5213)
);

BUFx6f_ASAP7_75t_L g5214 ( 
.A(n_4934),
.Y(n_5214)
);

INVx2_ASAP7_75t_L g5215 ( 
.A(n_5126),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_4966),
.Y(n_5216)
);

INVx1_ASAP7_75t_L g5217 ( 
.A(n_4977),
.Y(n_5217)
);

INVx2_ASAP7_75t_L g5218 ( 
.A(n_5126),
.Y(n_5218)
);

INVx2_ASAP7_75t_L g5219 ( 
.A(n_5043),
.Y(n_5219)
);

OAI21x1_ASAP7_75t_L g5220 ( 
.A1(n_5081),
.A2(n_4853),
.B(n_4865),
.Y(n_5220)
);

OR2x2_ASAP7_75t_L g5221 ( 
.A(n_4879),
.B(n_4579),
.Y(n_5221)
);

INVx2_ASAP7_75t_L g5222 ( 
.A(n_5073),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_4954),
.Y(n_5223)
);

INVx2_ASAP7_75t_L g5224 ( 
.A(n_5083),
.Y(n_5224)
);

INVx2_ASAP7_75t_SL g5225 ( 
.A(n_4994),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_4919),
.Y(n_5226)
);

INVx2_ASAP7_75t_SL g5227 ( 
.A(n_4880),
.Y(n_5227)
);

OAI21xp33_ASAP7_75t_SL g5228 ( 
.A1(n_5086),
.A2(n_5090),
.B(n_5089),
.Y(n_5228)
);

INVx2_ASAP7_75t_L g5229 ( 
.A(n_5124),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_4879),
.Y(n_5230)
);

INVx2_ASAP7_75t_L g5231 ( 
.A(n_5130),
.Y(n_5231)
);

INVx3_ASAP7_75t_L g5232 ( 
.A(n_4949),
.Y(n_5232)
);

INVx2_ASAP7_75t_L g5233 ( 
.A(n_5113),
.Y(n_5233)
);

INVx1_ASAP7_75t_L g5234 ( 
.A(n_4885),
.Y(n_5234)
);

NAND2x1p5_ASAP7_75t_L g5235 ( 
.A(n_4939),
.B(n_4594),
.Y(n_5235)
);

BUFx3_ASAP7_75t_L g5236 ( 
.A(n_4880),
.Y(n_5236)
);

BUFx2_ASAP7_75t_L g5237 ( 
.A(n_4947),
.Y(n_5237)
);

INVx2_ASAP7_75t_L g5238 ( 
.A(n_5114),
.Y(n_5238)
);

NAND2xp5_ASAP7_75t_L g5239 ( 
.A(n_4904),
.B(n_4591),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_4930),
.Y(n_5240)
);

AO21x2_ASAP7_75t_L g5241 ( 
.A1(n_5099),
.A2(n_4723),
.B(n_4728),
.Y(n_5241)
);

AND2x2_ASAP7_75t_L g5242 ( 
.A(n_4916),
.B(n_4579),
.Y(n_5242)
);

INVx2_ASAP7_75t_L g5243 ( 
.A(n_5116),
.Y(n_5243)
);

INVx2_ASAP7_75t_L g5244 ( 
.A(n_5104),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_5119),
.Y(n_5245)
);

NAND2x1p5_ASAP7_75t_L g5246 ( 
.A(n_4981),
.B(n_4836),
.Y(n_5246)
);

INVx2_ASAP7_75t_L g5247 ( 
.A(n_5122),
.Y(n_5247)
);

INVx2_ASAP7_75t_L g5248 ( 
.A(n_5093),
.Y(n_5248)
);

BUFx3_ASAP7_75t_L g5249 ( 
.A(n_4880),
.Y(n_5249)
);

OAI21x1_ASAP7_75t_L g5250 ( 
.A1(n_5097),
.A2(n_4701),
.B(n_4845),
.Y(n_5250)
);

NAND2xp5_ASAP7_75t_L g5251 ( 
.A(n_4996),
.B(n_4591),
.Y(n_5251)
);

NAND2xp5_ASAP7_75t_L g5252 ( 
.A(n_4996),
.B(n_5040),
.Y(n_5252)
);

AND2x4_ASAP7_75t_L g5253 ( 
.A(n_4915),
.B(n_4845),
.Y(n_5253)
);

HB1xp67_ASAP7_75t_L g5254 ( 
.A(n_4937),
.Y(n_5254)
);

HB1xp67_ASAP7_75t_L g5255 ( 
.A(n_4937),
.Y(n_5255)
);

OAI33xp33_ASAP7_75t_L g5256 ( 
.A1(n_5084),
.A2(n_148),
.A3(n_150),
.B1(n_146),
.B2(n_147),
.B3(n_149),
.Y(n_5256)
);

NAND2xp5_ASAP7_75t_L g5257 ( 
.A(n_4911),
.B(n_4591),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_5072),
.Y(n_5258)
);

INVx1_ASAP7_75t_L g5259 ( 
.A(n_5059),
.Y(n_5259)
);

BUFx10_ASAP7_75t_L g5260 ( 
.A(n_4934),
.Y(n_5260)
);

OAI21x1_ASAP7_75t_L g5261 ( 
.A1(n_5026),
.A2(n_4593),
.B(n_4627),
.Y(n_5261)
);

OAI21x1_ASAP7_75t_L g5262 ( 
.A1(n_5026),
.A2(n_4627),
.B(n_4624),
.Y(n_5262)
);

HB1xp67_ASAP7_75t_L g5263 ( 
.A(n_4900),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_4995),
.Y(n_5264)
);

AOI21x1_ASAP7_75t_L g5265 ( 
.A1(n_5084),
.A2(n_2258),
.B(n_2255),
.Y(n_5265)
);

INVx2_ASAP7_75t_L g5266 ( 
.A(n_5100),
.Y(n_5266)
);

INVx3_ASAP7_75t_L g5267 ( 
.A(n_4981),
.Y(n_5267)
);

HB1xp67_ASAP7_75t_L g5268 ( 
.A(n_4900),
.Y(n_5268)
);

BUFx2_ASAP7_75t_L g5269 ( 
.A(n_5101),
.Y(n_5269)
);

INVx2_ASAP7_75t_L g5270 ( 
.A(n_5121),
.Y(n_5270)
);

INVx2_ASAP7_75t_L g5271 ( 
.A(n_5132),
.Y(n_5271)
);

BUFx2_ASAP7_75t_L g5272 ( 
.A(n_5088),
.Y(n_5272)
);

INVx2_ASAP7_75t_SL g5273 ( 
.A(n_4929),
.Y(n_5273)
);

INVx3_ASAP7_75t_L g5274 ( 
.A(n_5011),
.Y(n_5274)
);

OR2x6_ASAP7_75t_L g5275 ( 
.A(n_4961),
.B(n_4698),
.Y(n_5275)
);

AND2x4_ASAP7_75t_L g5276 ( 
.A(n_4905),
.B(n_4698),
.Y(n_5276)
);

NAND3x1_ASAP7_75t_L g5277 ( 
.A(n_4896),
.B(n_147),
.C(n_148),
.Y(n_5277)
);

BUFx2_ASAP7_75t_L g5278 ( 
.A(n_4902),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5038),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_5041),
.Y(n_5280)
);

OAI22xp5_ASAP7_75t_L g5281 ( 
.A1(n_5000),
.A2(n_2269),
.B1(n_2271),
.B2(n_2255),
.Y(n_5281)
);

INVx2_ASAP7_75t_L g5282 ( 
.A(n_4927),
.Y(n_5282)
);

INVx2_ASAP7_75t_L g5283 ( 
.A(n_4927),
.Y(n_5283)
);

INVx2_ASAP7_75t_L g5284 ( 
.A(n_5017),
.Y(n_5284)
);

INVx2_ASAP7_75t_L g5285 ( 
.A(n_5017),
.Y(n_5285)
);

A2O1A1Ixp33_ASAP7_75t_L g5286 ( 
.A1(n_5027),
.A2(n_153),
.B(n_150),
.C(n_152),
.Y(n_5286)
);

INVx2_ASAP7_75t_L g5287 ( 
.A(n_5019),
.Y(n_5287)
);

INVx2_ASAP7_75t_L g5288 ( 
.A(n_5019),
.Y(n_5288)
);

INVx2_ASAP7_75t_L g5289 ( 
.A(n_5057),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_5011),
.Y(n_5290)
);

INVx3_ASAP7_75t_L g5291 ( 
.A(n_4929),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_5014),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_5014),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_5031),
.Y(n_5294)
);

AOI22xp33_ASAP7_75t_L g5295 ( 
.A1(n_5079),
.A2(n_157),
.B1(n_152),
.B2(n_154),
.Y(n_5295)
);

AOI21x1_ASAP7_75t_L g5296 ( 
.A1(n_5085),
.A2(n_2282),
.B(n_2281),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_5064),
.Y(n_5297)
);

NAND2xp5_ASAP7_75t_L g5298 ( 
.A(n_4917),
.B(n_4889),
.Y(n_5298)
);

OR2x2_ASAP7_75t_L g5299 ( 
.A(n_5010),
.B(n_158),
.Y(n_5299)
);

NAND2xp5_ASAP7_75t_L g5300 ( 
.A(n_4917),
.B(n_159),
.Y(n_5300)
);

NAND2x1p5_ASAP7_75t_L g5301 ( 
.A(n_4987),
.B(n_4993),
.Y(n_5301)
);

INVx3_ASAP7_75t_L g5302 ( 
.A(n_4934),
.Y(n_5302)
);

INVx1_ASAP7_75t_L g5303 ( 
.A(n_5064),
.Y(n_5303)
);

OAI21x1_ASAP7_75t_L g5304 ( 
.A1(n_5057),
.A2(n_2282),
.B(n_2281),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_5115),
.Y(n_5305)
);

INVx3_ASAP7_75t_L g5306 ( 
.A(n_5037),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_5115),
.Y(n_5307)
);

BUFx3_ASAP7_75t_L g5308 ( 
.A(n_5036),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_5007),
.Y(n_5309)
);

INVx2_ASAP7_75t_L g5310 ( 
.A(n_5110),
.Y(n_5310)
);

AND2x2_ASAP7_75t_L g5311 ( 
.A(n_4951),
.B(n_161),
.Y(n_5311)
);

INVx1_ASAP7_75t_L g5312 ( 
.A(n_5007),
.Y(n_5312)
);

AND2x2_ASAP7_75t_L g5313 ( 
.A(n_4983),
.B(n_163),
.Y(n_5313)
);

OAI21x1_ASAP7_75t_L g5314 ( 
.A1(n_5058),
.A2(n_2302),
.B(n_2283),
.Y(n_5314)
);

INVx2_ASAP7_75t_SL g5315 ( 
.A(n_5095),
.Y(n_5315)
);

BUFx8_ASAP7_75t_SL g5316 ( 
.A(n_4940),
.Y(n_5316)
);

HB1xp67_ASAP7_75t_L g5317 ( 
.A(n_5018),
.Y(n_5317)
);

OR2x2_ASAP7_75t_L g5318 ( 
.A(n_4893),
.B(n_164),
.Y(n_5318)
);

HB1xp67_ASAP7_75t_L g5319 ( 
.A(n_5018),
.Y(n_5319)
);

INVx2_ASAP7_75t_L g5320 ( 
.A(n_5058),
.Y(n_5320)
);

OR2x2_ASAP7_75t_L g5321 ( 
.A(n_4888),
.B(n_165),
.Y(n_5321)
);

INVx2_ASAP7_75t_L g5322 ( 
.A(n_5118),
.Y(n_5322)
);

INVx2_ASAP7_75t_L g5323 ( 
.A(n_5105),
.Y(n_5323)
);

INVx1_ASAP7_75t_L g5324 ( 
.A(n_4922),
.Y(n_5324)
);

BUFx2_ASAP7_75t_L g5325 ( 
.A(n_4920),
.Y(n_5325)
);

BUFx3_ASAP7_75t_L g5326 ( 
.A(n_5008),
.Y(n_5326)
);

NAND2x1p5_ASAP7_75t_L g5327 ( 
.A(n_4978),
.B(n_1714),
.Y(n_5327)
);

INVx1_ASAP7_75t_SL g5328 ( 
.A(n_4882),
.Y(n_5328)
);

NOR2x1_ASAP7_75t_SL g5329 ( 
.A(n_5129),
.B(n_5085),
.Y(n_5329)
);

INVx2_ASAP7_75t_L g5330 ( 
.A(n_5129),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_4922),
.Y(n_5331)
);

HB1xp67_ASAP7_75t_L g5332 ( 
.A(n_5129),
.Y(n_5332)
);

INVx2_ASAP7_75t_L g5333 ( 
.A(n_5095),
.Y(n_5333)
);

INVx1_ASAP7_75t_L g5334 ( 
.A(n_5051),
.Y(n_5334)
);

BUFx6f_ASAP7_75t_L g5335 ( 
.A(n_5034),
.Y(n_5335)
);

INVx3_ASAP7_75t_L g5336 ( 
.A(n_4920),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_4906),
.Y(n_5337)
);

AND2x2_ASAP7_75t_L g5338 ( 
.A(n_4877),
.B(n_167),
.Y(n_5338)
);

AOI22xp33_ASAP7_75t_L g5339 ( 
.A1(n_5111),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_5339)
);

AND2x4_ASAP7_75t_L g5340 ( 
.A(n_4970),
.B(n_4920),
.Y(n_5340)
);

INVx1_ASAP7_75t_L g5341 ( 
.A(n_5049),
.Y(n_5341)
);

INVx5_ASAP7_75t_L g5342 ( 
.A(n_5030),
.Y(n_5342)
);

HB1xp67_ASAP7_75t_L g5343 ( 
.A(n_5086),
.Y(n_5343)
);

INVx2_ASAP7_75t_L g5344 ( 
.A(n_5070),
.Y(n_5344)
);

INVx3_ASAP7_75t_L g5345 ( 
.A(n_5045),
.Y(n_5345)
);

INVx2_ASAP7_75t_L g5346 ( 
.A(n_5075),
.Y(n_5346)
);

AOI22xp33_ASAP7_75t_L g5347 ( 
.A1(n_5343),
.A2(n_5009),
.B1(n_5094),
.B2(n_5090),
.Y(n_5347)
);

INVx2_ASAP7_75t_L g5348 ( 
.A(n_5171),
.Y(n_5348)
);

OAI22xp5_ASAP7_75t_L g5349 ( 
.A1(n_5145),
.A2(n_5094),
.B1(n_4909),
.B2(n_5022),
.Y(n_5349)
);

OAI21xp5_ASAP7_75t_L g5350 ( 
.A1(n_5228),
.A2(n_5103),
.B(n_5112),
.Y(n_5350)
);

NAND2xp5_ASAP7_75t_L g5351 ( 
.A(n_5178),
.B(n_5047),
.Y(n_5351)
);

OAI22xp5_ASAP7_75t_L g5352 ( 
.A1(n_5175),
.A2(n_5339),
.B1(n_5295),
.B2(n_5300),
.Y(n_5352)
);

OAI22xp5_ASAP7_75t_L g5353 ( 
.A1(n_5339),
.A2(n_4909),
.B1(n_4924),
.B2(n_4913),
.Y(n_5353)
);

AO221x1_ASAP7_75t_L g5354 ( 
.A1(n_5297),
.A2(n_4953),
.B1(n_4897),
.B2(n_4936),
.C(n_5061),
.Y(n_5354)
);

AOI22xp5_ASAP7_75t_L g5355 ( 
.A1(n_5324),
.A2(n_4936),
.B1(n_5123),
.B2(n_4897),
.Y(n_5355)
);

OAI211xp5_ASAP7_75t_L g5356 ( 
.A1(n_5295),
.A2(n_5331),
.B(n_5298),
.C(n_5255),
.Y(n_5356)
);

CKINVDCx8_ASAP7_75t_R g5357 ( 
.A(n_5135),
.Y(n_5357)
);

AOI22xp33_ASAP7_75t_SL g5358 ( 
.A1(n_5329),
.A2(n_5120),
.B1(n_5077),
.B2(n_5108),
.Y(n_5358)
);

CKINVDCx5p33_ASAP7_75t_R g5359 ( 
.A(n_5316),
.Y(n_5359)
);

CKINVDCx5p33_ASAP7_75t_R g5360 ( 
.A(n_5316),
.Y(n_5360)
);

AOI22xp33_ASAP7_75t_L g5361 ( 
.A1(n_5256),
.A2(n_4941),
.B1(n_5098),
.B2(n_5056),
.Y(n_5361)
);

O2A1O1Ixp33_ASAP7_75t_L g5362 ( 
.A1(n_5286),
.A2(n_5077),
.B(n_5066),
.C(n_5071),
.Y(n_5362)
);

AOI22xp5_ASAP7_75t_L g5363 ( 
.A1(n_5277),
.A2(n_5123),
.B1(n_5106),
.B2(n_4938),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_5202),
.Y(n_5364)
);

AND2x2_ASAP7_75t_L g5365 ( 
.A(n_5163),
.B(n_4956),
.Y(n_5365)
);

BUFx5_ASAP7_75t_L g5366 ( 
.A(n_5260),
.Y(n_5366)
);

AOI22xp33_ASAP7_75t_L g5367 ( 
.A1(n_5259),
.A2(n_5055),
.B1(n_4984),
.B2(n_5024),
.Y(n_5367)
);

AOI22xp33_ASAP7_75t_L g5368 ( 
.A1(n_5137),
.A2(n_5055),
.B1(n_5024),
.B2(n_5067),
.Y(n_5368)
);

OA21x2_ASAP7_75t_L g5369 ( 
.A1(n_5215),
.A2(n_4945),
.B(n_4878),
.Y(n_5369)
);

AOI21x1_ASAP7_75t_L g5370 ( 
.A1(n_5278),
.A2(n_5076),
.B(n_5066),
.Y(n_5370)
);

AOI21xp33_ASAP7_75t_L g5371 ( 
.A1(n_5257),
.A2(n_5071),
.B(n_5061),
.Y(n_5371)
);

AOI22xp33_ASAP7_75t_L g5372 ( 
.A1(n_5281),
.A2(n_5067),
.B1(n_5044),
.B2(n_5065),
.Y(n_5372)
);

INVx2_ASAP7_75t_L g5373 ( 
.A(n_5138),
.Y(n_5373)
);

OAI22xp33_ASAP7_75t_L g5374 ( 
.A1(n_5139),
.A2(n_4933),
.B1(n_4883),
.B2(n_4990),
.Y(n_5374)
);

AOI211xp5_ASAP7_75t_L g5375 ( 
.A1(n_5193),
.A2(n_5054),
.B(n_4991),
.C(n_5042),
.Y(n_5375)
);

AOI221xp5_ASAP7_75t_L g5376 ( 
.A1(n_5254),
.A2(n_5134),
.B1(n_5078),
.B2(n_4979),
.C(n_5102),
.Y(n_5376)
);

OAI22xp33_ASAP7_75t_L g5377 ( 
.A1(n_5303),
.A2(n_4938),
.B1(n_4932),
.B2(n_4969),
.Y(n_5377)
);

AND2x2_ASAP7_75t_L g5378 ( 
.A(n_5201),
.B(n_5237),
.Y(n_5378)
);

OAI211xp5_ASAP7_75t_L g5379 ( 
.A1(n_5254),
.A2(n_4903),
.B(n_4968),
.C(n_4892),
.Y(n_5379)
);

AOI21xp5_ASAP7_75t_L g5380 ( 
.A1(n_5189),
.A2(n_4972),
.B(n_4931),
.Y(n_5380)
);

INVx2_ASAP7_75t_L g5381 ( 
.A(n_5138),
.Y(n_5381)
);

OR2x6_ASAP7_75t_L g5382 ( 
.A(n_5235),
.B(n_4932),
.Y(n_5382)
);

AND2x4_ASAP7_75t_L g5383 ( 
.A(n_5201),
.B(n_5074),
.Y(n_5383)
);

AO21x2_ASAP7_75t_L g5384 ( 
.A1(n_5263),
.A2(n_5046),
.B(n_5082),
.Y(n_5384)
);

INVx2_ASAP7_75t_L g5385 ( 
.A(n_5140),
.Y(n_5385)
);

OAI21xp5_ASAP7_75t_L g5386 ( 
.A1(n_5277),
.A2(n_4935),
.B(n_4914),
.Y(n_5386)
);

AOI22xp33_ASAP7_75t_L g5387 ( 
.A1(n_5258),
.A2(n_4985),
.B1(n_4946),
.B2(n_5092),
.Y(n_5387)
);

OAI22xp5_ASAP7_75t_L g5388 ( 
.A1(n_5318),
.A2(n_4887),
.B1(n_4901),
.B2(n_4976),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_5207),
.Y(n_5389)
);

AOI22xp33_ASAP7_75t_L g5390 ( 
.A1(n_5279),
.A2(n_5063),
.B1(n_4870),
.B2(n_4928),
.Y(n_5390)
);

OAI22xp5_ASAP7_75t_L g5391 ( 
.A1(n_5321),
.A2(n_4975),
.B1(n_5074),
.B2(n_5003),
.Y(n_5391)
);

AOI22xp33_ASAP7_75t_L g5392 ( 
.A1(n_5280),
.A2(n_5107),
.B1(n_5002),
.B2(n_5117),
.Y(n_5392)
);

OAI33xp33_ASAP7_75t_L g5393 ( 
.A1(n_5251),
.A2(n_5060),
.A3(n_5050),
.B1(n_5091),
.B2(n_173),
.B3(n_175),
.Y(n_5393)
);

OA211x2_ASAP7_75t_L g5394 ( 
.A1(n_5239),
.A2(n_5033),
.B(n_5016),
.C(n_5005),
.Y(n_5394)
);

OAI221xp5_ASAP7_75t_L g5395 ( 
.A1(n_5210),
.A2(n_5048),
.B1(n_5004),
.B2(n_5006),
.C(n_5020),
.Y(n_5395)
);

OAI221xp5_ASAP7_75t_L g5396 ( 
.A1(n_5210),
.A2(n_5068),
.B1(n_5001),
.B2(n_5023),
.C(n_5062),
.Y(n_5396)
);

OAI221xp5_ASAP7_75t_L g5397 ( 
.A1(n_5264),
.A2(n_5087),
.B1(n_5080),
.B2(n_5128),
.C(n_5109),
.Y(n_5397)
);

INVx4_ASAP7_75t_L g5398 ( 
.A(n_5156),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_5148),
.Y(n_5399)
);

INVx2_ASAP7_75t_L g5400 ( 
.A(n_5140),
.Y(n_5400)
);

AOI321xp33_ASAP7_75t_L g5401 ( 
.A1(n_5341),
.A2(n_173),
.A3(n_176),
.B1(n_169),
.B2(n_172),
.C(n_174),
.Y(n_5401)
);

AOI22xp33_ASAP7_75t_L g5402 ( 
.A1(n_5231),
.A2(n_5030),
.B1(n_5016),
.B2(n_5045),
.Y(n_5402)
);

AOI22xp33_ASAP7_75t_L g5403 ( 
.A1(n_5337),
.A2(n_5029),
.B1(n_5133),
.B2(n_2186),
.Y(n_5403)
);

OAI221xp5_ASAP7_75t_L g5404 ( 
.A1(n_5305),
.A2(n_5307),
.B1(n_5334),
.B2(n_5252),
.C(n_5294),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5153),
.Y(n_5405)
);

AOI22xp33_ASAP7_75t_L g5406 ( 
.A1(n_5274),
.A2(n_5029),
.B1(n_2186),
.B2(n_1899),
.Y(n_5406)
);

OAI221xp5_ASAP7_75t_L g5407 ( 
.A1(n_5240),
.A2(n_180),
.B1(n_177),
.B2(n_179),
.C(n_182),
.Y(n_5407)
);

OR2x2_ASAP7_75t_L g5408 ( 
.A(n_5204),
.B(n_179),
.Y(n_5408)
);

AOI22xp33_ASAP7_75t_L g5409 ( 
.A1(n_5274),
.A2(n_1899),
.B1(n_1880),
.B2(n_2179),
.Y(n_5409)
);

OAI21xp5_ASAP7_75t_SL g5410 ( 
.A1(n_5338),
.A2(n_5205),
.B(n_5156),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_5160),
.Y(n_5411)
);

AOI22xp33_ASAP7_75t_L g5412 ( 
.A1(n_5274),
.A2(n_1899),
.B1(n_1880),
.B2(n_2179),
.Y(n_5412)
);

AND2x4_ASAP7_75t_L g5413 ( 
.A(n_5340),
.B(n_183),
.Y(n_5413)
);

OR2x2_ASAP7_75t_L g5414 ( 
.A(n_5204),
.B(n_186),
.Y(n_5414)
);

INVx2_ASAP7_75t_L g5415 ( 
.A(n_5213),
.Y(n_5415)
);

AOI221xp5_ASAP7_75t_L g5416 ( 
.A1(n_5268),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.C(n_192),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_5213),
.Y(n_5417)
);

AOI221xp5_ASAP7_75t_L g5418 ( 
.A1(n_5268),
.A2(n_5162),
.B1(n_5158),
.B2(n_5209),
.C(n_5208),
.Y(n_5418)
);

AOI221xp5_ASAP7_75t_SL g5419 ( 
.A1(n_5142),
.A2(n_194),
.B1(n_197),
.B2(n_190),
.C(n_196),
.Y(n_5419)
);

AOI22xp33_ASAP7_75t_L g5420 ( 
.A1(n_5344),
.A2(n_1899),
.B1(n_1880),
.B2(n_2179),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_5164),
.Y(n_5421)
);

AOI22xp33_ASAP7_75t_L g5422 ( 
.A1(n_5344),
.A2(n_5346),
.B1(n_5290),
.B2(n_5293),
.Y(n_5422)
);

NAND2xp5_ASAP7_75t_L g5423 ( 
.A(n_5216),
.B(n_198),
.Y(n_5423)
);

OAI21xp5_ASAP7_75t_L g5424 ( 
.A1(n_5187),
.A2(n_5296),
.B(n_5265),
.Y(n_5424)
);

AOI22xp33_ASAP7_75t_L g5425 ( 
.A1(n_5346),
.A2(n_1899),
.B1(n_1880),
.B2(n_1615),
.Y(n_5425)
);

AOI22xp33_ASAP7_75t_L g5426 ( 
.A1(n_5292),
.A2(n_1880),
.B1(n_1631),
.B2(n_1644),
.Y(n_5426)
);

AOI221xp5_ASAP7_75t_L g5427 ( 
.A1(n_5158),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.C(n_202),
.Y(n_5427)
);

OR2x2_ASAP7_75t_L g5428 ( 
.A(n_5180),
.B(n_200),
.Y(n_5428)
);

INVx1_ASAP7_75t_L g5429 ( 
.A(n_5165),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_5167),
.Y(n_5430)
);

AOI221xp5_ASAP7_75t_L g5431 ( 
.A1(n_5162),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.C(n_206),
.Y(n_5431)
);

OAI22xp5_ASAP7_75t_L g5432 ( 
.A1(n_5203),
.A2(n_208),
.B1(n_203),
.B2(n_207),
.Y(n_5432)
);

AOI22xp33_ASAP7_75t_SL g5433 ( 
.A1(n_5156),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_5433)
);

INVx4_ASAP7_75t_L g5434 ( 
.A(n_5156),
.Y(n_5434)
);

OAI221xp5_ASAP7_75t_L g5435 ( 
.A1(n_5273),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.C(n_212),
.Y(n_5435)
);

AOI221xp5_ASAP7_75t_L g5436 ( 
.A1(n_5200),
.A2(n_215),
.B1(n_210),
.B2(n_213),
.C(n_216),
.Y(n_5436)
);

AOI22xp33_ASAP7_75t_L g5437 ( 
.A1(n_5242),
.A2(n_1644),
.B1(n_1651),
.B2(n_1587),
.Y(n_5437)
);

INVx2_ASAP7_75t_L g5438 ( 
.A(n_5146),
.Y(n_5438)
);

BUFx2_ASAP7_75t_L g5439 ( 
.A(n_5272),
.Y(n_5439)
);

INVx2_ASAP7_75t_L g5440 ( 
.A(n_5146),
.Y(n_5440)
);

BUFx6f_ASAP7_75t_L g5441 ( 
.A(n_5205),
.Y(n_5441)
);

OAI211xp5_ASAP7_75t_L g5442 ( 
.A1(n_5185),
.A2(n_223),
.B(n_219),
.C(n_220),
.Y(n_5442)
);

AOI22xp5_ASAP7_75t_L g5443 ( 
.A1(n_5284),
.A2(n_1663),
.B1(n_1686),
.B2(n_1657),
.Y(n_5443)
);

AOI21xp5_ASAP7_75t_L g5444 ( 
.A1(n_5275),
.A2(n_1663),
.B(n_1657),
.Y(n_5444)
);

INVx1_ASAP7_75t_L g5445 ( 
.A(n_5169),
.Y(n_5445)
);

OAI221xp5_ASAP7_75t_L g5446 ( 
.A1(n_5273),
.A2(n_229),
.B1(n_226),
.B2(n_228),
.C(n_230),
.Y(n_5446)
);

AND2x4_ASAP7_75t_L g5447 ( 
.A(n_5336),
.B(n_229),
.Y(n_5447)
);

CKINVDCx20_ASAP7_75t_R g5448 ( 
.A(n_5196),
.Y(n_5448)
);

OAI22xp5_ASAP7_75t_SL g5449 ( 
.A1(n_5326),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_5449)
);

AOI22xp33_ASAP7_75t_L g5450 ( 
.A1(n_5285),
.A2(n_5287),
.B1(n_5288),
.B2(n_5226),
.Y(n_5450)
);

INVx1_ASAP7_75t_L g5451 ( 
.A(n_5170),
.Y(n_5451)
);

AOI22xp5_ASAP7_75t_L g5452 ( 
.A1(n_5285),
.A2(n_1686),
.B1(n_1712),
.B2(n_1691),
.Y(n_5452)
);

O2A1O1Ixp33_ASAP7_75t_SL g5453 ( 
.A1(n_5191),
.A2(n_234),
.B(n_232),
.C(n_233),
.Y(n_5453)
);

NOR2x1_ASAP7_75t_R g5454 ( 
.A(n_5326),
.B(n_233),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_5177),
.Y(n_5455)
);

OAI221xp5_ASAP7_75t_L g5456 ( 
.A1(n_5151),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.C(n_237),
.Y(n_5456)
);

NAND3xp33_ASAP7_75t_L g5457 ( 
.A(n_5282),
.B(n_235),
.C(n_236),
.Y(n_5457)
);

AOI221xp5_ASAP7_75t_L g5458 ( 
.A1(n_5230),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.C(n_241),
.Y(n_5458)
);

OAI221xp5_ASAP7_75t_L g5459 ( 
.A1(n_5221),
.A2(n_242),
.B1(n_239),
.B2(n_241),
.C(n_244),
.Y(n_5459)
);

INVx2_ASAP7_75t_SL g5460 ( 
.A(n_5184),
.Y(n_5460)
);

AO21x2_ASAP7_75t_L g5461 ( 
.A1(n_5282),
.A2(n_245),
.B(n_248),
.Y(n_5461)
);

OAI22xp5_ASAP7_75t_L g5462 ( 
.A1(n_5327),
.A2(n_256),
.B1(n_253),
.B2(n_255),
.Y(n_5462)
);

NAND2xp5_ASAP7_75t_L g5463 ( 
.A(n_5217),
.B(n_255),
.Y(n_5463)
);

AOI22xp33_ASAP7_75t_L g5464 ( 
.A1(n_5223),
.A2(n_1744),
.B1(n_1756),
.B2(n_1740),
.Y(n_5464)
);

AOI211xp5_ASAP7_75t_L g5465 ( 
.A1(n_5299),
.A2(n_258),
.B(n_256),
.C(n_257),
.Y(n_5465)
);

AND2x2_ASAP7_75t_L g5466 ( 
.A(n_5325),
.B(n_257),
.Y(n_5466)
);

OAI221xp5_ASAP7_75t_SL g5467 ( 
.A1(n_5283),
.A2(n_5190),
.B1(n_5212),
.B2(n_5152),
.C(n_5147),
.Y(n_5467)
);

AND2x2_ASAP7_75t_L g5468 ( 
.A(n_5173),
.B(n_259),
.Y(n_5468)
);

AND2x2_ASAP7_75t_L g5469 ( 
.A(n_5173),
.B(n_260),
.Y(n_5469)
);

OAI221xp5_ASAP7_75t_L g5470 ( 
.A1(n_5191),
.A2(n_267),
.B1(n_262),
.B2(n_264),
.C(n_268),
.Y(n_5470)
);

A2O1A1Ixp33_ASAP7_75t_L g5471 ( 
.A1(n_5199),
.A2(n_271),
.B(n_268),
.C(n_269),
.Y(n_5471)
);

AND2x2_ASAP7_75t_L g5472 ( 
.A(n_5269),
.B(n_269),
.Y(n_5472)
);

OR2x6_ASAP7_75t_L g5473 ( 
.A(n_5199),
.B(n_272),
.Y(n_5473)
);

OAI22xp33_ASAP7_75t_L g5474 ( 
.A1(n_5342),
.A2(n_5199),
.B1(n_5225),
.B2(n_5232),
.Y(n_5474)
);

AOI221xp5_ASAP7_75t_L g5475 ( 
.A1(n_5234),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.C(n_277),
.Y(n_5475)
);

OAI332xp33_ASAP7_75t_L g5476 ( 
.A1(n_5283),
.A2(n_283),
.A3(n_282),
.B1(n_279),
.B2(n_285),
.B3(n_273),
.C1(n_274),
.C2(n_281),
.Y(n_5476)
);

OAI221xp5_ASAP7_75t_L g5477 ( 
.A1(n_5192),
.A2(n_289),
.B1(n_286),
.B2(n_287),
.C(n_290),
.Y(n_5477)
);

OAI22xp5_ASAP7_75t_L g5478 ( 
.A1(n_5205),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_5478)
);

AOI22xp33_ASAP7_75t_L g5479 ( 
.A1(n_5205),
.A2(n_1716),
.B1(n_1727),
.B2(n_1720),
.Y(n_5479)
);

AOI221xp5_ASAP7_75t_SL g5480 ( 
.A1(n_5245),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.C(n_297),
.Y(n_5480)
);

OAI22xp5_ASAP7_75t_L g5481 ( 
.A1(n_5342),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_5481)
);

OAI221xp5_ASAP7_75t_L g5482 ( 
.A1(n_5301),
.A2(n_5328),
.B1(n_5291),
.B2(n_5312),
.C(n_5309),
.Y(n_5482)
);

OAI21x1_ASAP7_75t_L g5483 ( 
.A1(n_5261),
.A2(n_1750),
.B(n_1714),
.Y(n_5483)
);

INVx4_ASAP7_75t_L g5484 ( 
.A(n_5214),
.Y(n_5484)
);

OAI22xp5_ASAP7_75t_L g5485 ( 
.A1(n_5301),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_5485)
);

OAI22xp33_ASAP7_75t_L g5486 ( 
.A1(n_5232),
.A2(n_5336),
.B1(n_5291),
.B2(n_5214),
.Y(n_5486)
);

NOR2xp33_ASAP7_75t_L g5487 ( 
.A(n_5308),
.B(n_301),
.Y(n_5487)
);

INVx2_ASAP7_75t_L g5488 ( 
.A(n_5154),
.Y(n_5488)
);

AOI22xp33_ASAP7_75t_L g5489 ( 
.A1(n_5211),
.A2(n_1716),
.B1(n_1727),
.B2(n_1720),
.Y(n_5489)
);

OAI22xp5_ASAP7_75t_L g5490 ( 
.A1(n_5236),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.Y(n_5490)
);

AOI221xp5_ASAP7_75t_L g5491 ( 
.A1(n_5218),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.C(n_308),
.Y(n_5491)
);

NAND4xp25_ASAP7_75t_L g5492 ( 
.A(n_5311),
.B(n_310),
.C(n_308),
.D(n_309),
.Y(n_5492)
);

AOI221xp5_ASAP7_75t_L g5493 ( 
.A1(n_5218),
.A2(n_315),
.B1(n_311),
.B2(n_314),
.C(n_316),
.Y(n_5493)
);

OAI22xp5_ASAP7_75t_L g5494 ( 
.A1(n_5249),
.A2(n_317),
.B1(n_311),
.B2(n_316),
.Y(n_5494)
);

OAI22xp33_ASAP7_75t_L g5495 ( 
.A1(n_5214),
.A2(n_321),
.B1(n_318),
.B2(n_319),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5155),
.Y(n_5496)
);

AOI22xp33_ASAP7_75t_L g5497 ( 
.A1(n_5330),
.A2(n_1727),
.B1(n_1735),
.B2(n_1720),
.Y(n_5497)
);

OAI211xp5_ASAP7_75t_L g5498 ( 
.A1(n_5317),
.A2(n_324),
.B(n_319),
.C(n_322),
.Y(n_5498)
);

INVx2_ASAP7_75t_L g5499 ( 
.A(n_5155),
.Y(n_5499)
);

AOI211xp5_ASAP7_75t_L g5500 ( 
.A1(n_5313),
.A2(n_5335),
.B(n_5332),
.C(n_5319),
.Y(n_5500)
);

NAND2xp5_ASAP7_75t_L g5501 ( 
.A(n_5182),
.B(n_322),
.Y(n_5501)
);

OAI21xp5_ASAP7_75t_L g5502 ( 
.A1(n_5149),
.A2(n_325),
.B(n_326),
.Y(n_5502)
);

OAI221xp5_ASAP7_75t_L g5503 ( 
.A1(n_5227),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.C(n_335),
.Y(n_5503)
);

BUFx2_ASAP7_75t_L g5504 ( 
.A(n_5439),
.Y(n_5504)
);

NAND2xp5_ASAP7_75t_L g5505 ( 
.A(n_5455),
.B(n_5179),
.Y(n_5505)
);

AND2x2_ASAP7_75t_L g5506 ( 
.A(n_5378),
.B(n_5333),
.Y(n_5506)
);

AND2x2_ASAP7_75t_L g5507 ( 
.A(n_5365),
.B(n_5267),
.Y(n_5507)
);

INVxp67_ASAP7_75t_L g5508 ( 
.A(n_5454),
.Y(n_5508)
);

INVx2_ASAP7_75t_L g5509 ( 
.A(n_5441),
.Y(n_5509)
);

AND2x2_ASAP7_75t_L g5510 ( 
.A(n_5383),
.B(n_5315),
.Y(n_5510)
);

AOI22xp33_ASAP7_75t_SL g5511 ( 
.A1(n_5354),
.A2(n_5352),
.B1(n_5349),
.B2(n_5350),
.Y(n_5511)
);

OAI222xp33_ASAP7_75t_L g5512 ( 
.A1(n_5358),
.A2(n_5315),
.B1(n_5302),
.B2(n_5159),
.C1(n_5197),
.C2(n_5174),
.Y(n_5512)
);

INVx2_ASAP7_75t_L g5513 ( 
.A(n_5441),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_5399),
.Y(n_5514)
);

INVx2_ASAP7_75t_L g5515 ( 
.A(n_5484),
.Y(n_5515)
);

BUFx6f_ASAP7_75t_L g5516 ( 
.A(n_5473),
.Y(n_5516)
);

INVx1_ASAP7_75t_L g5517 ( 
.A(n_5405),
.Y(n_5517)
);

INVx3_ASAP7_75t_L g5518 ( 
.A(n_5398),
.Y(n_5518)
);

INVx2_ASAP7_75t_L g5519 ( 
.A(n_5415),
.Y(n_5519)
);

INVx2_ASAP7_75t_L g5520 ( 
.A(n_5417),
.Y(n_5520)
);

AO22x1_ASAP7_75t_L g5521 ( 
.A1(n_5350),
.A2(n_5150),
.B1(n_5136),
.B2(n_5144),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_5411),
.Y(n_5522)
);

INVx2_ASAP7_75t_L g5523 ( 
.A(n_5348),
.Y(n_5523)
);

NAND2xp5_ASAP7_75t_L g5524 ( 
.A(n_5418),
.B(n_5188),
.Y(n_5524)
);

INVx1_ASAP7_75t_L g5525 ( 
.A(n_5421),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_5429),
.Y(n_5526)
);

INVx2_ASAP7_75t_L g5527 ( 
.A(n_5373),
.Y(n_5527)
);

INVx2_ASAP7_75t_L g5528 ( 
.A(n_5381),
.Y(n_5528)
);

INVx2_ASAP7_75t_L g5529 ( 
.A(n_5385),
.Y(n_5529)
);

INVx3_ASAP7_75t_L g5530 ( 
.A(n_5434),
.Y(n_5530)
);

NAND2xp5_ASAP7_75t_L g5531 ( 
.A(n_5430),
.B(n_5157),
.Y(n_5531)
);

NAND2xp5_ASAP7_75t_L g5532 ( 
.A(n_5445),
.B(n_5157),
.Y(n_5532)
);

HB1xp67_ASAP7_75t_L g5533 ( 
.A(n_5364),
.Y(n_5533)
);

AOI33xp33_ASAP7_75t_L g5534 ( 
.A1(n_5347),
.A2(n_5198),
.A3(n_5194),
.B1(n_5247),
.B2(n_5181),
.B3(n_5186),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_5451),
.Y(n_5535)
);

NAND2xp5_ASAP7_75t_L g5536 ( 
.A(n_5389),
.B(n_5161),
.Y(n_5536)
);

INVx2_ASAP7_75t_L g5537 ( 
.A(n_5400),
.Y(n_5537)
);

NOR2xp33_ASAP7_75t_R g5538 ( 
.A(n_5448),
.B(n_5260),
.Y(n_5538)
);

INVx1_ASAP7_75t_L g5539 ( 
.A(n_5496),
.Y(n_5539)
);

NAND2xp5_ASAP7_75t_L g5540 ( 
.A(n_5371),
.B(n_5161),
.Y(n_5540)
);

INVxp67_ASAP7_75t_SL g5541 ( 
.A(n_5500),
.Y(n_5541)
);

BUFx2_ASAP7_75t_L g5542 ( 
.A(n_5434),
.Y(n_5542)
);

AND2x2_ASAP7_75t_L g5543 ( 
.A(n_5500),
.B(n_5323),
.Y(n_5543)
);

INVx2_ASAP7_75t_L g5544 ( 
.A(n_5438),
.Y(n_5544)
);

OR2x2_ASAP7_75t_L g5545 ( 
.A(n_5408),
.B(n_5414),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_5440),
.Y(n_5546)
);

INVx2_ASAP7_75t_L g5547 ( 
.A(n_5413),
.Y(n_5547)
);

NOR2xp33_ASAP7_75t_L g5548 ( 
.A(n_5356),
.B(n_5150),
.Y(n_5548)
);

AND2x2_ASAP7_75t_L g5549 ( 
.A(n_5460),
.B(n_5176),
.Y(n_5549)
);

NAND2xp5_ASAP7_75t_L g5550 ( 
.A(n_5488),
.B(n_5143),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_5499),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5428),
.Y(n_5552)
);

CKINVDCx20_ASAP7_75t_R g5553 ( 
.A(n_5359),
.Y(n_5553)
);

AND2x2_ASAP7_75t_L g5554 ( 
.A(n_5450),
.B(n_5322),
.Y(n_5554)
);

AND2x2_ASAP7_75t_L g5555 ( 
.A(n_5422),
.B(n_5382),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_5461),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_5461),
.Y(n_5557)
);

INVx1_ASAP7_75t_L g5558 ( 
.A(n_5501),
.Y(n_5558)
);

AOI22xp33_ASAP7_75t_L g5559 ( 
.A1(n_5376),
.A2(n_5368),
.B1(n_5353),
.B2(n_5363),
.Y(n_5559)
);

NAND2xp5_ASAP7_75t_L g5560 ( 
.A(n_5423),
.B(n_5143),
.Y(n_5560)
);

INVx2_ASAP7_75t_L g5561 ( 
.A(n_5447),
.Y(n_5561)
);

INVx2_ASAP7_75t_L g5562 ( 
.A(n_5468),
.Y(n_5562)
);

AOI22xp33_ASAP7_75t_L g5563 ( 
.A1(n_5361),
.A2(n_5393),
.B1(n_5367),
.B2(n_5355),
.Y(n_5563)
);

NOR2x1_ASAP7_75t_L g5564 ( 
.A(n_5410),
.B(n_5306),
.Y(n_5564)
);

OR2x2_ASAP7_75t_L g5565 ( 
.A(n_5404),
.B(n_5369),
.Y(n_5565)
);

INVx1_ASAP7_75t_L g5566 ( 
.A(n_5469),
.Y(n_5566)
);

BUFx6f_ASAP7_75t_L g5567 ( 
.A(n_5473),
.Y(n_5567)
);

INVx2_ASAP7_75t_L g5568 ( 
.A(n_5370),
.Y(n_5568)
);

AOI211xp5_ASAP7_75t_L g5569 ( 
.A1(n_5380),
.A2(n_5206),
.B(n_5330),
.C(n_5253),
.Y(n_5569)
);

INVx2_ASAP7_75t_L g5570 ( 
.A(n_5366),
.Y(n_5570)
);

INVx3_ASAP7_75t_L g5571 ( 
.A(n_5357),
.Y(n_5571)
);

HB1xp67_ASAP7_75t_L g5572 ( 
.A(n_5384),
.Y(n_5572)
);

NAND2xp5_ASAP7_75t_L g5573 ( 
.A(n_5463),
.B(n_5229),
.Y(n_5573)
);

INVx2_ASAP7_75t_L g5574 ( 
.A(n_5366),
.Y(n_5574)
);

NAND2xp5_ASAP7_75t_L g5575 ( 
.A(n_5351),
.B(n_5233),
.Y(n_5575)
);

OAI22xp5_ASAP7_75t_L g5576 ( 
.A1(n_5375),
.A2(n_5320),
.B1(n_5246),
.B2(n_5345),
.Y(n_5576)
);

INVx1_ASAP7_75t_L g5577 ( 
.A(n_5472),
.Y(n_5577)
);

OA21x2_ASAP7_75t_L g5578 ( 
.A1(n_5480),
.A2(n_5238),
.B(n_5233),
.Y(n_5578)
);

AO21x2_ASAP7_75t_L g5579 ( 
.A1(n_5486),
.A2(n_5474),
.B(n_5457),
.Y(n_5579)
);

INVx3_ASAP7_75t_SL g5580 ( 
.A(n_5360),
.Y(n_5580)
);

NAND2xp5_ASAP7_75t_L g5581 ( 
.A(n_5377),
.B(n_5238),
.Y(n_5581)
);

INVx2_ASAP7_75t_L g5582 ( 
.A(n_5366),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_5379),
.Y(n_5583)
);

NAND2xp5_ASAP7_75t_L g5584 ( 
.A(n_5502),
.B(n_5243),
.Y(n_5584)
);

OR2x2_ASAP7_75t_L g5585 ( 
.A(n_5482),
.B(n_5266),
.Y(n_5585)
);

INVx2_ASAP7_75t_SL g5586 ( 
.A(n_5466),
.Y(n_5586)
);

INVx2_ASAP7_75t_L g5587 ( 
.A(n_5366),
.Y(n_5587)
);

OR2x2_ASAP7_75t_L g5588 ( 
.A(n_5467),
.B(n_5266),
.Y(n_5588)
);

AOI22xp33_ASAP7_75t_L g5589 ( 
.A1(n_5456),
.A2(n_5183),
.B1(n_5310),
.B2(n_5320),
.Y(n_5589)
);

AOI22xp33_ASAP7_75t_L g5590 ( 
.A1(n_5458),
.A2(n_5183),
.B1(n_5310),
.B2(n_5241),
.Y(n_5590)
);

AND2x4_ASAP7_75t_L g5591 ( 
.A(n_5386),
.B(n_5253),
.Y(n_5591)
);

AND2x2_ASAP7_75t_L g5592 ( 
.A(n_5390),
.B(n_5345),
.Y(n_5592)
);

AOI21xp33_ASAP7_75t_L g5593 ( 
.A1(n_5362),
.A2(n_5271),
.B(n_5270),
.Y(n_5593)
);

AND2x4_ASAP7_75t_L g5594 ( 
.A(n_5386),
.B(n_5276),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_5457),
.Y(n_5595)
);

INVx3_ASAP7_75t_L g5596 ( 
.A(n_5483),
.Y(n_5596)
);

INVxp67_ASAP7_75t_SL g5597 ( 
.A(n_5465),
.Y(n_5597)
);

AND2x2_ASAP7_75t_L g5598 ( 
.A(n_5387),
.B(n_5260),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_5394),
.Y(n_5599)
);

INVx2_ASAP7_75t_L g5600 ( 
.A(n_5443),
.Y(n_5600)
);

AND2x2_ASAP7_75t_L g5601 ( 
.A(n_5402),
.B(n_5276),
.Y(n_5601)
);

BUFx2_ASAP7_75t_L g5602 ( 
.A(n_5424),
.Y(n_5602)
);

AND2x2_ASAP7_75t_L g5603 ( 
.A(n_5391),
.B(n_5246),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_5452),
.Y(n_5604)
);

AOI22xp33_ASAP7_75t_L g5605 ( 
.A1(n_5475),
.A2(n_5416),
.B1(n_5372),
.B2(n_5427),
.Y(n_5605)
);

AND2x4_ASAP7_75t_L g5606 ( 
.A(n_5424),
.B(n_5244),
.Y(n_5606)
);

INVx1_ASAP7_75t_L g5607 ( 
.A(n_5388),
.Y(n_5607)
);

NAND2x1_ASAP7_75t_L g5608 ( 
.A(n_5481),
.B(n_5248),
.Y(n_5608)
);

INVx1_ASAP7_75t_L g5609 ( 
.A(n_5388),
.Y(n_5609)
);

INVx2_ASAP7_75t_L g5610 ( 
.A(n_5487),
.Y(n_5610)
);

INVx1_ASAP7_75t_L g5611 ( 
.A(n_5459),
.Y(n_5611)
);

INVx2_ASAP7_75t_L g5612 ( 
.A(n_5481),
.Y(n_5612)
);

AND2x2_ASAP7_75t_L g5613 ( 
.A(n_5437),
.B(n_5195),
.Y(n_5613)
);

INVx2_ASAP7_75t_L g5614 ( 
.A(n_5485),
.Y(n_5614)
);

AND2x2_ASAP7_75t_L g5615 ( 
.A(n_5375),
.B(n_5195),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_5442),
.Y(n_5616)
);

BUFx6f_ASAP7_75t_L g5617 ( 
.A(n_5476),
.Y(n_5617)
);

BUFx2_ASAP7_75t_L g5618 ( 
.A(n_5492),
.Y(n_5618)
);

INVx1_ASAP7_75t_L g5619 ( 
.A(n_5374),
.Y(n_5619)
);

INVx1_ASAP7_75t_L g5620 ( 
.A(n_5465),
.Y(n_5620)
);

INVx2_ASAP7_75t_L g5621 ( 
.A(n_5432),
.Y(n_5621)
);

INVx2_ASAP7_75t_L g5622 ( 
.A(n_5435),
.Y(n_5622)
);

NAND2xp5_ASAP7_75t_L g5623 ( 
.A(n_5436),
.B(n_5219),
.Y(n_5623)
);

INVx2_ASAP7_75t_L g5624 ( 
.A(n_5446),
.Y(n_5624)
);

HB1xp67_ASAP7_75t_L g5625 ( 
.A(n_5444),
.Y(n_5625)
);

INVxp67_ASAP7_75t_L g5626 ( 
.A(n_5449),
.Y(n_5626)
);

NAND2xp5_ASAP7_75t_L g5627 ( 
.A(n_5419),
.B(n_5222),
.Y(n_5627)
);

NAND2xp5_ASAP7_75t_L g5628 ( 
.A(n_5419),
.B(n_5222),
.Y(n_5628)
);

INVx3_ASAP7_75t_L g5629 ( 
.A(n_5476),
.Y(n_5629)
);

INVx2_ASAP7_75t_L g5630 ( 
.A(n_5407),
.Y(n_5630)
);

INVx2_ASAP7_75t_L g5631 ( 
.A(n_5470),
.Y(n_5631)
);

OR2x6_ASAP7_75t_L g5632 ( 
.A(n_5498),
.B(n_5172),
.Y(n_5632)
);

BUFx3_ASAP7_75t_L g5633 ( 
.A(n_5477),
.Y(n_5633)
);

INVx2_ASAP7_75t_L g5634 ( 
.A(n_5503),
.Y(n_5634)
);

AND2x2_ASAP7_75t_L g5635 ( 
.A(n_5392),
.B(n_5224),
.Y(n_5635)
);

INVx2_ASAP7_75t_L g5636 ( 
.A(n_5490),
.Y(n_5636)
);

AOI33xp33_ASAP7_75t_L g5637 ( 
.A1(n_5433),
.A2(n_5289),
.A3(n_338),
.B1(n_341),
.B2(n_335),
.B3(n_337),
.Y(n_5637)
);

OR2x2_ASAP7_75t_L g5638 ( 
.A(n_5420),
.B(n_5220),
.Y(n_5638)
);

AND2x2_ASAP7_75t_L g5639 ( 
.A(n_5497),
.B(n_5262),
.Y(n_5639)
);

INVx1_ASAP7_75t_L g5640 ( 
.A(n_5494),
.Y(n_5640)
);

OR2x2_ASAP7_75t_L g5641 ( 
.A(n_5425),
.B(n_5220),
.Y(n_5641)
);

AOI22xp33_ASAP7_75t_L g5642 ( 
.A1(n_5617),
.A2(n_5493),
.B1(n_5491),
.B2(n_5431),
.Y(n_5642)
);

OR2x6_ASAP7_75t_L g5643 ( 
.A(n_5516),
.B(n_5567),
.Y(n_5643)
);

AOI21xp5_ASAP7_75t_L g5644 ( 
.A1(n_5597),
.A2(n_5453),
.B(n_5471),
.Y(n_5644)
);

OAI211xp5_ASAP7_75t_SL g5645 ( 
.A1(n_5511),
.A2(n_5401),
.B(n_5495),
.C(n_5478),
.Y(n_5645)
);

NAND2xp5_ASAP7_75t_L g5646 ( 
.A(n_5595),
.B(n_5462),
.Y(n_5646)
);

AOI21xp33_ASAP7_75t_L g5647 ( 
.A1(n_5511),
.A2(n_5395),
.B(n_5396),
.Y(n_5647)
);

OAI31xp33_ASAP7_75t_L g5648 ( 
.A1(n_5597),
.A2(n_5397),
.A3(n_5406),
.B(n_5403),
.Y(n_5648)
);

AND2x2_ASAP7_75t_L g5649 ( 
.A(n_5510),
.B(n_5489),
.Y(n_5649)
);

AOI322xp5_ASAP7_75t_L g5650 ( 
.A1(n_5559),
.A2(n_5412),
.A3(n_5409),
.B1(n_5426),
.B2(n_5479),
.C1(n_339),
.C2(n_343),
.Y(n_5650)
);

A2O1A1Ixp33_ASAP7_75t_L g5651 ( 
.A1(n_5629),
.A2(n_5172),
.B(n_5166),
.C(n_5261),
.Y(n_5651)
);

AND2x2_ASAP7_75t_L g5652 ( 
.A(n_5507),
.B(n_5262),
.Y(n_5652)
);

OAI321xp33_ASAP7_75t_L g5653 ( 
.A1(n_5541),
.A2(n_5464),
.A3(n_341),
.B1(n_343),
.B2(n_337),
.C(n_338),
.Y(n_5653)
);

OAI21xp33_ASAP7_75t_L g5654 ( 
.A1(n_5559),
.A2(n_5141),
.B(n_5250),
.Y(n_5654)
);

AND2x2_ASAP7_75t_L g5655 ( 
.A(n_5504),
.B(n_5314),
.Y(n_5655)
);

AOI221xp5_ASAP7_75t_L g5656 ( 
.A1(n_5629),
.A2(n_345),
.B1(n_342),
.B2(n_344),
.C(n_346),
.Y(n_5656)
);

AOI221xp5_ASAP7_75t_L g5657 ( 
.A1(n_5583),
.A2(n_5609),
.B1(n_5607),
.B2(n_5602),
.C(n_5620),
.Y(n_5657)
);

NAND4xp25_ASAP7_75t_SL g5658 ( 
.A(n_5605),
.B(n_347),
.C(n_344),
.D(n_346),
.Y(n_5658)
);

NAND2xp33_ASAP7_75t_R g5659 ( 
.A(n_5538),
.B(n_348),
.Y(n_5659)
);

OA21x2_ASAP7_75t_L g5660 ( 
.A1(n_5512),
.A2(n_5304),
.B(n_5168),
.Y(n_5660)
);

NOR2xp33_ASAP7_75t_L g5661 ( 
.A(n_5571),
.B(n_5580),
.Y(n_5661)
);

OAI221xp5_ASAP7_75t_L g5662 ( 
.A1(n_5563),
.A2(n_353),
.B1(n_350),
.B2(n_351),
.C(n_354),
.Y(n_5662)
);

NAND3xp33_ASAP7_75t_L g5663 ( 
.A(n_5605),
.B(n_353),
.C(n_354),
.Y(n_5663)
);

OAI33xp33_ASAP7_75t_L g5664 ( 
.A1(n_5576),
.A2(n_359),
.A3(n_361),
.B1(n_356),
.B2(n_358),
.B3(n_360),
.Y(n_5664)
);

OAI221xp5_ASAP7_75t_L g5665 ( 
.A1(n_5589),
.A2(n_365),
.B1(n_362),
.B2(n_364),
.C(n_366),
.Y(n_5665)
);

AOI211xp5_ASAP7_75t_L g5666 ( 
.A1(n_5626),
.A2(n_367),
.B(n_365),
.C(n_366),
.Y(n_5666)
);

OAI221xp5_ASAP7_75t_L g5667 ( 
.A1(n_5626),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.C(n_376),
.Y(n_5667)
);

OA21x2_ASAP7_75t_L g5668 ( 
.A1(n_5572),
.A2(n_5568),
.B(n_5548),
.Y(n_5668)
);

AND2x4_ASAP7_75t_L g5669 ( 
.A(n_5564),
.B(n_378),
.Y(n_5669)
);

AO21x2_ASAP7_75t_L g5670 ( 
.A1(n_5572),
.A2(n_380),
.B(n_382),
.Y(n_5670)
);

NOR3xp33_ASAP7_75t_L g5671 ( 
.A(n_5615),
.B(n_383),
.C(n_384),
.Y(n_5671)
);

AND2x4_ASAP7_75t_L g5672 ( 
.A(n_5542),
.B(n_387),
.Y(n_5672)
);

AND2x2_ASAP7_75t_L g5673 ( 
.A(n_5506),
.B(n_388),
.Y(n_5673)
);

AND2x4_ASAP7_75t_L g5674 ( 
.A(n_5515),
.B(n_389),
.Y(n_5674)
);

NAND2xp5_ASAP7_75t_L g5675 ( 
.A(n_5612),
.B(n_391),
.Y(n_5675)
);

OAI33xp33_ASAP7_75t_L g5676 ( 
.A1(n_5616),
.A2(n_401),
.A3(n_404),
.B1(n_392),
.B2(n_394),
.B3(n_402),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_5533),
.Y(n_5677)
);

INVxp67_ASAP7_75t_SL g5678 ( 
.A(n_5608),
.Y(n_5678)
);

AOI22xp33_ASAP7_75t_L g5679 ( 
.A1(n_5633),
.A2(n_5619),
.B1(n_5630),
.B2(n_5611),
.Y(n_5679)
);

OAI21xp33_ASAP7_75t_SL g5680 ( 
.A1(n_5534),
.A2(n_408),
.B(n_409),
.Y(n_5680)
);

OAI322xp33_ASAP7_75t_L g5681 ( 
.A1(n_5630),
.A2(n_408),
.A3(n_410),
.B1(n_411),
.B2(n_412),
.C1(n_413),
.C2(n_414),
.Y(n_5681)
);

CKINVDCx5p33_ASAP7_75t_R g5682 ( 
.A(n_5553),
.Y(n_5682)
);

NAND3xp33_ASAP7_75t_L g5683 ( 
.A(n_5637),
.B(n_410),
.C(n_411),
.Y(n_5683)
);

AOI33xp33_ASAP7_75t_L g5684 ( 
.A1(n_5590),
.A2(n_417),
.A3(n_420),
.B1(n_415),
.B2(n_416),
.B3(n_418),
.Y(n_5684)
);

OAI22xp33_ASAP7_75t_L g5685 ( 
.A1(n_5632),
.A2(n_421),
.B1(n_418),
.B2(n_420),
.Y(n_5685)
);

AOI22xp33_ASAP7_75t_L g5686 ( 
.A1(n_5618),
.A2(n_1737),
.B1(n_1741),
.B2(n_1735),
.Y(n_5686)
);

INVx2_ASAP7_75t_L g5687 ( 
.A(n_5516),
.Y(n_5687)
);

NOR3xp33_ASAP7_75t_L g5688 ( 
.A(n_5521),
.B(n_421),
.C(n_423),
.Y(n_5688)
);

NOR4xp25_ASAP7_75t_L g5689 ( 
.A(n_5622),
.B(n_429),
.C(n_426),
.D(n_428),
.Y(n_5689)
);

INVx2_ASAP7_75t_L g5690 ( 
.A(n_5567),
.Y(n_5690)
);

A2O1A1Ixp33_ASAP7_75t_SL g5691 ( 
.A1(n_5590),
.A2(n_432),
.B(n_430),
.C(n_431),
.Y(n_5691)
);

AOI22xp33_ASAP7_75t_L g5692 ( 
.A1(n_5624),
.A2(n_5591),
.B1(n_5631),
.B2(n_5634),
.Y(n_5692)
);

OR2x2_ASAP7_75t_L g5693 ( 
.A(n_5540),
.B(n_435),
.Y(n_5693)
);

AND2x4_ASAP7_75t_L g5694 ( 
.A(n_5518),
.B(n_437),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_5514),
.Y(n_5695)
);

OAI22xp5_ASAP7_75t_L g5696 ( 
.A1(n_5640),
.A2(n_440),
.B1(n_438),
.B2(n_439),
.Y(n_5696)
);

AND2x2_ASAP7_75t_L g5697 ( 
.A(n_5543),
.B(n_438),
.Y(n_5697)
);

AND2x4_ASAP7_75t_L g5698 ( 
.A(n_5530),
.B(n_439),
.Y(n_5698)
);

INVx5_ASAP7_75t_L g5699 ( 
.A(n_5509),
.Y(n_5699)
);

NAND2xp5_ASAP7_75t_L g5700 ( 
.A(n_5636),
.B(n_5621),
.Y(n_5700)
);

OAI221xp5_ASAP7_75t_L g5701 ( 
.A1(n_5508),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.C(n_446),
.Y(n_5701)
);

INVx2_ASAP7_75t_L g5702 ( 
.A(n_5561),
.Y(n_5702)
);

AOI22xp33_ASAP7_75t_L g5703 ( 
.A1(n_5591),
.A2(n_5621),
.B1(n_5594),
.B2(n_5579),
.Y(n_5703)
);

AOI22xp33_ASAP7_75t_L g5704 ( 
.A1(n_5579),
.A2(n_1761),
.B1(n_1764),
.B2(n_1745),
.Y(n_5704)
);

OAI22xp33_ASAP7_75t_L g5705 ( 
.A1(n_5565),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_5517),
.Y(n_5706)
);

INVx2_ASAP7_75t_L g5707 ( 
.A(n_5547),
.Y(n_5707)
);

AOI22xp33_ASAP7_75t_SL g5708 ( 
.A1(n_5578),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.Y(n_5708)
);

INVx1_ASAP7_75t_L g5709 ( 
.A(n_5522),
.Y(n_5709)
);

INVx1_ASAP7_75t_L g5710 ( 
.A(n_5525),
.Y(n_5710)
);

OR2x2_ASAP7_75t_L g5711 ( 
.A(n_5575),
.B(n_450),
.Y(n_5711)
);

NAND3xp33_ASAP7_75t_L g5712 ( 
.A(n_5637),
.B(n_5557),
.C(n_5556),
.Y(n_5712)
);

AOI221xp5_ASAP7_75t_L g5713 ( 
.A1(n_5623),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.C(n_455),
.Y(n_5713)
);

AOI211xp5_ASAP7_75t_L g5714 ( 
.A1(n_5614),
.A2(n_459),
.B(n_457),
.C(n_458),
.Y(n_5714)
);

OAI211xp5_ASAP7_75t_SL g5715 ( 
.A1(n_5558),
.A2(n_461),
.B(n_457),
.C(n_460),
.Y(n_5715)
);

OA21x2_ASAP7_75t_L g5716 ( 
.A1(n_5581),
.A2(n_462),
.B(n_463),
.Y(n_5716)
);

NAND4xp75_ASAP7_75t_L g5717 ( 
.A(n_5603),
.B(n_465),
.C(n_463),
.D(n_464),
.Y(n_5717)
);

AOI21xp5_ASAP7_75t_L g5718 ( 
.A1(n_5627),
.A2(n_466),
.B(n_467),
.Y(n_5718)
);

OA21x2_ASAP7_75t_L g5719 ( 
.A1(n_5581),
.A2(n_469),
.B(n_470),
.Y(n_5719)
);

AOI22xp33_ASAP7_75t_L g5720 ( 
.A1(n_5599),
.A2(n_1764),
.B1(n_1767),
.B2(n_1761),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_5526),
.Y(n_5721)
);

OAI221xp5_ASAP7_75t_L g5722 ( 
.A1(n_5569),
.A2(n_472),
.B1(n_470),
.B2(n_471),
.C(n_473),
.Y(n_5722)
);

AND2x2_ASAP7_75t_L g5723 ( 
.A(n_5549),
.B(n_474),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_5535),
.Y(n_5724)
);

AOI221xp5_ASAP7_75t_L g5725 ( 
.A1(n_5627),
.A2(n_490),
.B1(n_487),
.B2(n_489),
.C(n_491),
.Y(n_5725)
);

OAI21xp5_ASAP7_75t_SL g5726 ( 
.A1(n_5555),
.A2(n_489),
.B(n_490),
.Y(n_5726)
);

AOI221xp5_ASAP7_75t_L g5727 ( 
.A1(n_5628),
.A2(n_5524),
.B1(n_5593),
.B2(n_5584),
.C(n_5606),
.Y(n_5727)
);

OAI33xp33_ASAP7_75t_L g5728 ( 
.A1(n_5628),
.A2(n_491),
.A3(n_492),
.B1(n_493),
.B2(n_494),
.B3(n_495),
.Y(n_5728)
);

AOI221xp5_ASAP7_75t_L g5729 ( 
.A1(n_5524),
.A2(n_498),
.B1(n_499),
.B2(n_501),
.C(n_502),
.Y(n_5729)
);

OR2x6_ASAP7_75t_L g5730 ( 
.A(n_5586),
.B(n_499),
.Y(n_5730)
);

OA21x2_ASAP7_75t_L g5731 ( 
.A1(n_5570),
.A2(n_5587),
.B(n_5582),
.Y(n_5731)
);

OAI21xp5_ASAP7_75t_L g5732 ( 
.A1(n_5598),
.A2(n_5592),
.B(n_5638),
.Y(n_5732)
);

AOI22xp33_ASAP7_75t_L g5733 ( 
.A1(n_5601),
.A2(n_5635),
.B1(n_5552),
.B2(n_5610),
.Y(n_5733)
);

INVx2_ASAP7_75t_L g5734 ( 
.A(n_5513),
.Y(n_5734)
);

AND2x2_ASAP7_75t_L g5735 ( 
.A(n_5554),
.B(n_503),
.Y(n_5735)
);

OA21x2_ASAP7_75t_L g5736 ( 
.A1(n_5570),
.A2(n_505),
.B(n_506),
.Y(n_5736)
);

OAI33xp33_ASAP7_75t_L g5737 ( 
.A1(n_5560),
.A2(n_507),
.A3(n_511),
.B1(n_512),
.B2(n_515),
.B3(n_518),
.Y(n_5737)
);

OR2x6_ASAP7_75t_L g5738 ( 
.A(n_5562),
.B(n_511),
.Y(n_5738)
);

NAND3xp33_ASAP7_75t_L g5739 ( 
.A(n_5641),
.B(n_518),
.C(n_519),
.Y(n_5739)
);

AOI22xp5_ASAP7_75t_L g5740 ( 
.A1(n_5604),
.A2(n_525),
.B1(n_521),
.B2(n_522),
.Y(n_5740)
);

OAI22xp5_ASAP7_75t_L g5741 ( 
.A1(n_5600),
.A2(n_532),
.B1(n_529),
.B2(n_531),
.Y(n_5741)
);

CKINVDCx5p33_ASAP7_75t_R g5742 ( 
.A(n_5625),
.Y(n_5742)
);

NAND4xp25_ASAP7_75t_L g5743 ( 
.A(n_5534),
.B(n_537),
.C(n_532),
.D(n_536),
.Y(n_5743)
);

NAND2xp5_ASAP7_75t_L g5744 ( 
.A(n_5566),
.B(n_538),
.Y(n_5744)
);

INVxp67_ASAP7_75t_L g5745 ( 
.A(n_5545),
.Y(n_5745)
);

NOR2xp67_ASAP7_75t_L g5746 ( 
.A(n_5669),
.B(n_5585),
.Y(n_5746)
);

INVxp33_ASAP7_75t_L g5747 ( 
.A(n_5661),
.Y(n_5747)
);

INVx2_ASAP7_75t_L g5748 ( 
.A(n_5699),
.Y(n_5748)
);

INVx2_ASAP7_75t_L g5749 ( 
.A(n_5699),
.Y(n_5749)
);

INVx2_ASAP7_75t_L g5750 ( 
.A(n_5699),
.Y(n_5750)
);

AND2x4_ASAP7_75t_L g5751 ( 
.A(n_5643),
.B(n_5577),
.Y(n_5751)
);

INVx2_ASAP7_75t_SL g5752 ( 
.A(n_5682),
.Y(n_5752)
);

NAND2xp5_ASAP7_75t_L g5753 ( 
.A(n_5716),
.B(n_5573),
.Y(n_5753)
);

HB1xp67_ASAP7_75t_L g5754 ( 
.A(n_5670),
.Y(n_5754)
);

AND2x2_ASAP7_75t_L g5755 ( 
.A(n_5649),
.B(n_5574),
.Y(n_5755)
);

HB1xp67_ASAP7_75t_SL g5756 ( 
.A(n_5656),
.Y(n_5756)
);

INVx2_ASAP7_75t_L g5757 ( 
.A(n_5687),
.Y(n_5757)
);

INVx2_ASAP7_75t_L g5758 ( 
.A(n_5690),
.Y(n_5758)
);

INVx1_ASAP7_75t_SL g5759 ( 
.A(n_5742),
.Y(n_5759)
);

NAND2xp5_ASAP7_75t_L g5760 ( 
.A(n_5719),
.B(n_5539),
.Y(n_5760)
);

INVx1_ASAP7_75t_SL g5761 ( 
.A(n_5672),
.Y(n_5761)
);

INVxp67_ASAP7_75t_L g5762 ( 
.A(n_5659),
.Y(n_5762)
);

INVx1_ASAP7_75t_L g5763 ( 
.A(n_5677),
.Y(n_5763)
);

AND2x2_ASAP7_75t_L g5764 ( 
.A(n_5678),
.B(n_5519),
.Y(n_5764)
);

AND2x2_ASAP7_75t_L g5765 ( 
.A(n_5702),
.B(n_5520),
.Y(n_5765)
);

INVx3_ASAP7_75t_L g5766 ( 
.A(n_5694),
.Y(n_5766)
);

NAND2xp5_ASAP7_75t_L g5767 ( 
.A(n_5718),
.B(n_5523),
.Y(n_5767)
);

INVx3_ASAP7_75t_L g5768 ( 
.A(n_5698),
.Y(n_5768)
);

NAND2xp5_ASAP7_75t_L g5769 ( 
.A(n_5727),
.B(n_5642),
.Y(n_5769)
);

NAND2xp5_ASAP7_75t_L g5770 ( 
.A(n_5644),
.B(n_5523),
.Y(n_5770)
);

INVx2_ASAP7_75t_L g5771 ( 
.A(n_5731),
.Y(n_5771)
);

OR2x2_ASAP7_75t_L g5772 ( 
.A(n_5700),
.B(n_5588),
.Y(n_5772)
);

OR2x2_ASAP7_75t_L g5773 ( 
.A(n_5707),
.B(n_5505),
.Y(n_5773)
);

INVxp67_ASAP7_75t_SL g5774 ( 
.A(n_5668),
.Y(n_5774)
);

INVx5_ASAP7_75t_L g5775 ( 
.A(n_5738),
.Y(n_5775)
);

INVx2_ASAP7_75t_L g5776 ( 
.A(n_5731),
.Y(n_5776)
);

NAND2xp5_ASAP7_75t_L g5777 ( 
.A(n_5712),
.B(n_5527),
.Y(n_5777)
);

HB1xp67_ASAP7_75t_L g5778 ( 
.A(n_5736),
.Y(n_5778)
);

INVx1_ASAP7_75t_L g5779 ( 
.A(n_5695),
.Y(n_5779)
);

NAND2xp5_ASAP7_75t_L g5780 ( 
.A(n_5712),
.B(n_5527),
.Y(n_5780)
);

INVx1_ASAP7_75t_L g5781 ( 
.A(n_5706),
.Y(n_5781)
);

NAND2xp5_ASAP7_75t_L g5782 ( 
.A(n_5697),
.B(n_5528),
.Y(n_5782)
);

INVx1_ASAP7_75t_L g5783 ( 
.A(n_5709),
.Y(n_5783)
);

INVx1_ASAP7_75t_L g5784 ( 
.A(n_5710),
.Y(n_5784)
);

AND2x4_ASAP7_75t_L g5785 ( 
.A(n_5734),
.B(n_5546),
.Y(n_5785)
);

NAND2xp5_ASAP7_75t_L g5786 ( 
.A(n_5745),
.B(n_5529),
.Y(n_5786)
);

INVx1_ASAP7_75t_L g5787 ( 
.A(n_5721),
.Y(n_5787)
);

HB1xp67_ASAP7_75t_L g5788 ( 
.A(n_5736),
.Y(n_5788)
);

INVx2_ASAP7_75t_L g5789 ( 
.A(n_5674),
.Y(n_5789)
);

HB1xp67_ASAP7_75t_L g5790 ( 
.A(n_5668),
.Y(n_5790)
);

NAND2xp5_ASAP7_75t_L g5791 ( 
.A(n_5657),
.B(n_5703),
.Y(n_5791)
);

NAND2xp5_ASAP7_75t_L g5792 ( 
.A(n_5679),
.B(n_5529),
.Y(n_5792)
);

HB1xp67_ASAP7_75t_L g5793 ( 
.A(n_5738),
.Y(n_5793)
);

NAND2xp5_ASAP7_75t_L g5794 ( 
.A(n_5680),
.B(n_5537),
.Y(n_5794)
);

AND2x2_ASAP7_75t_L g5795 ( 
.A(n_5723),
.B(n_5551),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5724),
.Y(n_5796)
);

AND2x2_ASAP7_75t_L g5797 ( 
.A(n_5735),
.B(n_5537),
.Y(n_5797)
);

INVx2_ASAP7_75t_SL g5798 ( 
.A(n_5730),
.Y(n_5798)
);

INVxp67_ASAP7_75t_SL g5799 ( 
.A(n_5685),
.Y(n_5799)
);

AND2x4_ASAP7_75t_L g5800 ( 
.A(n_5730),
.B(n_5688),
.Y(n_5800)
);

INVx1_ASAP7_75t_L g5801 ( 
.A(n_5711),
.Y(n_5801)
);

AOI22xp33_ASAP7_75t_SL g5802 ( 
.A1(n_5683),
.A2(n_5639),
.B1(n_5613),
.B2(n_5596),
.Y(n_5802)
);

NAND2xp5_ASAP7_75t_L g5803 ( 
.A(n_5680),
.B(n_5708),
.Y(n_5803)
);

INVx1_ASAP7_75t_L g5804 ( 
.A(n_5675),
.Y(n_5804)
);

AND2x2_ASAP7_75t_L g5805 ( 
.A(n_5733),
.B(n_5544),
.Y(n_5805)
);

NAND2xp5_ASAP7_75t_L g5806 ( 
.A(n_5693),
.B(n_5646),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_5744),
.Y(n_5807)
);

NAND2xp5_ASAP7_75t_L g5808 ( 
.A(n_5689),
.B(n_5544),
.Y(n_5808)
);

INVx2_ASAP7_75t_L g5809 ( 
.A(n_5655),
.Y(n_5809)
);

NAND2xp5_ASAP7_75t_L g5810 ( 
.A(n_5671),
.B(n_5531),
.Y(n_5810)
);

AND2x4_ASAP7_75t_L g5811 ( 
.A(n_5673),
.B(n_5732),
.Y(n_5811)
);

AND2x2_ASAP7_75t_L g5812 ( 
.A(n_5692),
.B(n_5536),
.Y(n_5812)
);

NAND2xp5_ASAP7_75t_L g5813 ( 
.A(n_5739),
.B(n_5531),
.Y(n_5813)
);

INVx1_ASAP7_75t_SL g5814 ( 
.A(n_5717),
.Y(n_5814)
);

AND2x2_ASAP7_75t_L g5815 ( 
.A(n_5652),
.B(n_5532),
.Y(n_5815)
);

AND2x4_ASAP7_75t_L g5816 ( 
.A(n_5683),
.B(n_5550),
.Y(n_5816)
);

NOR2xp33_ASAP7_75t_L g5817 ( 
.A(n_5647),
.B(n_5596),
.Y(n_5817)
);

OR2x2_ASAP7_75t_L g5818 ( 
.A(n_5743),
.B(n_541),
.Y(n_5818)
);

NAND2xp5_ASAP7_75t_L g5819 ( 
.A(n_5705),
.B(n_543),
.Y(n_5819)
);

NOR2xp67_ASAP7_75t_L g5820 ( 
.A(n_5663),
.B(n_546),
.Y(n_5820)
);

NAND2xp5_ASAP7_75t_L g5821 ( 
.A(n_5725),
.B(n_5729),
.Y(n_5821)
);

INVx2_ASAP7_75t_L g5822 ( 
.A(n_5660),
.Y(n_5822)
);

AND2x2_ASAP7_75t_L g5823 ( 
.A(n_5726),
.B(n_547),
.Y(n_5823)
);

NOR2xp67_ASAP7_75t_L g5824 ( 
.A(n_5775),
.B(n_5663),
.Y(n_5824)
);

INVx1_ASAP7_75t_SL g5825 ( 
.A(n_5761),
.Y(n_5825)
);

AO21x2_ASAP7_75t_L g5826 ( 
.A1(n_5774),
.A2(n_5651),
.B(n_5654),
.Y(n_5826)
);

INVx1_ASAP7_75t_L g5827 ( 
.A(n_5790),
.Y(n_5827)
);

INVx3_ASAP7_75t_L g5828 ( 
.A(n_5766),
.Y(n_5828)
);

HB1xp67_ASAP7_75t_L g5829 ( 
.A(n_5775),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_5790),
.Y(n_5830)
);

AND2x2_ASAP7_75t_L g5831 ( 
.A(n_5752),
.B(n_5704),
.Y(n_5831)
);

AND2x4_ASAP7_75t_L g5832 ( 
.A(n_5775),
.B(n_5740),
.Y(n_5832)
);

INVx1_ASAP7_75t_SL g5833 ( 
.A(n_5761),
.Y(n_5833)
);

NAND4xp25_ASAP7_75t_L g5834 ( 
.A(n_5769),
.B(n_5666),
.C(n_5713),
.D(n_5662),
.Y(n_5834)
);

NAND2xp5_ASAP7_75t_L g5835 ( 
.A(n_5762),
.B(n_5714),
.Y(n_5835)
);

NOR2xp33_ASAP7_75t_L g5836 ( 
.A(n_5747),
.B(n_5645),
.Y(n_5836)
);

INVx2_ASAP7_75t_L g5837 ( 
.A(n_5768),
.Y(n_5837)
);

INVx1_ASAP7_75t_L g5838 ( 
.A(n_5793),
.Y(n_5838)
);

OR2x2_ASAP7_75t_L g5839 ( 
.A(n_5794),
.B(n_5772),
.Y(n_5839)
);

NAND2xp5_ASAP7_75t_L g5840 ( 
.A(n_5798),
.B(n_5666),
.Y(n_5840)
);

AOI33xp33_ASAP7_75t_L g5841 ( 
.A1(n_5802),
.A2(n_5814),
.A3(n_5816),
.B1(n_5800),
.B2(n_5812),
.B3(n_5805),
.Y(n_5841)
);

INVxp67_ASAP7_75t_SL g5842 ( 
.A(n_5746),
.Y(n_5842)
);

OAI211xp5_ASAP7_75t_SL g5843 ( 
.A1(n_5791),
.A2(n_5648),
.B(n_5684),
.C(n_5722),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_5754),
.Y(n_5844)
);

AOI222xp33_ASAP7_75t_L g5845 ( 
.A1(n_5820),
.A2(n_5728),
.B1(n_5664),
.B2(n_5676),
.C1(n_5737),
.C2(n_5665),
.Y(n_5845)
);

AOI21xp5_ASAP7_75t_SL g5846 ( 
.A1(n_5803),
.A2(n_5658),
.B(n_5681),
.Y(n_5846)
);

INVx2_ASAP7_75t_L g5847 ( 
.A(n_5748),
.Y(n_5847)
);

INVx2_ASAP7_75t_SL g5848 ( 
.A(n_5749),
.Y(n_5848)
);

NAND3xp33_ASAP7_75t_L g5849 ( 
.A(n_5777),
.B(n_5667),
.C(n_5701),
.Y(n_5849)
);

INVx1_ASAP7_75t_L g5850 ( 
.A(n_5778),
.Y(n_5850)
);

INVx3_ASAP7_75t_L g5851 ( 
.A(n_5750),
.Y(n_5851)
);

INVx3_ASAP7_75t_L g5852 ( 
.A(n_5751),
.Y(n_5852)
);

INVx1_ASAP7_75t_L g5853 ( 
.A(n_5788),
.Y(n_5853)
);

OAI21xp5_ASAP7_75t_L g5854 ( 
.A1(n_5821),
.A2(n_5691),
.B(n_5653),
.Y(n_5854)
);

OR2x2_ASAP7_75t_L g5855 ( 
.A(n_5794),
.B(n_5696),
.Y(n_5855)
);

AOI22xp5_ASAP7_75t_L g5856 ( 
.A1(n_5756),
.A2(n_5715),
.B1(n_5741),
.B2(n_5720),
.Y(n_5856)
);

NAND3xp33_ASAP7_75t_L g5857 ( 
.A(n_5777),
.B(n_5650),
.C(n_5686),
.Y(n_5857)
);

HB1xp67_ASAP7_75t_L g5858 ( 
.A(n_5788),
.Y(n_5858)
);

AOI322xp5_ASAP7_75t_L g5859 ( 
.A1(n_5799),
.A2(n_548),
.A3(n_549),
.B1(n_550),
.B2(n_551),
.C1(n_552),
.C2(n_553),
.Y(n_5859)
);

INVx3_ASAP7_75t_L g5860 ( 
.A(n_5751),
.Y(n_5860)
);

NOR2xp33_ASAP7_75t_L g5861 ( 
.A(n_5759),
.B(n_548),
.Y(n_5861)
);

INVx2_ASAP7_75t_L g5862 ( 
.A(n_5789),
.Y(n_5862)
);

NAND4xp25_ASAP7_75t_L g5863 ( 
.A(n_5817),
.B(n_5780),
.C(n_5806),
.D(n_5818),
.Y(n_5863)
);

INVx1_ASAP7_75t_L g5864 ( 
.A(n_5774),
.Y(n_5864)
);

OR2x2_ASAP7_75t_L g5865 ( 
.A(n_5770),
.B(n_5808),
.Y(n_5865)
);

INVx2_ASAP7_75t_L g5866 ( 
.A(n_5764),
.Y(n_5866)
);

OR2x2_ASAP7_75t_L g5867 ( 
.A(n_5770),
.B(n_556),
.Y(n_5867)
);

AND2x2_ASAP7_75t_L g5868 ( 
.A(n_5797),
.B(n_557),
.Y(n_5868)
);

OR2x2_ASAP7_75t_L g5869 ( 
.A(n_5792),
.B(n_558),
.Y(n_5869)
);

NAND2xp5_ASAP7_75t_L g5870 ( 
.A(n_5811),
.B(n_559),
.Y(n_5870)
);

AND2x2_ASAP7_75t_L g5871 ( 
.A(n_5755),
.B(n_560),
.Y(n_5871)
);

NAND4xp25_ASAP7_75t_L g5872 ( 
.A(n_5780),
.B(n_563),
.C(n_561),
.D(n_562),
.Y(n_5872)
);

INVx2_ASAP7_75t_L g5873 ( 
.A(n_5757),
.Y(n_5873)
);

HB1xp67_ASAP7_75t_L g5874 ( 
.A(n_5771),
.Y(n_5874)
);

INVx2_ASAP7_75t_L g5875 ( 
.A(n_5758),
.Y(n_5875)
);

OAI221xp5_ASAP7_75t_L g5876 ( 
.A1(n_5810),
.A2(n_564),
.B1(n_565),
.B2(n_566),
.C(n_567),
.Y(n_5876)
);

INVx1_ASAP7_75t_L g5877 ( 
.A(n_5782),
.Y(n_5877)
);

AND2x2_ASAP7_75t_L g5878 ( 
.A(n_5795),
.B(n_568),
.Y(n_5878)
);

OR2x2_ASAP7_75t_L g5879 ( 
.A(n_5792),
.B(n_570),
.Y(n_5879)
);

INVx1_ASAP7_75t_L g5880 ( 
.A(n_5786),
.Y(n_5880)
);

INVx2_ASAP7_75t_L g5881 ( 
.A(n_5852),
.Y(n_5881)
);

HB1xp67_ASAP7_75t_L g5882 ( 
.A(n_5829),
.Y(n_5882)
);

AOI32xp33_ASAP7_75t_L g5883 ( 
.A1(n_5843),
.A2(n_5823),
.A3(n_5813),
.B1(n_5767),
.B2(n_5819),
.Y(n_5883)
);

OR2x2_ASAP7_75t_L g5884 ( 
.A(n_5825),
.B(n_5833),
.Y(n_5884)
);

INVx3_ASAP7_75t_L g5885 ( 
.A(n_5860),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5858),
.Y(n_5886)
);

NAND2xp5_ASAP7_75t_L g5887 ( 
.A(n_5842),
.B(n_5801),
.Y(n_5887)
);

INVx1_ASAP7_75t_L g5888 ( 
.A(n_5874),
.Y(n_5888)
);

NAND2xp5_ASAP7_75t_L g5889 ( 
.A(n_5828),
.B(n_5804),
.Y(n_5889)
);

OR2x2_ASAP7_75t_L g5890 ( 
.A(n_5835),
.B(n_5840),
.Y(n_5890)
);

NAND2x1_ASAP7_75t_L g5891 ( 
.A(n_5832),
.B(n_5776),
.Y(n_5891)
);

INVx1_ASAP7_75t_L g5892 ( 
.A(n_5838),
.Y(n_5892)
);

NAND2xp5_ASAP7_75t_L g5893 ( 
.A(n_5824),
.B(n_5807),
.Y(n_5893)
);

INVx2_ASAP7_75t_L g5894 ( 
.A(n_5851),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_5827),
.Y(n_5895)
);

INVx1_ASAP7_75t_L g5896 ( 
.A(n_5830),
.Y(n_5896)
);

INVx2_ASAP7_75t_L g5897 ( 
.A(n_5837),
.Y(n_5897)
);

INVx1_ASAP7_75t_L g5898 ( 
.A(n_5864),
.Y(n_5898)
);

AND2x2_ASAP7_75t_L g5899 ( 
.A(n_5866),
.B(n_5765),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5850),
.Y(n_5900)
);

INVx1_ASAP7_75t_L g5901 ( 
.A(n_5853),
.Y(n_5901)
);

NOR5xp2_ASAP7_75t_L g5902 ( 
.A(n_5857),
.B(n_5849),
.C(n_5863),
.D(n_5834),
.E(n_5876),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5844),
.Y(n_5903)
);

INVx2_ASAP7_75t_SL g5904 ( 
.A(n_5848),
.Y(n_5904)
);

INVx2_ASAP7_75t_L g5905 ( 
.A(n_5847),
.Y(n_5905)
);

OR2x2_ASAP7_75t_L g5906 ( 
.A(n_5839),
.B(n_5753),
.Y(n_5906)
);

NAND2x1_ASAP7_75t_L g5907 ( 
.A(n_5846),
.B(n_5785),
.Y(n_5907)
);

NOR2x1p5_ASAP7_75t_SL g5908 ( 
.A(n_5865),
.B(n_5822),
.Y(n_5908)
);

INVx1_ASAP7_75t_L g5909 ( 
.A(n_5862),
.Y(n_5909)
);

NAND2xp5_ASAP7_75t_L g5910 ( 
.A(n_5841),
.B(n_5763),
.Y(n_5910)
);

HB1xp67_ASAP7_75t_SL g5911 ( 
.A(n_5861),
.Y(n_5911)
);

AND2x2_ASAP7_75t_L g5912 ( 
.A(n_5871),
.B(n_5831),
.Y(n_5912)
);

OR2x2_ASAP7_75t_L g5913 ( 
.A(n_5855),
.B(n_5869),
.Y(n_5913)
);

INVx1_ASAP7_75t_L g5914 ( 
.A(n_5868),
.Y(n_5914)
);

OR2x2_ASAP7_75t_L g5915 ( 
.A(n_5879),
.B(n_5867),
.Y(n_5915)
);

INVx1_ASAP7_75t_SL g5916 ( 
.A(n_5878),
.Y(n_5916)
);

NOR2x1p5_ASAP7_75t_L g5917 ( 
.A(n_5870),
.B(n_5760),
.Y(n_5917)
);

INVx4_ASAP7_75t_L g5918 ( 
.A(n_5873),
.Y(n_5918)
);

OR2x2_ASAP7_75t_L g5919 ( 
.A(n_5875),
.B(n_5773),
.Y(n_5919)
);

NAND2xp5_ASAP7_75t_L g5920 ( 
.A(n_5836),
.B(n_5779),
.Y(n_5920)
);

NAND2xp5_ASAP7_75t_L g5921 ( 
.A(n_5845),
.B(n_5781),
.Y(n_5921)
);

BUFx2_ASAP7_75t_L g5922 ( 
.A(n_5880),
.Y(n_5922)
);

BUFx2_ASAP7_75t_L g5923 ( 
.A(n_5877),
.Y(n_5923)
);

AND2x2_ASAP7_75t_L g5924 ( 
.A(n_5854),
.B(n_5809),
.Y(n_5924)
);

NAND2xp5_ASAP7_75t_L g5925 ( 
.A(n_5859),
.B(n_5783),
.Y(n_5925)
);

OR2x2_ASAP7_75t_L g5926 ( 
.A(n_5849),
.B(n_5784),
.Y(n_5926)
);

OR2x6_ASAP7_75t_L g5927 ( 
.A(n_5854),
.B(n_5787),
.Y(n_5927)
);

HB1xp67_ASAP7_75t_L g5928 ( 
.A(n_5826),
.Y(n_5928)
);

AND2x2_ASAP7_75t_L g5929 ( 
.A(n_5856),
.B(n_5815),
.Y(n_5929)
);

INVx3_ASAP7_75t_L g5930 ( 
.A(n_5826),
.Y(n_5930)
);

INVx1_ASAP7_75t_L g5931 ( 
.A(n_5928),
.Y(n_5931)
);

OR2x2_ASAP7_75t_L g5932 ( 
.A(n_5884),
.B(n_5872),
.Y(n_5932)
);

AND2x4_ASAP7_75t_L g5933 ( 
.A(n_5885),
.B(n_5796),
.Y(n_5933)
);

INVx1_ASAP7_75t_L g5934 ( 
.A(n_5882),
.Y(n_5934)
);

INVx1_ASAP7_75t_L g5935 ( 
.A(n_5886),
.Y(n_5935)
);

INVx1_ASAP7_75t_L g5936 ( 
.A(n_5886),
.Y(n_5936)
);

INVx1_ASAP7_75t_L g5937 ( 
.A(n_5887),
.Y(n_5937)
);

INVx1_ASAP7_75t_L g5938 ( 
.A(n_5930),
.Y(n_5938)
);

NAND4xp25_ASAP7_75t_L g5939 ( 
.A(n_5902),
.B(n_575),
.C(n_576),
.D(n_577),
.Y(n_5939)
);

INVx1_ASAP7_75t_L g5940 ( 
.A(n_5908),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_5891),
.Y(n_5941)
);

INVxp67_ASAP7_75t_L g5942 ( 
.A(n_5911),
.Y(n_5942)
);

NAND2xp5_ASAP7_75t_L g5943 ( 
.A(n_5881),
.B(n_577),
.Y(n_5943)
);

OR2x2_ASAP7_75t_L g5944 ( 
.A(n_5916),
.B(n_579),
.Y(n_5944)
);

AND2x4_ASAP7_75t_L g5945 ( 
.A(n_5894),
.B(n_580),
.Y(n_5945)
);

INVx1_ASAP7_75t_L g5946 ( 
.A(n_5895),
.Y(n_5946)
);

NAND2xp5_ASAP7_75t_L g5947 ( 
.A(n_5904),
.B(n_582),
.Y(n_5947)
);

INVx1_ASAP7_75t_L g5948 ( 
.A(n_5896),
.Y(n_5948)
);

OR2x6_ASAP7_75t_L g5949 ( 
.A(n_5907),
.B(n_582),
.Y(n_5949)
);

OR2x2_ASAP7_75t_L g5950 ( 
.A(n_5913),
.B(n_584),
.Y(n_5950)
);

AND2x2_ASAP7_75t_L g5951 ( 
.A(n_5912),
.B(n_585),
.Y(n_5951)
);

NAND2x1_ASAP7_75t_L g5952 ( 
.A(n_5918),
.B(n_586),
.Y(n_5952)
);

INVx1_ASAP7_75t_L g5953 ( 
.A(n_5900),
.Y(n_5953)
);

NAND2xp5_ASAP7_75t_L g5954 ( 
.A(n_5883),
.B(n_589),
.Y(n_5954)
);

OAI31xp33_ASAP7_75t_L g5955 ( 
.A1(n_5921),
.A2(n_591),
.A3(n_592),
.B(n_594),
.Y(n_5955)
);

INVx1_ASAP7_75t_L g5956 ( 
.A(n_5900),
.Y(n_5956)
);

INVx1_ASAP7_75t_L g5957 ( 
.A(n_5901),
.Y(n_5957)
);

HB1xp67_ASAP7_75t_L g5958 ( 
.A(n_5888),
.Y(n_5958)
);

BUFx2_ASAP7_75t_L g5959 ( 
.A(n_5918),
.Y(n_5959)
);

OR2x2_ASAP7_75t_L g5960 ( 
.A(n_5890),
.B(n_597),
.Y(n_5960)
);

AND2x2_ASAP7_75t_L g5961 ( 
.A(n_5899),
.B(n_5924),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5898),
.Y(n_5962)
);

AOI32xp33_ASAP7_75t_L g5963 ( 
.A1(n_5925),
.A2(n_602),
.A3(n_604),
.B1(n_605),
.B2(n_606),
.Y(n_5963)
);

INVx1_ASAP7_75t_L g5964 ( 
.A(n_5926),
.Y(n_5964)
);

NAND3xp33_ASAP7_75t_L g5965 ( 
.A(n_5910),
.B(n_607),
.C(n_609),
.Y(n_5965)
);

NAND2xp5_ASAP7_75t_L g5966 ( 
.A(n_5929),
.B(n_607),
.Y(n_5966)
);

NAND2x1p5_ASAP7_75t_L g5967 ( 
.A(n_5915),
.B(n_610),
.Y(n_5967)
);

AND2x2_ASAP7_75t_L g5968 ( 
.A(n_5914),
.B(n_611),
.Y(n_5968)
);

INVx2_ASAP7_75t_L g5969 ( 
.A(n_5897),
.Y(n_5969)
);

INVxp67_ASAP7_75t_L g5970 ( 
.A(n_5923),
.Y(n_5970)
);

INVx3_ASAP7_75t_L g5971 ( 
.A(n_5905),
.Y(n_5971)
);

NAND2xp5_ASAP7_75t_L g5972 ( 
.A(n_5892),
.B(n_5917),
.Y(n_5972)
);

INVx3_ASAP7_75t_L g5973 ( 
.A(n_5919),
.Y(n_5973)
);

OA211x2_ASAP7_75t_L g5974 ( 
.A1(n_5952),
.A2(n_5893),
.B(n_5920),
.C(n_5889),
.Y(n_5974)
);

NOR2x1_ASAP7_75t_L g5975 ( 
.A(n_5949),
.B(n_5927),
.Y(n_5975)
);

NAND2xp5_ASAP7_75t_L g5976 ( 
.A(n_5942),
.B(n_5909),
.Y(n_5976)
);

NAND2xp5_ASAP7_75t_L g5977 ( 
.A(n_5961),
.B(n_5909),
.Y(n_5977)
);

NAND2xp5_ASAP7_75t_L g5978 ( 
.A(n_5973),
.B(n_5922),
.Y(n_5978)
);

OR2x2_ASAP7_75t_L g5979 ( 
.A(n_5932),
.B(n_5906),
.Y(n_5979)
);

BUFx3_ASAP7_75t_L g5980 ( 
.A(n_5959),
.Y(n_5980)
);

INVx3_ASAP7_75t_L g5981 ( 
.A(n_5933),
.Y(n_5981)
);

INVx1_ASAP7_75t_L g5982 ( 
.A(n_5938),
.Y(n_5982)
);

INVx1_ASAP7_75t_L g5983 ( 
.A(n_5951),
.Y(n_5983)
);

INVx1_ASAP7_75t_L g5984 ( 
.A(n_5958),
.Y(n_5984)
);

INVx1_ASAP7_75t_L g5985 ( 
.A(n_5931),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5931),
.Y(n_5986)
);

INVx1_ASAP7_75t_L g5987 ( 
.A(n_5934),
.Y(n_5987)
);

INVx1_ASAP7_75t_L g5988 ( 
.A(n_5967),
.Y(n_5988)
);

CKINVDCx5p33_ASAP7_75t_R g5989 ( 
.A(n_5949),
.Y(n_5989)
);

INVxp67_ASAP7_75t_SL g5990 ( 
.A(n_5940),
.Y(n_5990)
);

NAND2xp33_ASAP7_75t_R g5991 ( 
.A(n_5964),
.B(n_5903),
.Y(n_5991)
);

INVx2_ASAP7_75t_L g5992 ( 
.A(n_5941),
.Y(n_5992)
);

NAND2xp5_ASAP7_75t_L g5993 ( 
.A(n_5970),
.B(n_616),
.Y(n_5993)
);

OR2x2_ASAP7_75t_L g5994 ( 
.A(n_5966),
.B(n_617),
.Y(n_5994)
);

INVx1_ASAP7_75t_SL g5995 ( 
.A(n_5941),
.Y(n_5995)
);

OR2x2_ASAP7_75t_L g5996 ( 
.A(n_5950),
.B(n_619),
.Y(n_5996)
);

OR2x2_ASAP7_75t_L g5997 ( 
.A(n_5944),
.B(n_5972),
.Y(n_5997)
);

NAND2xp5_ASAP7_75t_L g5998 ( 
.A(n_5963),
.B(n_619),
.Y(n_5998)
);

NAND2x1_ASAP7_75t_L g5999 ( 
.A(n_5933),
.B(n_5971),
.Y(n_5999)
);

OR2x2_ASAP7_75t_L g6000 ( 
.A(n_5954),
.B(n_5960),
.Y(n_6000)
);

AND2x2_ASAP7_75t_L g6001 ( 
.A(n_5968),
.B(n_5937),
.Y(n_6001)
);

INVx1_ASAP7_75t_L g6002 ( 
.A(n_5953),
.Y(n_6002)
);

INVx1_ASAP7_75t_L g6003 ( 
.A(n_5953),
.Y(n_6003)
);

NOR2xp33_ASAP7_75t_L g6004 ( 
.A(n_5965),
.B(n_621),
.Y(n_6004)
);

INVx2_ASAP7_75t_SL g6005 ( 
.A(n_5945),
.Y(n_6005)
);

INVx3_ASAP7_75t_L g6006 ( 
.A(n_5971),
.Y(n_6006)
);

INVx1_ASAP7_75t_L g6007 ( 
.A(n_5956),
.Y(n_6007)
);

HB1xp67_ASAP7_75t_L g6008 ( 
.A(n_5999),
.Y(n_6008)
);

NAND2xp5_ASAP7_75t_L g6009 ( 
.A(n_6006),
.B(n_5990),
.Y(n_6009)
);

AND2x4_ASAP7_75t_L g6010 ( 
.A(n_5981),
.B(n_5935),
.Y(n_6010)
);

NAND2xp5_ASAP7_75t_L g6011 ( 
.A(n_6006),
.B(n_5939),
.Y(n_6011)
);

OR2x2_ASAP7_75t_L g6012 ( 
.A(n_6005),
.B(n_5969),
.Y(n_6012)
);

OR2x2_ASAP7_75t_L g6013 ( 
.A(n_5978),
.B(n_5947),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_5980),
.Y(n_6014)
);

NAND2xp5_ASAP7_75t_L g6015 ( 
.A(n_5995),
.B(n_5936),
.Y(n_6015)
);

NAND2xp5_ASAP7_75t_SL g6016 ( 
.A(n_5989),
.B(n_5955),
.Y(n_6016)
);

INVx1_ASAP7_75t_L g6017 ( 
.A(n_5977),
.Y(n_6017)
);

NAND3xp33_ASAP7_75t_L g6018 ( 
.A(n_5991),
.B(n_5957),
.C(n_5956),
.Y(n_6018)
);

INVx2_ASAP7_75t_L g6019 ( 
.A(n_5992),
.Y(n_6019)
);

NAND2xp5_ASAP7_75t_L g6020 ( 
.A(n_5984),
.B(n_5983),
.Y(n_6020)
);

INVx2_ASAP7_75t_L g6021 ( 
.A(n_5996),
.Y(n_6021)
);

NAND2xp5_ASAP7_75t_L g6022 ( 
.A(n_5975),
.B(n_5946),
.Y(n_6022)
);

AND2x4_ASAP7_75t_L g6023 ( 
.A(n_5988),
.B(n_5957),
.Y(n_6023)
);

OR2x2_ASAP7_75t_L g6024 ( 
.A(n_5979),
.B(n_5943),
.Y(n_6024)
);

AND2x2_ASAP7_75t_L g6025 ( 
.A(n_6001),
.B(n_5948),
.Y(n_6025)
);

INVx1_ASAP7_75t_L g6026 ( 
.A(n_5976),
.Y(n_6026)
);

AND2x2_ASAP7_75t_L g6027 ( 
.A(n_5987),
.B(n_5962),
.Y(n_6027)
);

NAND2xp5_ASAP7_75t_L g6028 ( 
.A(n_6004),
.B(n_626),
.Y(n_6028)
);

OAI31xp33_ASAP7_75t_L g6029 ( 
.A1(n_5998),
.A2(n_5986),
.A3(n_5985),
.B(n_5993),
.Y(n_6029)
);

NAND2xp5_ASAP7_75t_L g6030 ( 
.A(n_5982),
.B(n_629),
.Y(n_6030)
);

NAND2xp5_ASAP7_75t_L g6031 ( 
.A(n_6002),
.B(n_629),
.Y(n_6031)
);

NAND2x1p5_ASAP7_75t_L g6032 ( 
.A(n_5997),
.B(n_630),
.Y(n_6032)
);

INVx2_ASAP7_75t_L g6033 ( 
.A(n_5994),
.Y(n_6033)
);

AND2x2_ASAP7_75t_L g6034 ( 
.A(n_6000),
.B(n_631),
.Y(n_6034)
);

NAND2xp5_ASAP7_75t_L g6035 ( 
.A(n_6008),
.B(n_6010),
.Y(n_6035)
);

INVx2_ASAP7_75t_SL g6036 ( 
.A(n_6010),
.Y(n_6036)
);

OAI21xp33_ASAP7_75t_L g6037 ( 
.A1(n_6011),
.A2(n_6014),
.B(n_6016),
.Y(n_6037)
);

INVx1_ASAP7_75t_L g6038 ( 
.A(n_6032),
.Y(n_6038)
);

INVx1_ASAP7_75t_L g6039 ( 
.A(n_6009),
.Y(n_6039)
);

OAI31xp33_ASAP7_75t_L g6040 ( 
.A1(n_6018),
.A2(n_6007),
.A3(n_6003),
.B(n_5974),
.Y(n_6040)
);

INVx2_ASAP7_75t_L g6041 ( 
.A(n_6012),
.Y(n_6041)
);

HB1xp67_ASAP7_75t_L g6042 ( 
.A(n_6015),
.Y(n_6042)
);

INVx2_ASAP7_75t_SL g6043 ( 
.A(n_6023),
.Y(n_6043)
);

AOI21xp5_ASAP7_75t_L g6044 ( 
.A1(n_6022),
.A2(n_633),
.B(n_634),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_6025),
.Y(n_6045)
);

NAND4xp25_ASAP7_75t_SL g6046 ( 
.A(n_6029),
.B(n_638),
.C(n_639),
.D(n_640),
.Y(n_6046)
);

CKINVDCx16_ASAP7_75t_R g6047 ( 
.A(n_6024),
.Y(n_6047)
);

AOI22xp33_ASAP7_75t_SL g6048 ( 
.A1(n_6017),
.A2(n_638),
.B1(n_640),
.B2(n_641),
.Y(n_6048)
);

OAI322xp33_ASAP7_75t_L g6049 ( 
.A1(n_6020),
.A2(n_646),
.A3(n_647),
.B1(n_648),
.B2(n_649),
.C1(n_650),
.C2(n_1750),
.Y(n_6049)
);

NAND3x2_ASAP7_75t_L g6050 ( 
.A(n_6013),
.B(n_649),
.C(n_2065),
.Y(n_6050)
);

NAND2xp5_ASAP7_75t_L g6051 ( 
.A(n_6034),
.B(n_1755),
.Y(n_6051)
);

OA22x2_ASAP7_75t_L g6052 ( 
.A1(n_6019),
.A2(n_1755),
.B1(n_1701),
.B2(n_1697),
.Y(n_6052)
);

BUFx2_ASAP7_75t_L g6053 ( 
.A(n_6027),
.Y(n_6053)
);

NAND2xp5_ASAP7_75t_L g6054 ( 
.A(n_6021),
.B(n_1683),
.Y(n_6054)
);

INVx1_ASAP7_75t_L g6055 ( 
.A(n_6030),
.Y(n_6055)
);

OAI21xp33_ASAP7_75t_L g6056 ( 
.A1(n_6026),
.A2(n_2226),
.B(n_1959),
.Y(n_6056)
);

AOI22xp5_ASAP7_75t_L g6057 ( 
.A1(n_6028),
.A2(n_1959),
.B1(n_2309),
.B2(n_2177),
.Y(n_6057)
);

AO21x1_ASAP7_75t_L g6058 ( 
.A1(n_6031),
.A2(n_2153),
.B(n_2267),
.Y(n_6058)
);

INVx1_ASAP7_75t_L g6059 ( 
.A(n_6030),
.Y(n_6059)
);

INVx1_ASAP7_75t_SL g6060 ( 
.A(n_6053),
.Y(n_6060)
);

INVx1_ASAP7_75t_L g6061 ( 
.A(n_6036),
.Y(n_6061)
);

INVx1_ASAP7_75t_L g6062 ( 
.A(n_6043),
.Y(n_6062)
);

OR2x2_ASAP7_75t_L g6063 ( 
.A(n_6047),
.B(n_6033),
.Y(n_6063)
);

NAND2xp5_ASAP7_75t_L g6064 ( 
.A(n_6038),
.B(n_1945),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_6035),
.Y(n_6065)
);

INVx1_ASAP7_75t_L g6066 ( 
.A(n_6042),
.Y(n_6066)
);

AND2x2_ASAP7_75t_L g6067 ( 
.A(n_6041),
.B(n_1586),
.Y(n_6067)
);

INVx1_ASAP7_75t_L g6068 ( 
.A(n_6045),
.Y(n_6068)
);

XOR2x2_ASAP7_75t_L g6069 ( 
.A(n_6050),
.B(n_2153),
.Y(n_6069)
);

NAND2xp5_ASAP7_75t_L g6070 ( 
.A(n_6048),
.B(n_1594),
.Y(n_6070)
);

NAND2xp5_ASAP7_75t_L g6071 ( 
.A(n_6044),
.B(n_6040),
.Y(n_6071)
);

AND2x2_ASAP7_75t_L g6072 ( 
.A(n_6039),
.B(n_1594),
.Y(n_6072)
);

NAND2xp5_ASAP7_75t_L g6073 ( 
.A(n_6037),
.B(n_1945),
.Y(n_6073)
);

INVxp67_ASAP7_75t_L g6074 ( 
.A(n_6046),
.Y(n_6074)
);

INVx1_ASAP7_75t_L g6075 ( 
.A(n_6051),
.Y(n_6075)
);

NOR2x1_ASAP7_75t_L g6076 ( 
.A(n_6049),
.B(n_1945),
.Y(n_6076)
);

NAND2xp5_ASAP7_75t_L g6077 ( 
.A(n_6055),
.B(n_1595),
.Y(n_6077)
);

AND2x2_ASAP7_75t_L g6078 ( 
.A(n_6059),
.B(n_1595),
.Y(n_6078)
);

NAND2xp5_ASAP7_75t_L g6079 ( 
.A(n_6060),
.B(n_6056),
.Y(n_6079)
);

AOI21xp5_ASAP7_75t_L g6080 ( 
.A1(n_6060),
.A2(n_6054),
.B(n_6058),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_6062),
.Y(n_6081)
);

OAI21xp5_ASAP7_75t_L g6082 ( 
.A1(n_6071),
.A2(n_6057),
.B(n_6052),
.Y(n_6082)
);

INVxp67_ASAP7_75t_SL g6083 ( 
.A(n_6063),
.Y(n_6083)
);

NAND2xp5_ASAP7_75t_L g6084 ( 
.A(n_6061),
.B(n_6057),
.Y(n_6084)
);

A2O1A1Ixp33_ASAP7_75t_L g6085 ( 
.A1(n_6066),
.A2(n_2262),
.B(n_2223),
.C(n_1996),
.Y(n_6085)
);

NAND2xp5_ASAP7_75t_L g6086 ( 
.A(n_6074),
.B(n_1595),
.Y(n_6086)
);

INVx1_ASAP7_75t_L g6087 ( 
.A(n_6065),
.Y(n_6087)
);

AOI221xp5_ASAP7_75t_L g6088 ( 
.A1(n_6068),
.A2(n_1614),
.B1(n_1606),
.B2(n_1595),
.C(n_1599),
.Y(n_6088)
);

INVx2_ASAP7_75t_SL g6089 ( 
.A(n_6069),
.Y(n_6089)
);

INVx1_ASAP7_75t_L g6090 ( 
.A(n_6067),
.Y(n_6090)
);

OAI22xp33_ASAP7_75t_L g6091 ( 
.A1(n_6073),
.A2(n_1599),
.B1(n_1700),
.B2(n_1689),
.Y(n_6091)
);

AND2x2_ASAP7_75t_L g6092 ( 
.A(n_6075),
.B(n_1791),
.Y(n_6092)
);

NAND2xp5_ASAP7_75t_L g6093 ( 
.A(n_6076),
.B(n_1791),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_6083),
.Y(n_6094)
);

NAND2xp5_ASAP7_75t_SL g6095 ( 
.A(n_6081),
.B(n_6070),
.Y(n_6095)
);

INVx1_ASAP7_75t_L g6096 ( 
.A(n_6087),
.Y(n_6096)
);

OAI22xp5_ASAP7_75t_L g6097 ( 
.A1(n_6089),
.A2(n_6079),
.B1(n_6084),
.B2(n_6086),
.Y(n_6097)
);

INVx1_ASAP7_75t_L g6098 ( 
.A(n_6092),
.Y(n_6098)
);

AOI221xp5_ASAP7_75t_SL g6099 ( 
.A1(n_6080),
.A2(n_6064),
.B1(n_6077),
.B2(n_6072),
.C(n_6078),
.Y(n_6099)
);

INVx1_ASAP7_75t_L g6100 ( 
.A(n_6093),
.Y(n_6100)
);

INVx1_ASAP7_75t_L g6101 ( 
.A(n_6090),
.Y(n_6101)
);

AOI22xp5_ASAP7_75t_SL g6102 ( 
.A1(n_6082),
.A2(n_2182),
.B1(n_2157),
.B2(n_2147),
.Y(n_6102)
);

OAI22xp5_ASAP7_75t_L g6103 ( 
.A1(n_6085),
.A2(n_6091),
.B1(n_6088),
.B2(n_1996),
.Y(n_6103)
);

AO22x1_ASAP7_75t_L g6104 ( 
.A1(n_6083),
.A2(n_2157),
.B1(n_2147),
.B2(n_2142),
.Y(n_6104)
);

NOR2xp33_ASAP7_75t_L g6105 ( 
.A(n_6096),
.B(n_6101),
.Y(n_6105)
);

NOR3xp33_ASAP7_75t_L g6106 ( 
.A(n_6097),
.B(n_2292),
.C(n_2267),
.Y(n_6106)
);

OAI21xp5_ASAP7_75t_L g6107 ( 
.A1(n_6095),
.A2(n_2022),
.B(n_2031),
.Y(n_6107)
);

XOR2xp5_ASAP7_75t_L g6108 ( 
.A(n_6098),
.B(n_1660),
.Y(n_6108)
);

INVx1_ASAP7_75t_L g6109 ( 
.A(n_6102),
.Y(n_6109)
);

AOI211x1_ASAP7_75t_L g6110 ( 
.A1(n_6104),
.A2(n_6103),
.B(n_6100),
.C(n_6099),
.Y(n_6110)
);

NAND2x1p5_ASAP7_75t_L g6111 ( 
.A(n_6094),
.B(n_1660),
.Y(n_6111)
);

INVx2_ASAP7_75t_L g6112 ( 
.A(n_6094),
.Y(n_6112)
);

INVx2_ASAP7_75t_SL g6113 ( 
.A(n_6094),
.Y(n_6113)
);

INVx1_ASAP7_75t_L g6114 ( 
.A(n_6112),
.Y(n_6114)
);

INVx2_ASAP7_75t_L g6115 ( 
.A(n_6111),
.Y(n_6115)
);

INVx1_ASAP7_75t_L g6116 ( 
.A(n_6108),
.Y(n_6116)
);

OAI211xp5_ASAP7_75t_L g6117 ( 
.A1(n_6110),
.A2(n_2022),
.B(n_2292),
.C(n_2153),
.Y(n_6117)
);

AND2x2_ASAP7_75t_L g6118 ( 
.A(n_6109),
.B(n_1685),
.Y(n_6118)
);

NAND2xp5_ASAP7_75t_L g6119 ( 
.A(n_6106),
.B(n_1799),
.Y(n_6119)
);

NAND3xp33_ASAP7_75t_L g6120 ( 
.A(n_6107),
.B(n_1671),
.C(n_1670),
.Y(n_6120)
);

A2O1A1Ixp33_ASAP7_75t_SL g6121 ( 
.A1(n_6105),
.A2(n_1671),
.B(n_1670),
.C(n_1669),
.Y(n_6121)
);

AOI22xp5_ASAP7_75t_L g6122 ( 
.A1(n_6113),
.A2(n_1670),
.B1(n_1669),
.B2(n_1660),
.Y(n_6122)
);

NOR3x1_ASAP7_75t_L g6123 ( 
.A(n_6113),
.B(n_1845),
.C(n_1977),
.Y(n_6123)
);

AOI211xp5_ASAP7_75t_L g6124 ( 
.A1(n_6105),
.A2(n_2015),
.B(n_2287),
.C(n_2284),
.Y(n_6124)
);

INVxp33_ASAP7_75t_L g6125 ( 
.A(n_6114),
.Y(n_6125)
);

NOR3xp33_ASAP7_75t_L g6126 ( 
.A(n_6116),
.B(n_1845),
.C(n_2287),
.Y(n_6126)
);

NAND2xp5_ASAP7_75t_SL g6127 ( 
.A(n_6115),
.B(n_2015),
.Y(n_6127)
);

INVx2_ASAP7_75t_L g6128 ( 
.A(n_6118),
.Y(n_6128)
);

NOR2x1_ASAP7_75t_L g6129 ( 
.A(n_6117),
.B(n_6120),
.Y(n_6129)
);

OR5x1_ASAP7_75t_L g6130 ( 
.A(n_6123),
.B(n_2006),
.C(n_2278),
.D(n_2263),
.E(n_2242),
.Y(n_6130)
);

NAND3x1_ASAP7_75t_SL g6131 ( 
.A(n_6121),
.B(n_1999),
.C(n_2242),
.Y(n_6131)
);

NOR2x1_ASAP7_75t_L g6132 ( 
.A(n_6119),
.B(n_1999),
.Y(n_6132)
);

NAND3x1_ASAP7_75t_L g6133 ( 
.A(n_6122),
.B(n_1994),
.C(n_2242),
.Y(n_6133)
);

INVx1_ASAP7_75t_L g6134 ( 
.A(n_6124),
.Y(n_6134)
);

NAND2xp5_ASAP7_75t_L g6135 ( 
.A(n_6128),
.B(n_6125),
.Y(n_6135)
);

OAI222xp33_ASAP7_75t_L g6136 ( 
.A1(n_6129),
.A2(n_1958),
.B1(n_2019),
.B2(n_1597),
.C1(n_1616),
.C2(n_1577),
.Y(n_6136)
);

AO22x2_ASAP7_75t_L g6137 ( 
.A1(n_6134),
.A2(n_1981),
.B1(n_2206),
.B2(n_2205),
.Y(n_6137)
);

NOR3xp33_ASAP7_75t_L g6138 ( 
.A(n_6126),
.B(n_2215),
.C(n_2161),
.Y(n_6138)
);

AOI221xp5_ASAP7_75t_L g6139 ( 
.A1(n_6127),
.A2(n_2215),
.B1(n_2161),
.B2(n_2156),
.C(n_2128),
.Y(n_6139)
);

OAI211xp5_ASAP7_75t_SL g6140 ( 
.A1(n_6132),
.A2(n_1952),
.B(n_2123),
.C(n_2109),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_6135),
.Y(n_6141)
);

AND3x4_ASAP7_75t_L g6142 ( 
.A(n_6138),
.B(n_6130),
.C(n_6131),
.Y(n_6142)
);

INVx2_ASAP7_75t_L g6143 ( 
.A(n_6137),
.Y(n_6143)
);

NOR2x1_ASAP7_75t_L g6144 ( 
.A(n_6140),
.B(n_6133),
.Y(n_6144)
);

BUFx2_ASAP7_75t_L g6145 ( 
.A(n_6139),
.Y(n_6145)
);

XNOR2x1_ASAP7_75t_L g6146 ( 
.A(n_6136),
.B(n_1921),
.Y(n_6146)
);

NOR4xp25_ASAP7_75t_L g6147 ( 
.A(n_6141),
.B(n_1921),
.C(n_2102),
.D(n_2095),
.Y(n_6147)
);

INVx1_ASAP7_75t_L g6148 ( 
.A(n_6144),
.Y(n_6148)
);

INVx1_ASAP7_75t_L g6149 ( 
.A(n_6142),
.Y(n_6149)
);

INVxp67_ASAP7_75t_SL g6150 ( 
.A(n_6146),
.Y(n_6150)
);

INVx1_ASAP7_75t_L g6151 ( 
.A(n_6143),
.Y(n_6151)
);

NOR3xp33_ASAP7_75t_L g6152 ( 
.A(n_6145),
.B(n_1947),
.C(n_2102),
.Y(n_6152)
);

NAND3xp33_ASAP7_75t_SL g6153 ( 
.A(n_6141),
.B(n_1912),
.C(n_2094),
.Y(n_6153)
);

AOI22xp5_ASAP7_75t_L g6154 ( 
.A1(n_6148),
.A2(n_1907),
.B1(n_2094),
.B2(n_2088),
.Y(n_6154)
);

NAND2xp5_ASAP7_75t_L g6155 ( 
.A(n_6151),
.B(n_1907),
.Y(n_6155)
);

AOI211x1_ASAP7_75t_L g6156 ( 
.A1(n_6149),
.A2(n_1907),
.B(n_2094),
.C(n_2088),
.Y(n_6156)
);

AO22x1_ASAP7_75t_L g6157 ( 
.A1(n_6150),
.A2(n_2156),
.B1(n_1907),
.B2(n_1947),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_6152),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_6153),
.Y(n_6159)
);

INVx2_ASAP7_75t_L g6160 ( 
.A(n_6147),
.Y(n_6160)
);

AOI22xp5_ASAP7_75t_L g6161 ( 
.A1(n_6148),
.A2(n_2088),
.B1(n_2062),
.B2(n_2051),
.Y(n_6161)
);

AOI21xp5_ASAP7_75t_L g6162 ( 
.A1(n_6148),
.A2(n_2062),
.B(n_2051),
.Y(n_6162)
);

INVx1_ASAP7_75t_L g6163 ( 
.A(n_6148),
.Y(n_6163)
);

HB1xp67_ASAP7_75t_L g6164 ( 
.A(n_6163),
.Y(n_6164)
);

INVxp67_ASAP7_75t_L g6165 ( 
.A(n_6155),
.Y(n_6165)
);

AND3x4_ASAP7_75t_L g6166 ( 
.A(n_6160),
.B(n_2046),
.C(n_2027),
.Y(n_6166)
);

HB1xp67_ASAP7_75t_L g6167 ( 
.A(n_6159),
.Y(n_6167)
);

OAI22x1_ASAP7_75t_L g6168 ( 
.A1(n_6164),
.A2(n_6158),
.B1(n_6161),
.B2(n_6154),
.Y(n_6168)
);

AOI21xp5_ASAP7_75t_L g6169 ( 
.A1(n_6167),
.A2(n_6162),
.B(n_6157),
.Y(n_6169)
);

XNOR2xp5_ASAP7_75t_L g6170 ( 
.A(n_6166),
.B(n_6156),
.Y(n_6170)
);

OAI22xp5_ASAP7_75t_L g6171 ( 
.A1(n_6165),
.A2(n_1977),
.B1(n_2019),
.B2(n_1958),
.Y(n_6171)
);

INVx1_ASAP7_75t_L g6172 ( 
.A(n_6170),
.Y(n_6172)
);

OAI22xp5_ASAP7_75t_SL g6173 ( 
.A1(n_6172),
.A2(n_6168),
.B1(n_6171),
.B2(n_6169),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_6173),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_6174),
.Y(n_6175)
);

INVx1_ASAP7_75t_L g6176 ( 
.A(n_6175),
.Y(n_6176)
);

OA21x2_ASAP7_75t_L g6177 ( 
.A1(n_6176),
.A2(n_1573),
.B(n_1577),
.Y(n_6177)
);

AOI22x1_ASAP7_75t_L g6178 ( 
.A1(n_6177),
.A2(n_1573),
.B1(n_1616),
.B2(n_1629),
.Y(n_6178)
);

OR2x6_ASAP7_75t_L g6179 ( 
.A(n_6178),
.B(n_1616),
.Y(n_6179)
);

AOI221xp5_ASAP7_75t_L g6180 ( 
.A1(n_6179),
.A2(n_1616),
.B1(n_1629),
.B2(n_1635),
.C(n_1662),
.Y(n_6180)
);

AOI211xp5_ASAP7_75t_L g6181 ( 
.A1(n_6180),
.A2(n_1629),
.B(n_1635),
.C(n_1662),
.Y(n_6181)
);


endmodule