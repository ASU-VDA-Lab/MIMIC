module fake_jpeg_23630_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_39),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_36),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_53),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_34),
.A2(n_23),
.B1(n_33),
.B2(n_35),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_67),
.B1(n_23),
.B2(n_33),
.Y(n_83)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx2_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_61),
.C(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_39),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_20),
.B1(n_17),
.B2(n_23),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_53),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_70),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_69),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_20),
.B(n_17),
.Y(n_70)
);

HAxp5_ASAP7_75t_SL g107 ( 
.A(n_71),
.B(n_22),
.CON(n_107),
.SN(n_107)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_74),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_38),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_77),
.B(n_91),
.Y(n_108)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_87),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_18),
.B1(n_28),
.B2(n_31),
.Y(n_117)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_38),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_16),
.C(n_22),
.Y(n_111)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_64),
.B1(n_62),
.B2(n_55),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_37),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_30),
.B1(n_21),
.B2(n_24),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_109),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_45),
.B1(n_67),
.B2(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_42),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_111),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_57),
.B1(n_47),
.B2(n_16),
.Y(n_106)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_107),
.B(n_82),
.Y(n_140)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_47),
.B1(n_24),
.B2(n_28),
.Y(n_113)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_116),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_74),
.A2(n_18),
.B1(n_28),
.B2(n_31),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_120),
.B1(n_78),
.B2(n_72),
.Y(n_134)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_119),
.Y(n_144)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_28),
.B1(n_26),
.B2(n_31),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_122),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_123),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_68),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_129),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_126),
.B(n_133),
.Y(n_152)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_130),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_89),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_91),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_84),
.B1(n_95),
.B2(n_94),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_75),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_143),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_82),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_137),
.B(n_140),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_109),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_93),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_117),
.B1(n_112),
.B2(n_99),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_150),
.A2(n_160),
.B1(n_111),
.B2(n_73),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_114),
.B1(n_78),
.B2(n_72),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_153),
.A2(n_156),
.B1(n_165),
.B2(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_105),
.C(n_121),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_174),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_112),
.B(n_115),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_162),
.B(n_166),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_114),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_159),
.B(n_171),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_124),
.A2(n_102),
.B1(n_116),
.B2(n_84),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_102),
.Y(n_162)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_113),
.B1(n_120),
.B2(n_95),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_123),
.B(n_104),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_101),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_88),
.B1(n_90),
.B2(n_81),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_132),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_126),
.B(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_135),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_184),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_161),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_SL g224 ( 
.A(n_178),
.B(n_194),
.C(n_197),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_170),
.A2(n_142),
.B1(n_144),
.B2(n_129),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_179),
.A2(n_182),
.B1(n_183),
.B2(n_196),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_140),
.B1(n_148),
.B2(n_130),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_161),
.A2(n_129),
.B1(n_101),
.B2(n_81),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_188),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_154),
.B1(n_157),
.B2(n_162),
.Y(n_209)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_189),
.B(n_198),
.Y(n_226)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_193),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_150),
.A2(n_147),
.B1(n_148),
.B2(n_79),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_191),
.A2(n_158),
.B1(n_151),
.B2(n_168),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_192),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_73),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_SL g194 ( 
.A1(n_172),
.A2(n_18),
.B(n_26),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_148),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_199),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_79),
.B1(n_94),
.B2(n_128),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_0),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_138),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_145),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_138),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_201),
.B(n_169),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_222),
.B1(n_220),
.B2(n_184),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_168),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_207),
.B(n_190),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_154),
.C(n_162),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_214),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_209),
.B(n_223),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_177),
.B(n_162),
.CI(n_157),
.CON(n_214),
.SN(n_214)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_199),
.A2(n_166),
.B1(n_153),
.B2(n_152),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_215),
.A2(n_216),
.B1(n_219),
.B2(n_180),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_152),
.B1(n_159),
.B2(n_166),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_166),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_197),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_193),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_225),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_181),
.A2(n_151),
.B(n_169),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_220),
.A2(n_155),
.B1(n_185),
.B2(n_180),
.Y(n_241)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_155),
.B1(n_94),
.B2(n_145),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_51),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_51),
.Y(n_225)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_186),
.B(n_52),
.CI(n_29),
.CON(n_227),
.SN(n_227)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_187),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_200),
.Y(n_228)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

AOI211xp5_ASAP7_75t_SL g230 ( 
.A1(n_217),
.A2(n_197),
.B(n_182),
.C(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_231),
.A2(n_241),
.B1(n_244),
.B2(n_249),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_233),
.A2(n_211),
.B(n_205),
.Y(n_256)
);

OAI21x1_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_189),
.B(n_188),
.Y(n_235)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_242),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_215),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_239),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_202),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_204),
.A2(n_122),
.B1(n_93),
.B2(n_52),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_122),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_245),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_0),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_256),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_202),
.B1(n_216),
.B2(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_249),
.B1(n_248),
.B2(n_245),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_254),
.A2(n_261),
.B1(n_268),
.B2(n_228),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_239),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_259),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_237),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_211),
.B1(n_208),
.B2(n_225),
.Y(n_261)
);

XOR2x2_ASAP7_75t_SL g263 ( 
.A(n_230),
.B(n_214),
.Y(n_263)
);

XNOR2x1_ASAP7_75t_SL g286 ( 
.A(n_263),
.B(n_256),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_223),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_238),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_213),
.C(n_214),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_234),
.C(n_233),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_244),
.A2(n_227),
.B1(n_31),
.B2(n_29),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_275),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_246),
.Y(n_273)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_234),
.B1(n_236),
.B2(n_247),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_227),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_276),
.B(n_283),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_284),
.B1(n_262),
.B2(n_258),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_29),
.C(n_26),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_282),
.C(n_285),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_15),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_259),
.B(n_14),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_0),
.C(n_1),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_252),
.A2(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_1),
.C(n_2),
.Y(n_285)
);

OAI321xp33_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_13),
.A3(n_11),
.B1(n_10),
.B2(n_4),
.C(n_5),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_267),
.C(n_251),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_301),
.C(n_1),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_294),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_281),
.B(n_268),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_296),
.B(n_297),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_271),
.A2(n_263),
.B1(n_250),
.B2(n_265),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_275),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_282),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_284),
.C(n_11),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_280),
.A2(n_11),
.B(n_10),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_313),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_303),
.B(n_306),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

A2O1A1O1Ixp25_ASAP7_75t_L g307 ( 
.A1(n_288),
.A2(n_285),
.B(n_280),
.C(n_278),
.D(n_277),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_308),
.C(n_310),
.Y(n_315)
);

XNOR2x2_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_2),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_289),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_27),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_300),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_290),
.C(n_287),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_318),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_290),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_311),
.C(n_306),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_320),
.B(n_321),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_293),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_293),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_3),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_315),
.B1(n_319),
.B2(n_316),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_327),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_3),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_3),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_329),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_330),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_326),
.C(n_325),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_329),
.C(n_332),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_331),
.C(n_6),
.Y(n_336)
);

A2O1A1O1Ixp25_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_4),
.B(n_6),
.C(n_7),
.D(n_9),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_4),
.B(n_6),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_6),
.B(n_7),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_7),
.C(n_9),
.Y(n_340)
);


endmodule