module fake_netlist_6_382_n_1428 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_152, n_92, n_105, n_227, n_132, n_102, n_204, n_261, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_231, n_40, n_240, n_139, n_41, n_134, n_273, n_95, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1428);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_152;
input n_92;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_231;
input n_40;
input n_240;
input n_139;
input n_41;
input n_134;
input n_273;
input n_95;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1428;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_474;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1382;
wire n_1372;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_934;
wire n_482;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_859;
wire n_570;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_96),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_148),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_245),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_54),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_101),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_302),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_262),
.B(n_11),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_33),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_178),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_144),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_163),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_258),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_113),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_142),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_295),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_133),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_244),
.Y(n_327)
);

BUFx10_ASAP7_75t_L g328 ( 
.A(n_135),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_248),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_124),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_213),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_126),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_217),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_77),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_210),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_117),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_127),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_203),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_57),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_82),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_186),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_56),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_120),
.Y(n_343)
);

BUFx5_ASAP7_75t_L g344 ( 
.A(n_206),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_224),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_27),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_46),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_141),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_3),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_145),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_279),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_215),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_269),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_70),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_242),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_99),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_43),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_253),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_189),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_261),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_129),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_91),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_274),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_180),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_8),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_48),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_263),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_190),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_58),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_125),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_47),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_3),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_229),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_174),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_28),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_64),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_281),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_115),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_28),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_74),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_239),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_299),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_284),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_94),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_168),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_159),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_25),
.Y(n_388)
);

BUFx10_ASAP7_75t_L g389 ( 
.A(n_237),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_200),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_16),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_38),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_39),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_52),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_146),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_283),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_51),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_59),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_L g399 ( 
.A(n_187),
.B(n_193),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_289),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_118),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_236),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_181),
.B(n_121),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_54),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_241),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_191),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_162),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_266),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_300),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_78),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_264),
.Y(n_411)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_67),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_298),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_275),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_212),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_182),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_221),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_61),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_107),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_16),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_110),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_112),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_20),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_27),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_257),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_111),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_167),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_13),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_208),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_51),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_79),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_84),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_209),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_207),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_196),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_170),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_227),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_25),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_109),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_98),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_131),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_108),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_293),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_89),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_172),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_137),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_271),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_100),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_184),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_173),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_87),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_5),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_2),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_95),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_240),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_307),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_202),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_50),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_243),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_31),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_53),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_10),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_197),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_73),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_214),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_104),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_235),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_38),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_139),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_228),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_80),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_103),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_53),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_220),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_34),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_97),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_136),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_230),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_238),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_247),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_194),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_143),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_106),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_192),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_35),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_231),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_34),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_154),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_306),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_140),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_86),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_249),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_255),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_41),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_105),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_251),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_246),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_288),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_161),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_157),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_138),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_204),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_291),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_40),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_36),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_177),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_222),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_278),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_256),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_175),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_276),
.Y(n_511)
);

BUFx5_ASAP7_75t_L g512 ( 
.A(n_234),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_297),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_72),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_46),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_155),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_252),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_273),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_150),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_265),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_52),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_164),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_250),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_41),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_205),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_17),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_223),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_13),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_49),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_233),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_151),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_102),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_394),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_328),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_339),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_468),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_412),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_537)
);

BUFx12f_ASAP7_75t_L g538 ( 
.A(n_420),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_412),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_311),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_386),
.B(n_4),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_5),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_394),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_394),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_394),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_344),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_315),
.B(n_6),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_411),
.B(n_6),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_392),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_346),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_392),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_460),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_344),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_349),
.Y(n_554)
);

OAI22x1_ASAP7_75t_R g555 ( 
.A1(n_393),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_555)
);

BUFx12f_ASAP7_75t_L g556 ( 
.A(n_389),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_454),
.B(n_7),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_349),
.B(n_55),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_460),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_453),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_315),
.B(n_341),
.Y(n_561)
);

OAI22x1_ASAP7_75t_SL g562 ( 
.A1(n_423),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_349),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_349),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_398),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_398),
.Y(n_566)
);

BUFx12f_ASAP7_75t_L g567 ( 
.A(n_437),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_341),
.B(n_459),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_475),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_314),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g571 ( 
.A1(n_329),
.A2(n_378),
.B(n_364),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_398),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_459),
.B(n_12),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_367),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_355),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_398),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_466),
.B(n_60),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_494),
.Y(n_578)
);

OAI21x1_ASAP7_75t_L g579 ( 
.A1(n_390),
.A2(n_63),
.B(n_62),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_437),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_344),
.Y(n_581)
);

OAI22x1_ASAP7_75t_L g582 ( 
.A1(n_529),
.A2(n_376),
.B1(n_388),
.B2(n_373),
.Y(n_582)
);

AND2x6_ASAP7_75t_L g583 ( 
.A(n_466),
.B(n_65),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_391),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_347),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_502),
.B(n_12),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_408),
.B(n_14),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_529),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_451),
.B(n_14),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_466),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_466),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_501),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_318),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_397),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_470),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_404),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_451),
.B(n_15),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_501),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_501),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_501),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_428),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_502),
.B(n_15),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_312),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_430),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_344),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_532),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_532),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_344),
.Y(n_608)
);

BUFx8_ASAP7_75t_L g609 ( 
.A(n_452),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_313),
.B(n_17),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_344),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_461),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_512),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_462),
.Y(n_614)
);

AND2x6_ASAP7_75t_L g615 ( 
.A(n_323),
.B(n_370),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_448),
.B(n_18),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_350),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_358),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_471),
.B(n_18),
.Y(n_619)
);

BUFx12f_ASAP7_75t_L g620 ( 
.A(n_470),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_512),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_512),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_512),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_417),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_487),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_515),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_330),
.B(n_19),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_521),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_319),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_512),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_440),
.Y(n_631)
);

OAI22x1_ASAP7_75t_SL g632 ( 
.A1(n_366),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_632)
);

BUFx12f_ASAP7_75t_L g633 ( 
.A(n_476),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_476),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_490),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_490),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_512),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_316),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_410),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_481),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_499),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_508),
.B(n_21),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_511),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_372),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_327),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_380),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_335),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_340),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_343),
.B(n_22),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_345),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_351),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_354),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_356),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_357),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_360),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_362),
.Y(n_656)
);

OAI21x1_ASAP7_75t_L g657 ( 
.A1(n_374),
.A2(n_68),
.B(n_66),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_352),
.B(n_69),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_424),
.Y(n_659)
);

BUFx12f_ASAP7_75t_L g660 ( 
.A(n_438),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_SL g661 ( 
.A1(n_458),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_363),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_384),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_387),
.Y(n_664)
);

AND2x2_ASAP7_75t_SL g665 ( 
.A(n_402),
.B(n_23),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_407),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_413),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_320),
.Y(n_668)
);

OA21x2_ASAP7_75t_L g669 ( 
.A1(n_418),
.A2(n_24),
.B(n_26),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_330),
.B(n_26),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_467),
.B(n_29),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_321),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_473),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_431),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_432),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_434),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_439),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_444),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_400),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_485),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_504),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_445),
.B(n_30),
.Y(n_682)
);

CKINVDCx11_ASAP7_75t_R g683 ( 
.A(n_414),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_683),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_R g685 ( 
.A(n_540),
.B(n_603),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_563),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_533),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_SL g688 ( 
.A1(n_587),
.A2(n_616),
.B1(n_548),
.B2(n_557),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_549),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_543),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_544),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_668),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_R g693 ( 
.A(n_593),
.B(n_505),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_672),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_535),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_575),
.Y(n_696)
);

AND3x2_ASAP7_75t_L g697 ( 
.A(n_589),
.B(n_467),
.C(n_336),
.Y(n_697)
);

AOI21x1_ASAP7_75t_L g698 ( 
.A1(n_629),
.A2(n_463),
.B(n_446),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_544),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_641),
.B(n_382),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_662),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_679),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_545),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_545),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_549),
.Y(n_705)
);

AOI21x1_ASAP7_75t_L g706 ( 
.A1(n_629),
.A2(n_469),
.B(n_464),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_556),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_585),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_R g709 ( 
.A(n_580),
.B(n_435),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_567),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_620),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_551),
.Y(n_712)
);

AO21x2_ASAP7_75t_L g713 ( 
.A1(n_619),
.A2(n_317),
.B(n_399),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_R g714 ( 
.A(n_593),
.B(n_524),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_551),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_633),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_541),
.A2(n_526),
.B1(n_336),
.B2(n_495),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_660),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_552),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_563),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_552),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_564),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_564),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_566),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_680),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_559),
.Y(n_726)
);

BUFx10_ASAP7_75t_L g727 ( 
.A(n_634),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_617),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_538),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_617),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_566),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_572),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_638),
.Y(n_733)
);

BUFx10_ASAP7_75t_L g734 ( 
.A(n_634),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_641),
.Y(n_735)
);

NOR2xp67_ASAP7_75t_L g736 ( 
.A(n_641),
.B(n_472),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_636),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_R g738 ( 
.A(n_595),
.B(n_322),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_618),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_618),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_572),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_644),
.Y(n_742)
);

NOR2xp67_ASAP7_75t_L g743 ( 
.A(n_635),
.B(n_479),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_644),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_576),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_646),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_576),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_646),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_659),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_590),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_606),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_659),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_534),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_590),
.Y(n_754)
);

BUFx8_ASAP7_75t_L g755 ( 
.A(n_588),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_681),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_561),
.B(n_421),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_631),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_536),
.B(n_32),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_631),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_624),
.B(n_491),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_606),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_609),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_591),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_588),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_607),
.Y(n_766)
);

INVx5_ASAP7_75t_L g767 ( 
.A(n_558),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_561),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_568),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_591),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_598),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_598),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_609),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_599),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_599),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_600),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_578),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_689),
.Y(n_778)
);

INVxp67_ASAP7_75t_SL g779 ( 
.A(n_689),
.Y(n_779)
);

NOR3xp33_ASAP7_75t_SL g780 ( 
.A(n_693),
.B(n_661),
.C(n_627),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_764),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_691),
.B(n_571),
.Y(n_782)
);

BUFx6f_ASAP7_75t_SL g783 ( 
.A(n_727),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_727),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_725),
.B(n_597),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_717),
.A2(n_665),
.B1(n_539),
.B2(n_537),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_757),
.B(n_615),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_700),
.B(n_615),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_693),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_713),
.B(n_615),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_764),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_751),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_705),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_705),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_756),
.B(n_542),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_768),
.B(n_670),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_688),
.B(n_671),
.C(n_673),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_720),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_722),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_723),
.Y(n_800)
);

BUFx6f_ASAP7_75t_SL g801 ( 
.A(n_734),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_734),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_751),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_686),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_L g805 ( 
.A(n_769),
.B(n_658),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_713),
.B(n_643),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_732),
.Y(n_807)
);

AO221x1_ASAP7_75t_L g808 ( 
.A1(n_765),
.A2(n_582),
.B1(n_498),
.B2(n_509),
.C(n_503),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_741),
.Y(n_809)
);

NOR2xp67_ASAP7_75t_L g810 ( 
.A(n_767),
.B(n_554),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_697),
.B(n_643),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_737),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_697),
.B(n_643),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_733),
.B(n_554),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_770),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_709),
.Y(n_816)
);

NAND2xp33_ASAP7_75t_L g817 ( 
.A(n_767),
.B(n_658),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_774),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_686),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_685),
.Y(n_820)
);

NAND2xp33_ASAP7_75t_L g821 ( 
.A(n_767),
.B(n_658),
.Y(n_821)
);

AO221x1_ASAP7_75t_L g822 ( 
.A1(n_712),
.A2(n_522),
.B1(n_527),
.B2(n_525),
.C(n_492),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_687),
.B(n_554),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_762),
.B(n_610),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_776),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_699),
.B(n_592),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_724),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_724),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_703),
.B(n_592),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_704),
.B(n_592),
.Y(n_830)
);

NAND2x1p5_ASAP7_75t_L g831 ( 
.A(n_767),
.B(n_547),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_747),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_766),
.B(n_656),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_747),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_759),
.B(n_648),
.C(n_650),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_691),
.B(n_565),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_731),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_745),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_714),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_750),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_754),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_771),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_739),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_692),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_690),
.B(n_546),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_772),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_709),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_775),
.B(n_649),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_715),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_719),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_694),
.B(n_753),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_743),
.B(n_682),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_736),
.B(n_682),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_738),
.B(n_547),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_698),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_740),
.Y(n_856)
);

NAND2xp33_ASAP7_75t_L g857 ( 
.A(n_742),
.B(n_558),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_706),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_721),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_761),
.B(n_553),
.Y(n_860)
);

INVxp67_ASAP7_75t_SL g861 ( 
.A(n_726),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_758),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_760),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_854),
.A2(n_746),
.B1(n_748),
.B2(n_744),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_L g865 ( 
.A(n_789),
.B(n_752),
.C(n_749),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_833),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_778),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_793),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_794),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_797),
.A2(n_642),
.B1(n_573),
.B2(n_602),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_781),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_791),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_843),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_792),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_785),
.B(n_735),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_803),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_839),
.B(n_779),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_795),
.B(n_586),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_848),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_786),
.A2(n_808),
.B1(n_822),
.B2(n_790),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_827),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_796),
.B(n_852),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_798),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_792),
.Y(n_884)
);

NOR2x1p5_ASAP7_75t_L g885 ( 
.A(n_820),
.B(n_773),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_816),
.B(n_777),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_815),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_856),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_853),
.B(n_586),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_832),
.Y(n_890)
);

AND2x6_ASAP7_75t_L g891 ( 
.A(n_787),
.B(n_602),
.Y(n_891)
);

NAND2x1p5_ASAP7_75t_L g892 ( 
.A(n_844),
.B(n_657),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_828),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_847),
.B(n_695),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_834),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_812),
.B(n_696),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_788),
.B(n_718),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_792),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_799),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_838),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_786),
.A2(n_642),
.B1(n_714),
.B2(n_669),
.Y(n_901)
);

OAI21xp33_ASAP7_75t_L g902 ( 
.A1(n_780),
.A2(n_651),
.B(n_650),
.Y(n_902)
);

NOR2x2_ASAP7_75t_L g903 ( 
.A(n_863),
.B(n_555),
.Y(n_903)
);

INVxp33_ASAP7_75t_SL g904 ( 
.A(n_851),
.Y(n_904)
);

NOR2x2_ASAP7_75t_L g905 ( 
.A(n_859),
.B(n_562),
.Y(n_905)
);

AND2x6_ASAP7_75t_SL g906 ( 
.A(n_862),
.B(n_632),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_861),
.B(n_570),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_806),
.B(n_639),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_844),
.B(n_728),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_SL g910 ( 
.A1(n_784),
.A2(n_730),
.B1(n_701),
.B2(n_708),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_824),
.B(n_702),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_800),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_SL g913 ( 
.A1(n_802),
.A2(n_763),
.B1(n_684),
.B2(n_570),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_811),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_783),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_814),
.B(n_639),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_855),
.B(n_640),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_807),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_813),
.Y(n_919)
);

INVxp67_ASAP7_75t_SL g920 ( 
.A(n_836),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_809),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_835),
.B(n_707),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_835),
.B(n_710),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_831),
.B(n_711),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_818),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_825),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_804),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_845),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_782),
.B(n_676),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_840),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_841),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_842),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_837),
.B(n_716),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_782),
.A2(n_531),
.B1(n_403),
.B2(n_325),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_846),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_805),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_858),
.A2(n_669),
.B1(n_577),
.B2(n_583),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_845),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_804),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_849),
.Y(n_940)
);

INVx5_ASAP7_75t_L g941 ( 
.A(n_804),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_855),
.B(n_640),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_850),
.Y(n_943)
);

INVx4_ASAP7_75t_L g944 ( 
.A(n_837),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_860),
.B(n_558),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_857),
.A2(n_677),
.B1(n_652),
.B2(n_654),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_860),
.B(n_858),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_817),
.A2(n_652),
.B1(n_654),
.B2(n_651),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_819),
.Y(n_949)
);

BUFx12f_ASAP7_75t_L g950 ( 
.A(n_819),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_858),
.B(n_577),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_821),
.B(n_577),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_837),
.B(n_324),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_819),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_826),
.B(n_583),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_884),
.B(n_574),
.Y(n_956)
);

AOI21x1_ASAP7_75t_L g957 ( 
.A1(n_951),
.A2(n_830),
.B(n_829),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_947),
.A2(n_810),
.B(n_823),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_940),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_882),
.B(n_326),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_917),
.A2(n_810),
.B(n_579),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_943),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_928),
.A2(n_583),
.B1(n_666),
.B2(n_655),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_942),
.A2(n_600),
.B(n_581),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_888),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_866),
.B(n_729),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_879),
.A2(n_332),
.B1(n_333),
.B2(n_331),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_886),
.Y(n_968)
);

O2A1O1Ixp5_ASAP7_75t_SL g969 ( 
.A1(n_934),
.A2(n_666),
.B(n_655),
.C(n_574),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_883),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_904),
.B(n_755),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_878),
.B(n_755),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_920),
.A2(n_608),
.B(n_605),
.Y(n_973)
);

NOR2xp67_ASAP7_75t_L g974 ( 
.A(n_889),
.B(n_945),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_890),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_871),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_887),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_SL g978 ( 
.A1(n_955),
.A2(n_613),
.B(n_621),
.C(n_611),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_938),
.B(n_870),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_872),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_930),
.Y(n_981)
);

AOI21xp33_ASAP7_75t_L g982 ( 
.A1(n_877),
.A2(n_337),
.B(n_334),
.Y(n_982)
);

BUFx4f_ASAP7_75t_L g983 ( 
.A(n_950),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_870),
.B(n_338),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_936),
.A2(n_348),
.B1(n_353),
.B2(n_342),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_929),
.A2(n_623),
.B(n_622),
.Y(n_986)
);

AND2x2_ASAP7_75t_SL g987 ( 
.A(n_909),
.B(n_783),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_874),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_902),
.A2(n_637),
.B(n_630),
.C(n_584),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_874),
.Y(n_990)
);

CKINVDCx14_ASAP7_75t_R g991 ( 
.A(n_910),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_902),
.A2(n_936),
.B(n_914),
.C(n_908),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_867),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_868),
.A2(n_584),
.B(n_596),
.C(n_594),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_869),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_864),
.B(n_801),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_873),
.B(n_560),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_907),
.B(n_359),
.Y(n_998)
);

AOI22x1_ASAP7_75t_L g999 ( 
.A1(n_892),
.A2(n_365),
.B1(n_368),
.B2(n_361),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_873),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_875),
.B(n_369),
.Y(n_1001)
);

CKINVDCx16_ASAP7_75t_R g1002 ( 
.A(n_910),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_907),
.B(n_880),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_931),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_901),
.B(n_371),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_929),
.A2(n_377),
.B(n_375),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_890),
.A2(n_596),
.B(n_594),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_894),
.B(n_379),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_932),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_901),
.B(n_381),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_880),
.B(n_383),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_911),
.B(n_385),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_937),
.A2(n_396),
.B(n_395),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_944),
.A2(n_952),
.B(n_916),
.Y(n_1014)
);

AOI21x1_ASAP7_75t_L g1015 ( 
.A1(n_881),
.A2(n_604),
.B(n_601),
.Y(n_1015)
);

NOR2xp67_ASAP7_75t_SL g1016 ( 
.A(n_874),
.B(n_401),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_944),
.A2(n_406),
.B(n_405),
.Y(n_1017)
);

OAI21xp33_ASAP7_75t_L g1018 ( 
.A1(n_865),
.A2(n_604),
.B(n_601),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_891),
.B(n_409),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_SL g1020 ( 
.A1(n_953),
.A2(n_612),
.B(n_626),
.C(n_550),
.Y(n_1020)
);

NAND2xp33_ASAP7_75t_R g1021 ( 
.A(n_919),
.B(n_415),
.Y(n_1021)
);

CKINVDCx6p67_ASAP7_75t_R g1022 ( 
.A(n_876),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_892),
.A2(n_419),
.B(n_416),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_897),
.A2(n_612),
.B(n_626),
.C(n_550),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_896),
.B(n_422),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_935),
.B(n_425),
.Y(n_1026)
);

AOI221xp5_ASAP7_75t_L g1027 ( 
.A1(n_923),
.A2(n_614),
.B1(n_625),
.B2(n_628),
.C(n_569),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_895),
.A2(n_496),
.B(n_427),
.C(n_429),
.Y(n_1028)
);

INVx5_ASAP7_75t_L g1029 ( 
.A(n_891),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_899),
.A2(n_493),
.B(n_433),
.C(n_436),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_R g1031 ( 
.A(n_915),
.B(n_426),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_922),
.B(n_900),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_925),
.A2(n_918),
.B(n_921),
.C(n_912),
.Y(n_1033)
);

INVxp67_ASAP7_75t_L g1034 ( 
.A(n_933),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_961),
.A2(n_949),
.B(n_939),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_965),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_993),
.Y(n_1037)
);

AO21x2_ASAP7_75t_L g1038 ( 
.A1(n_974),
.A2(n_946),
.B(n_926),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_995),
.B(n_898),
.Y(n_1039)
);

INVx8_ASAP7_75t_L g1040 ( 
.A(n_988),
.Y(n_1040)
);

BUFx4f_ASAP7_75t_SL g1041 ( 
.A(n_1022),
.Y(n_1041)
);

AO21x2_ASAP7_75t_L g1042 ( 
.A1(n_974),
.A2(n_946),
.B(n_948),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_988),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_975),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_975),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_988),
.B(n_941),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_1000),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_997),
.Y(n_1048)
);

AND2x6_ASAP7_75t_L g1049 ( 
.A(n_979),
.B(n_948),
.Y(n_1049)
);

INVx6_ASAP7_75t_L g1050 ( 
.A(n_990),
.Y(n_1050)
);

INVx5_ASAP7_75t_SL g1051 ( 
.A(n_990),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_956),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_959),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_962),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_970),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_SL g1056 ( 
.A(n_987),
.Y(n_1056)
);

NAND2x1p5_ASAP7_75t_L g1057 ( 
.A(n_1029),
.B(n_941),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_977),
.Y(n_1058)
);

NAND2x1_ASAP7_75t_L g1059 ( 
.A(n_980),
.B(n_927),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_1003),
.A2(n_891),
.B1(n_893),
.B2(n_913),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_968),
.B(n_906),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_976),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_983),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_998),
.B(n_924),
.Y(n_1064)
);

AO21x2_ASAP7_75t_L g1065 ( 
.A1(n_1014),
.A2(n_891),
.B(n_954),
.Y(n_1065)
);

INVx6_ASAP7_75t_L g1066 ( 
.A(n_956),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_981),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_1034),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_1004),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_1009),
.Y(n_1070)
);

AO21x2_ASAP7_75t_L g1071 ( 
.A1(n_1007),
.A2(n_941),
.B(n_442),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1015),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_957),
.A2(n_885),
.B(n_75),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_1029),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_966),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_960),
.B(n_441),
.Y(n_1076)
);

AO21x2_ASAP7_75t_L g1077 ( 
.A1(n_958),
.A2(n_447),
.B(n_443),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_1033),
.A2(n_76),
.B(n_71),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1032),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_989),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_1029),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_972),
.B(n_81),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_1005),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1010),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_1031),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_1012),
.B(n_906),
.Y(n_1086)
);

BUFx2_ASAP7_75t_SL g1087 ( 
.A(n_1026),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1001),
.B(n_449),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_1011),
.Y(n_1089)
);

BUFx2_ASAP7_75t_SL g1090 ( 
.A(n_1023),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_994),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_973),
.A2(n_85),
.B(n_83),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_969),
.A2(n_999),
.B(n_964),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1019),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_984),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_986),
.A2(n_90),
.B(n_88),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_992),
.B(n_450),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_1025),
.B(n_913),
.Y(n_1098)
);

INVx6_ASAP7_75t_L g1099 ( 
.A(n_1002),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_982),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1024),
.Y(n_1101)
);

OA21x2_ASAP7_75t_L g1102 ( 
.A1(n_963),
.A2(n_456),
.B(n_455),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_971),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1083),
.A2(n_1016),
.B(n_1006),
.Y(n_1104)
);

NAND2x1p5_ASAP7_75t_L g1105 ( 
.A(n_1043),
.B(n_996),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_1081),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_1036),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_1099),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1037),
.Y(n_1109)
);

AO21x1_ASAP7_75t_L g1110 ( 
.A1(n_1098),
.A2(n_1030),
.B(n_1013),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_1040),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_1048),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1053),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1048),
.B(n_1008),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1098),
.A2(n_1018),
.B1(n_991),
.B2(n_1027),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1054),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1049),
.A2(n_664),
.B1(n_678),
.B2(n_675),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1086),
.A2(n_1021),
.B1(n_967),
.B2(n_985),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_1043),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1089),
.B(n_614),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1062),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1049),
.A2(n_663),
.B1(n_675),
.B2(n_645),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_1093),
.A2(n_1028),
.B(n_1017),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1055),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1067),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_1043),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1058),
.Y(n_1127)
);

INVx6_ASAP7_75t_L g1128 ( 
.A(n_1040),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_1047),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1070),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1070),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1049),
.A2(n_664),
.B1(n_647),
.B2(n_678),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1079),
.Y(n_1133)
);

CKINVDCx14_ASAP7_75t_R g1134 ( 
.A(n_1063),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1081),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_SL g1136 ( 
.A1(n_1086),
.A2(n_903),
.B1(n_905),
.B2(n_625),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1089),
.B(n_628),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1075),
.B(n_645),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_1068),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1083),
.A2(n_507),
.B1(n_465),
.B2(n_474),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1072),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1100),
.A2(n_1020),
.B1(n_510),
.B2(n_506),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1044),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1045),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1075),
.B(n_647),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1084),
.A2(n_1095),
.B(n_1088),
.Y(n_1146)
);

OAI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1100),
.A2(n_653),
.B1(n_663),
.B2(n_667),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1049),
.A2(n_653),
.B1(n_667),
.B2(n_674),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1045),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1052),
.B(n_457),
.Y(n_1150)
);

NAND2x1p5_ASAP7_75t_L g1151 ( 
.A(n_1081),
.B(n_978),
.Y(n_1151)
);

INVx4_ASAP7_75t_L g1152 ( 
.A(n_1040),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1049),
.A2(n_530),
.B1(n_523),
.B2(n_520),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1074),
.Y(n_1154)
);

OA21x2_ASAP7_75t_L g1155 ( 
.A1(n_1035),
.A2(n_1078),
.B(n_1073),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1069),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1085),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1039),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1060),
.A2(n_519),
.B1(n_518),
.B2(n_517),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_SL g1160 ( 
.A1(n_1056),
.A2(n_516),
.B1(n_514),
.B2(n_513),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1069),
.Y(n_1161)
);

BUFx12f_ASAP7_75t_L g1162 ( 
.A(n_1063),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_SL g1163 ( 
.A(n_1103),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_1099),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_SL g1165 ( 
.A1(n_1056),
.A2(n_500),
.B1(n_497),
.B2(n_489),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1118),
.A2(n_1115),
.B1(n_1153),
.B2(n_1114),
.Y(n_1166)
);

OAI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1164),
.A2(n_1103),
.B1(n_1064),
.B2(n_1088),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1116),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_R g1169 ( 
.A(n_1134),
.B(n_1041),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1146),
.A2(n_1065),
.B(n_1076),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_1163),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1120),
.B(n_1137),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1110),
.A2(n_1080),
.A3(n_1097),
.B(n_1101),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1157),
.Y(n_1174)
);

CKINVDCx16_ASAP7_75t_R g1175 ( 
.A(n_1162),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1115),
.A2(n_1082),
.B(n_1061),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1124),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1139),
.B(n_1061),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1107),
.B(n_1094),
.Y(n_1179)
);

NAND2xp33_ASAP7_75t_R g1180 ( 
.A(n_1158),
.B(n_1039),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_R g1181 ( 
.A(n_1134),
.B(n_1041),
.Y(n_1181)
);

NOR3xp33_ASAP7_75t_SL g1182 ( 
.A(n_1147),
.B(n_1076),
.C(n_1097),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1109),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1107),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1138),
.B(n_1066),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1119),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1112),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1113),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1121),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1108),
.B(n_1074),
.Y(n_1190)
);

NAND2xp33_ASAP7_75t_R g1191 ( 
.A(n_1129),
.B(n_1102),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_1163),
.Y(n_1192)
);

CKINVDCx11_ASAP7_75t_R g1193 ( 
.A(n_1111),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1145),
.B(n_1066),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1127),
.Y(n_1195)
);

INVxp67_ASAP7_75t_L g1196 ( 
.A(n_1112),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1125),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_1111),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1119),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1133),
.B(n_1087),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1159),
.A2(n_1066),
.B1(n_1091),
.B2(n_1051),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1141),
.Y(n_1202)
);

AO21x2_ASAP7_75t_L g1203 ( 
.A1(n_1104),
.A2(n_1065),
.B(n_1071),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1139),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1117),
.A2(n_1092),
.B(n_1096),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1150),
.B(n_1051),
.Y(n_1206)
);

OR2x6_ASAP7_75t_L g1207 ( 
.A(n_1105),
.B(n_1090),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1150),
.B(n_1051),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1152),
.B(n_1059),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1131),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_R g1211 ( 
.A(n_1128),
.B(n_1050),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1152),
.B(n_1042),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_R g1213 ( 
.A(n_1128),
.B(n_1050),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1153),
.A2(n_1042),
.B1(n_1077),
.B2(n_1038),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1130),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1143),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_SL g1217 ( 
.A1(n_1147),
.A2(n_1057),
.B(n_1038),
.C(n_1046),
.Y(n_1217)
);

NAND2xp33_ASAP7_75t_SL g1218 ( 
.A(n_1119),
.B(n_1077),
.Y(n_1218)
);

CKINVDCx16_ASAP7_75t_R g1219 ( 
.A(n_1156),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1144),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1160),
.B(n_1050),
.Y(n_1221)
);

CKINVDCx16_ASAP7_75t_R g1222 ( 
.A(n_1161),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1160),
.B(n_477),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1172),
.B(n_1171),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1166),
.A2(n_1159),
.B1(n_1165),
.B2(n_1132),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1183),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1187),
.B(n_1105),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_1170),
.A2(n_1155),
.A3(n_1149),
.B(n_1071),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1188),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1221),
.B(n_1154),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1192),
.B(n_1179),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1189),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1212),
.B(n_1207),
.Y(n_1233)
);

OR2x2_ASAP7_75t_L g1234 ( 
.A(n_1196),
.B(n_1140),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1197),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1185),
.B(n_1154),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1194),
.B(n_1184),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1176),
.A2(n_1165),
.B1(n_1122),
.B2(n_1132),
.Y(n_1238)
);

AO21x2_ASAP7_75t_L g1239 ( 
.A1(n_1205),
.A2(n_1203),
.B(n_1217),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1212),
.B(n_1106),
.Y(n_1240)
);

NAND4xp25_ASAP7_75t_L g1241 ( 
.A(n_1178),
.B(n_1136),
.C(n_1148),
.D(n_1117),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1167),
.B(n_1136),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1207),
.B(n_1135),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1198),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1173),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1206),
.B(n_1142),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1204),
.B(n_1210),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1207),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1219),
.B(n_1122),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1176),
.B(n_1148),
.Y(n_1250)
);

AOI222xp33_ASAP7_75t_L g1251 ( 
.A1(n_1223),
.A2(n_478),
.B1(n_480),
.B2(n_482),
.C1(n_483),
.C2(n_484),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1173),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_1174),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1168),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1173),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1202),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1215),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1222),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1200),
.B(n_1123),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1177),
.B(n_1123),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1195),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1186),
.Y(n_1262)
);

INVxp67_ASAP7_75t_L g1263 ( 
.A(n_1180),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1216),
.B(n_1151),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1203),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1208),
.B(n_1126),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1191),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1220),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1169),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1175),
.B(n_1155),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1186),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1193),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1199),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1199),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1190),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1182),
.B(n_486),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1214),
.B(n_1057),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1181),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1190),
.B(n_1201),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1218),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1205),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1233),
.B(n_1248),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_L g1283 ( 
.A(n_1225),
.B(n_1241),
.C(n_1238),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1232),
.Y(n_1284)
);

INVx2_ASAP7_75t_SL g1285 ( 
.A(n_1244),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1232),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1226),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1229),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1243),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1233),
.B(n_1209),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1256),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1230),
.B(n_1211),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1256),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1268),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1227),
.B(n_1213),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1235),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1224),
.B(n_36),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1237),
.B(n_37),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1240),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1244),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1267),
.B(n_37),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1270),
.B(n_1259),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1258),
.Y(n_1303)
);

INVxp67_ASAP7_75t_L g1304 ( 
.A(n_1254),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1231),
.B(n_39),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1268),
.Y(n_1306)
);

AND2x4_ASAP7_75t_SL g1307 ( 
.A(n_1236),
.B(n_92),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1247),
.B(n_42),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1257),
.Y(n_1309)
);

NAND2x1_ASAP7_75t_SL g1310 ( 
.A(n_1276),
.B(n_1280),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1253),
.B(n_1266),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1257),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1240),
.B(n_93),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1260),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1261),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1243),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_SL g1317 ( 
.A(n_1263),
.B(n_488),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1250),
.B(n_42),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1279),
.B(n_44),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1245),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1271),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1225),
.B(n_1251),
.C(n_1242),
.Y(n_1322)
);

NAND3xp33_ASAP7_75t_L g1323 ( 
.A(n_1281),
.B(n_45),
.C(n_48),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1246),
.B(n_45),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1302),
.B(n_1281),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1314),
.B(n_1265),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1287),
.Y(n_1327)
);

CKINVDCx14_ASAP7_75t_R g1328 ( 
.A(n_1303),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1285),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1316),
.B(n_1252),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1316),
.B(n_1255),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1288),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1296),
.B(n_1255),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1282),
.B(n_1239),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1284),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1286),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1291),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1282),
.B(n_1239),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1299),
.B(n_1243),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1309),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1322),
.A2(n_1283),
.B1(n_1323),
.B2(n_1324),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1312),
.B(n_1228),
.Y(n_1342)
);

INVx2_ASAP7_75t_SL g1343 ( 
.A(n_1299),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1304),
.B(n_1228),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1293),
.B(n_1228),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1317),
.A2(n_1249),
.B1(n_1272),
.B2(n_1275),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1294),
.B(n_1228),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1306),
.B(n_1264),
.Y(n_1348)
);

NAND3xp33_ASAP7_75t_L g1349 ( 
.A(n_1317),
.B(n_1318),
.C(n_1301),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1315),
.B(n_1273),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1326),
.B(n_1321),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1327),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1325),
.B(n_1319),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1349),
.B(n_1311),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1346),
.B(n_1295),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1328),
.B(n_1289),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1332),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1341),
.A2(n_1234),
.B1(n_1297),
.B2(n_1300),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1348),
.B(n_1310),
.Y(n_1359)
);

INVxp67_ASAP7_75t_L g1360 ( 
.A(n_1348),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1329),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1335),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1340),
.B(n_1320),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1334),
.A2(n_1272),
.B(n_1307),
.C(n_1313),
.Y(n_1364)
);

CKINVDCx16_ASAP7_75t_R g1365 ( 
.A(n_1339),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1336),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1350),
.B(n_1308),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1337),
.Y(n_1368)
);

AOI33xp33_ASAP7_75t_L g1369 ( 
.A1(n_1344),
.A2(n_1305),
.A3(n_1298),
.B1(n_1292),
.B2(n_1278),
.B3(n_1274),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1366),
.Y(n_1370)
);

AOI21xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1354),
.A2(n_1355),
.B(n_1358),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1352),
.Y(n_1372)
);

OAI21xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1359),
.A2(n_1338),
.B(n_1343),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_SL g1374 ( 
.A1(n_1364),
.A2(n_1329),
.B(n_1262),
.C(n_1277),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1365),
.B(n_1339),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1362),
.A2(n_1342),
.B(n_1345),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1356),
.B(n_1330),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1353),
.A2(n_1290),
.B1(n_1330),
.B2(n_1331),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1357),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1351),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1351),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1361),
.A2(n_1347),
.B1(n_1345),
.B2(n_1333),
.Y(n_1382)
);

OAI21xp33_ASAP7_75t_L g1383 ( 
.A1(n_1371),
.A2(n_1369),
.B(n_1367),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1370),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1374),
.A2(n_1363),
.B(n_1253),
.Y(n_1385)
);

NAND4xp25_ASAP7_75t_SL g1386 ( 
.A(n_1373),
.B(n_1269),
.C(n_1368),
.D(n_1333),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1372),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1379),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1375),
.B(n_1360),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1377),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1380),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1381),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1383),
.B(n_1377),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1390),
.B(n_1389),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1389),
.Y(n_1395)
);

AOI221xp5_ASAP7_75t_L g1396 ( 
.A1(n_1386),
.A2(n_1392),
.B1(n_1391),
.B2(n_1387),
.C(n_1388),
.Y(n_1396)
);

NOR3xp33_ASAP7_75t_L g1397 ( 
.A(n_1385),
.B(n_1382),
.C(n_1378),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1384),
.B(n_1376),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1397),
.A2(n_114),
.B1(n_116),
.B2(n_119),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_SL g1400 ( 
.A(n_1395),
.B(n_122),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1393),
.A2(n_123),
.B1(n_128),
.B2(n_130),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1396),
.A2(n_132),
.B(n_134),
.Y(n_1402)
);

NAND2x1_ASAP7_75t_SL g1403 ( 
.A(n_1394),
.B(n_1398),
.Y(n_1403)
);

OAI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1399),
.A2(n_147),
.B1(n_149),
.B2(n_152),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1402),
.A2(n_153),
.B1(n_156),
.B2(n_158),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_SL g1406 ( 
.A(n_1400),
.B(n_160),
.Y(n_1406)
);

OAI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1403),
.A2(n_165),
.B1(n_166),
.B2(n_169),
.C(n_171),
.Y(n_1407)
);

NOR2x1_ASAP7_75t_L g1408 ( 
.A(n_1407),
.B(n_1401),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1406),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1405),
.Y(n_1410)
);

NAND2x1p5_ASAP7_75t_L g1411 ( 
.A(n_1409),
.B(n_1404),
.Y(n_1411)
);

NAND5xp2_ASAP7_75t_L g1412 ( 
.A(n_1410),
.B(n_176),
.C(n_179),
.D(n_183),
.E(n_185),
.Y(n_1412)
);

OAI221xp5_ASAP7_75t_L g1413 ( 
.A1(n_1408),
.A2(n_188),
.B1(n_195),
.B2(n_198),
.C(n_199),
.Y(n_1413)
);

CKINVDCx16_ASAP7_75t_R g1414 ( 
.A(n_1412),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1411),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1415),
.A2(n_1413),
.B1(n_211),
.B2(n_216),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1414),
.A2(n_201),
.B1(n_218),
.B2(n_219),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1417),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1416),
.A2(n_225),
.B1(n_226),
.B2(n_232),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1419),
.A2(n_254),
.B1(n_259),
.B2(n_260),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1418),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_SL g1422 ( 
.A1(n_1421),
.A2(n_267),
.B1(n_268),
.B2(n_270),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1420),
.A2(n_272),
.B1(n_277),
.B2(n_280),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1422),
.A2(n_282),
.B1(n_285),
.B2(n_286),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1423),
.A2(n_287),
.B(n_290),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1425),
.A2(n_292),
.B1(n_294),
.B2(n_296),
.Y(n_1426)
);

AOI221xp5_ASAP7_75t_L g1427 ( 
.A1(n_1426),
.A2(n_1424),
.B1(n_301),
.B2(n_303),
.C(n_304),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1427),
.A2(n_305),
.B1(n_308),
.B2(n_309),
.Y(n_1428)
);


endmodule