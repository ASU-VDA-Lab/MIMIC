module real_jpeg_18065_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_620;
wire n_456;
wire n_578;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_634;
wire n_153;
wire n_104;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_638;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_572;
wire n_412;
wire n_405;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_602;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_1),
.A2(n_138),
.B1(n_141),
.B2(n_142),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_1),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_1),
.A2(n_141),
.B1(n_174),
.B2(n_178),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_1),
.A2(n_141),
.B1(n_246),
.B2(n_252),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_1),
.A2(n_93),
.B1(n_141),
.B2(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_2),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_2),
.A2(n_65),
.B1(n_106),
.B2(n_157),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_2),
.A2(n_65),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_2),
.A2(n_65),
.B1(n_301),
.B2(n_304),
.Y(n_300)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_3),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_3),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_3),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_4),
.B(n_337),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_4),
.A2(n_336),
.B(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_4),
.Y(n_436)
);

OAI32xp33_ASAP7_75t_L g477 ( 
.A1(n_4),
.A2(n_469),
.A3(n_478),
.B1(n_482),
.B2(n_484),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_4),
.A2(n_158),
.B1(n_436),
.B2(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_4),
.B(n_188),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_4),
.A2(n_193),
.B1(n_598),
.B2(n_606),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_5),
.A2(n_98),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_5),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_5),
.A2(n_360),
.B1(n_395),
.B2(n_396),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_5),
.A2(n_360),
.B1(n_512),
.B2(n_515),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_SL g573 ( 
.A1(n_5),
.A2(n_360),
.B1(n_574),
.B2(n_577),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_6),
.Y(n_82)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_6),
.Y(n_330)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_21),
.B(n_23),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_9),
.Y(n_251)
);

BUFx4f_ASAP7_75t_L g255 ( 
.A(n_9),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_10),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_10),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_10),
.A2(n_106),
.B1(n_264),
.B2(n_316),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_10),
.A2(n_264),
.B1(n_467),
.B2(n_470),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_10),
.A2(n_264),
.B1(n_559),
.B2(n_562),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_11),
.A2(n_105),
.B1(n_110),
.B2(n_111),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_11),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_11),
.A2(n_110),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_11),
.A2(n_110),
.B1(n_212),
.B2(n_216),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_11),
.A2(n_110),
.B1(n_347),
.B2(n_350),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_12),
.A2(n_98),
.B1(n_100),
.B2(n_102),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_12),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_12),
.A2(n_102),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_12),
.A2(n_102),
.B1(n_174),
.B2(n_238),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_12),
.A2(n_102),
.B1(n_342),
.B2(n_345),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_13),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_13),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_13),
.A2(n_223),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_13),
.A2(n_223),
.B1(n_408),
.B2(n_410),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_13),
.A2(n_223),
.B1(n_488),
.B2(n_492),
.Y(n_487)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_14),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_14),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_14),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_15),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_15),
.Y(n_215)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_15),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_15),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_16),
.A2(n_355),
.B1(n_357),
.B2(n_358),
.Y(n_354)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_16),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_16),
.A2(n_358),
.B1(n_422),
.B2(n_426),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_16),
.A2(n_174),
.B1(n_358),
.B2(n_554),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_16),
.A2(n_358),
.B1(n_599),
.B2(n_602),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_17),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_18),
.A2(n_89),
.B1(n_93),
.B2(n_95),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_18),
.A2(n_95),
.B1(n_269),
.B2(n_272),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_18),
.A2(n_95),
.B1(n_370),
.B2(n_375),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_18),
.A2(n_95),
.B1(n_431),
.B2(n_433),
.Y(n_430)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_19),
.Y(n_292)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_19),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_637),
.B(n_640),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_309),
.B(n_630),
.Y(n_25)
);

NOR3xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_279),
.C(n_297),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_225),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21x1_ASAP7_75t_SL g632 ( 
.A1(n_29),
.A2(n_633),
.B(n_634),
.Y(n_632)
);

NOR2xp67_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_164),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_30),
.B(n_164),
.Y(n_634)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_146),
.Y(n_30)
);

INVxp33_ASAP7_75t_SL g296 ( 
.A(n_31),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_69),
.C(n_103),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_32),
.A2(n_155),
.B1(n_161),
.B2(n_162),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_32),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_32),
.B(n_103),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_32),
.B(n_148),
.C(n_162),
.Y(n_293)
);

OA21x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_46),
.B(n_59),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_33),
.A2(n_46),
.B1(n_59),
.B2(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_33),
.B(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_33),
.A2(n_46),
.B1(n_237),
.B2(n_369),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_33),
.A2(n_46),
.B1(n_466),
.B2(n_511),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_33),
.A2(n_46),
.B1(n_549),
.B2(n_553),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_33),
.A2(n_46),
.B1(n_511),
.B2(n_553),
.Y(n_567)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_34),
.A2(n_173),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_34),
.A2(n_210),
.B1(n_407),
.B2(n_411),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_34),
.A2(n_210),
.B1(n_407),
.B2(n_465),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_34),
.B(n_436),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_41),
.B2(n_44),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_40),
.Y(n_200)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_40),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_40),
.Y(n_206)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_40),
.Y(n_344)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_40),
.Y(n_351)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_40),
.Y(n_434)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_40),
.Y(n_546)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_41),
.Y(n_494)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_42),
.Y(n_592)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_43),
.Y(n_536)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_43),
.Y(n_601)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_46),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_46),
.B(n_237),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B1(n_54),
.B2(n_58),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_49),
.Y(n_133)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_50),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_50),
.Y(n_514)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_56),
.Y(n_538)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_64),
.Y(n_469)
);

BUFx12f_ASAP7_75t_L g552 ( 
.A(n_64),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_67),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_68),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_69),
.A2(n_70),
.B1(n_147),
.B2(n_163),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_69),
.A2(n_70),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_70),
.B(n_295),
.C(n_296),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_88),
.B1(n_96),
.B2(n_97),
.Y(n_70)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_71),
.A2(n_88),
.B1(n_96),
.B2(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_71),
.A2(n_96),
.B1(n_221),
.B2(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_71),
.A2(n_96),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_71),
.A2(n_96),
.B1(n_287),
.B2(n_300),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_71),
.A2(n_96),
.B1(n_354),
.B2(n_359),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_71),
.A2(n_96),
.B1(n_261),
.B2(n_359),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_71),
.A2(n_96),
.B1(n_354),
.B2(n_403),
.Y(n_402)
);

AO21x2_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_76),
.B(n_81),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_72),
.A2(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_73),
.Y(n_263)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_81),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g638 ( 
.A1(n_81),
.A2(n_150),
.B(n_639),
.Y(n_638)
);

AO22x2_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_84),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_85),
.Y(n_319)
);

BUFx5_ASAP7_75t_L g335 ( 
.A(n_85),
.Y(n_335)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_86),
.Y(n_427)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_89),
.Y(n_361)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_91),
.Y(n_266)
);

INVx8_ASAP7_75t_L g356 ( 
.A(n_91),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_92),
.Y(n_307)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_96),
.B(n_436),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_98),
.Y(n_224)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_101),
.Y(n_405)
);

OAI22x1_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_115),
.B1(n_137),
.B2(n_145),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_108),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_114),
.Y(n_425)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_114),
.Y(n_527)
);

OAI22x1_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_137),
.B1(n_145),
.B2(n_156),
.Y(n_155)
);

OAI22x1_ASAP7_75t_SL g267 ( 
.A1(n_115),
.A2(n_145),
.B1(n_183),
.B2(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_115),
.A2(n_145),
.B1(n_268),
.B2(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_115),
.A2(n_145),
.B1(n_394),
.B2(n_401),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_115),
.A2(n_145),
.B1(n_394),
.B2(n_421),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_115),
.A2(n_145),
.B1(n_421),
.B2(n_523),
.Y(n_522)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_116),
.A2(n_182),
.B1(n_188),
.B2(n_189),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_116),
.A2(n_188),
.B(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_116),
.A2(n_188),
.B1(n_315),
.B2(n_320),
.Y(n_314)
);

OA21x2_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_124),
.B(n_129),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_123),
.Y(n_481)
);

INVxp33_ASAP7_75t_L g484 ( 
.A(n_124),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g400 ( 
.A(n_128),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_132),
.B1(n_134),
.B2(n_136),
.Y(n_129)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_139),
.Y(n_322)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_147),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_154),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_151),
.Y(n_286)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_156),
.Y(n_284)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.C(n_190),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_166),
.A2(n_169),
.B1(n_170),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_166),
.Y(n_278)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_170),
.A2(n_171),
.B(n_181),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_181),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_186),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_190),
.B(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_207),
.B(n_220),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_192),
.B1(n_220),
.B2(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_191),
.A2(n_192),
.B1(n_209),
.B2(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_201),
.B(n_204),
.Y(n_192)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_193),
.A2(n_201),
.B1(n_340),
.B2(n_346),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_193),
.A2(n_245),
.B1(n_346),
.B2(n_379),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_193),
.A2(n_257),
.B1(n_558),
.B2(n_563),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_193),
.A2(n_573),
.B1(n_598),
.B2(n_610),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_194),
.A2(n_243),
.B1(n_341),
.B2(n_430),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_194),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_196),
.Y(n_381)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_196),
.Y(n_612)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_197),
.Y(n_258)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_200),
.Y(n_576)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_203),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_204),
.Y(n_259)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_206),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_207),
.A2(n_208),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_209),
.Y(n_444)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_215),
.Y(n_409)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_276),
.Y(n_225)
);

NAND2x1_ASAP7_75t_SL g633 ( 
.A(n_226),
.B(n_276),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_232),
.C(n_234),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_228),
.B(n_233),
.Y(n_452)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_234),
.B(n_452),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_260),
.C(n_267),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_235),
.B(n_446),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_240),
.B(n_242),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_236),
.B(n_240),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_242),
.B(n_364),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_256),
.B2(n_259),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_243),
.A2(n_430),
.B1(n_487),
.B2(n_495),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_243),
.A2(n_572),
.B1(n_581),
.B2(n_582),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_250),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_251),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_254),
.Y(n_605)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_255),
.Y(n_561)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_260),
.B(n_267),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_263),
.Y(n_357)
);

INVx3_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_272),
.Y(n_395)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

A2O1A1O1Ixp25_ASAP7_75t_L g631 ( 
.A1(n_280),
.A2(n_298),
.B(n_632),
.C(n_635),
.D(n_636),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_294),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_281),
.B(n_294),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_293),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_285),
.C(n_293),
.Y(n_308)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_308),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_299),
.B(n_308),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_299),
.B(n_638),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_299),
.B(n_638),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_300),
.Y(n_639)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_455),
.B(n_625),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_437),
.C(n_450),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_386),
.B(n_412),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_312),
.B(n_386),
.C(n_627),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_362),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_313),
.B(n_363),
.C(n_365),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_323),
.C(n_352),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_314),
.A2(n_352),
.B1(n_353),
.B2(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_315),
.Y(n_401)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_323),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_339),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_324),
.B(n_339),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_331),
.B(n_336),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_344),
.Y(n_580)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_349),
.Y(n_432)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_349),
.Y(n_562)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx6_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_382),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_366),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_378),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_367),
.A2(n_368),
.B1(n_378),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_369),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_372),
.Y(n_483)
);

INVx5_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_374),
.Y(n_377)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_374),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_374),
.Y(n_555)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_378),
.Y(n_391)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_383),
.B(n_440),
.C(n_441),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_384),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_390),
.C(n_392),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_387),
.B(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_392),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_402),
.C(n_406),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_406),
.Y(n_417)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_402),
.B(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_415),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_413),
.B(n_415),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.C(n_419),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_416),
.B(n_458),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_418),
.B(n_419),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_428),
.C(n_435),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_420),
.B(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

INVx6_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx6_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_428),
.A2(n_429),
.B1(n_435),
.B2(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_435),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_436),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_436),
.B(n_540),
.Y(n_539)
);

OAI21xp33_ASAP7_75t_SL g549 ( 
.A1(n_436),
.A2(n_539),
.B(n_550),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_436),
.B(n_594),
.Y(n_593)
);

A2O1A1O1Ixp25_ASAP7_75t_L g625 ( 
.A1(n_437),
.A2(n_450),
.B(n_626),
.C(n_628),
.D(n_629),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_438),
.B(n_449),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_438),
.B(n_449),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_442),
.Y(n_438)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_439),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_445),
.B1(n_447),
.B2(n_448),
.Y(n_442)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_443),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_448),
.C(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_445),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_453),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_451),
.B(n_453),
.Y(n_629)
);

AOI21x1_ASAP7_75t_L g455 ( 
.A1(n_456),
.A2(n_501),
.B(n_624),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_459),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_457),
.B(n_459),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_464),
.C(n_475),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_460),
.A2(n_461),
.B1(n_504),
.B2(n_505),
.Y(n_503)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_464),
.A2(n_475),
.B1(n_476),
.B2(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_464),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_473),
.Y(n_534)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_485),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_477),
.A2(n_485),
.B1(n_486),
.B2(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_477),
.Y(n_509)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_487),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_500),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_528),
.B(n_623),
.Y(n_501)
);

NOR2xp67_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_507),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_503),
.B(n_507),
.Y(n_623)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_510),
.C(n_521),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_508),
.B(n_620),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_510),
.A2(n_521),
.B1(n_522),
.B2(n_621),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_510),
.Y(n_621)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_519),
.Y(n_540)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_525),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_527),
.Y(n_526)
);

AOI21x1_ASAP7_75t_SL g528 ( 
.A1(n_529),
.A2(n_617),
.B(n_622),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_530),
.A2(n_569),
.B(n_616),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_556),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_531),
.B(n_556),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_547),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_532),
.A2(n_547),
.B1(n_548),
.B2(n_584),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_532),
.Y(n_584)
);

OAI32xp33_ASAP7_75t_L g532 ( 
.A1(n_533),
.A2(n_535),
.A3(n_537),
.B1(n_539),
.B2(n_541),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_537),
.Y(n_542)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_543),
.Y(n_541)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_564),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_557),
.B(n_566),
.C(n_568),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_558),
.Y(n_582)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_565),
.A2(n_566),
.B1(n_567),
.B2(n_568),
.Y(n_564)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_565),
.Y(n_568)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_570),
.A2(n_585),
.B(n_615),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_571),
.B(n_583),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_571),
.B(n_583),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_586),
.A2(n_608),
.B(n_614),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_587),
.B(n_597),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_588),
.B(n_593),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_609),
.B(n_613),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_609),
.B(n_613),
.Y(n_614)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_618),
.B(n_619),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_SL g622 ( 
.A(n_618),
.B(n_619),
.Y(n_622)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_641),
.Y(n_640)
);


endmodule