module real_jpeg_21577_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_40),
.B1(n_42),
.B2(n_53),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_1),
.A2(n_5),
.B1(n_44),
.B2(n_53),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_3),
.B1(n_19),
.B2(n_20),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_2),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_2),
.A2(n_19),
.B1(n_40),
.B2(n_42),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_5),
.B1(n_19),
.B2(n_44),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_3),
.A2(n_7),
.B1(n_20),
.B2(n_28),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_3),
.A2(n_25),
.B(n_28),
.C(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_4),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_5),
.A2(n_10),
.B1(n_41),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_5),
.B(n_73),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_5),
.A2(n_8),
.B1(n_44),
.B2(n_46),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_5),
.A2(n_7),
.B1(n_28),
.B2(n_44),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_5),
.A2(n_7),
.B(n_10),
.Y(n_173)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_7),
.A2(n_28),
.B1(n_40),
.B2(n_42),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_7),
.A2(n_24),
.B(n_31),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_7),
.B(n_21),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_7),
.A2(n_42),
.B(n_49),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_8),
.A2(n_40),
.B1(n_42),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_46),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_9),
.A2(n_20),
.B(n_22),
.C(n_30),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_10),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_11),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_100),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_98),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_83),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_15),
.B(n_83),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_61),
.C(n_67),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_16),
.B(n_61),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_60),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_17),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_17),
.A2(n_60),
.B1(n_85),
.B2(n_96),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_17),
.B(n_117),
.C(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_17),
.A2(n_60),
.B1(n_151),
.B2(n_154),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_17),
.A2(n_60),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_17),
.B(n_228),
.C(n_230),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_21),
.B(n_26),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_18),
.A2(n_21),
.B1(n_81),
.B2(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_22),
.B(n_29),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_23),
.A2(n_48),
.B(n_49),
.C(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_49),
.Y(n_58)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_24),
.A2(n_28),
.B(n_50),
.C(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_27),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_28),
.A2(n_41),
.B(n_42),
.C(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_28),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_28),
.B(n_43),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_28),
.B(n_48),
.Y(n_188)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_47),
.B2(n_59),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_34),
.A2(n_35),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_34),
.B(n_59),
.C(n_60),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_45),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_37),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_43),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_43),
.B1(n_45),
.B2(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_38),
.B(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_38),
.A2(n_43),
.B1(n_79),
.B2(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_43),
.Y(n_38)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_42),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_63),
.B(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_43),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_44),
.B(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_54),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_56),
.B1(n_57),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_55),
.A2(n_66),
.B(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_56),
.B(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_61),
.A2(n_62),
.B(n_64),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_64),
.A2(n_86),
.B1(n_87),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_64),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_64),
.B(n_158),
.C(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_64),
.A2(n_142),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_67),
.A2(n_68),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_75),
.B(n_80),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_80),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_69),
.A2(n_76),
.B1(n_105),
.B2(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_71),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_74),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_72),
.B(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_72),
.A2(n_73),
.B1(n_136),
.B2(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_76),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_78),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_79),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_97),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_86),
.A2(n_87),
.B1(n_117),
.B2(n_153),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_110),
.C(n_117),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_87),
.B(n_142),
.C(n_143),
.Y(n_233)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_93),
.B(n_94),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_121),
.B(n_254),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_118),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_102),
.B(n_118),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.C(n_108),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_103),
.B(n_107),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_108),
.A2(n_109),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_110),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_111),
.A2(n_115),
.B1(n_189),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_111),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_113),
.B(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_114),
.A2(n_135),
.B(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_115),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_115),
.B(n_147),
.C(n_188),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_115),
.A2(n_189),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_115),
.B(n_207),
.C(n_212),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_138),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_117),
.A2(n_128),
.B1(n_129),
.B2(n_153),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_117),
.B(n_129),
.C(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_248),
.B(n_253),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_236),
.B(n_247),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_163),
.B(n_220),
.C(n_235),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_149),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_125),
.B(n_149),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_140),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_137),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_127),
.B(n_137),
.C(n_140),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_129),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_128),
.B(n_133),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_129),
.B(n_172),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

NOR2x1_ASAP7_75t_R g179 ( 
.A(n_147),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_180),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_147),
.A2(n_156),
.B1(n_186),
.B2(n_190),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.C(n_157),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_150),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_155),
.B(n_157),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_170),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_219),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_214),
.B(n_218),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_204),
.B(n_213),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_192),
.B(n_203),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_183),
.B(n_191),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_174),
.B(n_182),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_179),
.B(n_181),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_185),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_194),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_196),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_201),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_206),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_211),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_216),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_221),
.B(n_222),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_233),
.B2(n_234),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_227),
.C(n_234),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_233),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_237),
.B(n_238),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_246),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_244),
.C(n_246),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_250),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);


endmodule