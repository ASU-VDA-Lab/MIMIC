module real_aes_4752_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_1034, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_1035, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_1036, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_1034;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_1035;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_1036;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1016;
wire n_908;
wire n_549;
wire n_376;
wire n_571;
wire n_308;
wire n_491;
wire n_694;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_932;
wire n_1021;
wire n_399;
wire n_700;
wire n_948;
wire n_958;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_994;
wire n_372;
wire n_528;
wire n_495;
wire n_892;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_559;
wire n_976;
wire n_466;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_931;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_284;
wire n_656;
wire n_532;
wire n_1025;
wire n_316;
wire n_755;
wire n_409;
wire n_748;
wire n_860;
wire n_909;
wire n_523;
wire n_996;
wire n_298;
wire n_781;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1008;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_954;
wire n_296;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_1003;
wire n_1028;
wire n_533;
wire n_1000;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_397;
wire n_293;
wire n_749;
wire n_385;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_1001;
wire n_494;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_633;
wire n_520;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_0), .A2(n_679), .B(n_682), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_1), .A2(n_145), .B1(n_406), .B2(n_506), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_2), .A2(n_95), .B1(n_440), .B2(n_457), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_3), .A2(n_53), .B1(n_770), .B2(n_771), .Y(n_769) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_4), .Y(n_722) );
AND2x4_ASAP7_75t_L g733 ( .A(n_4), .B(n_274), .Y(n_733) );
AND2x4_ASAP7_75t_L g738 ( .A(n_4), .B(n_739), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_5), .A2(n_231), .B1(n_420), .B2(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g434 ( .A(n_6), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_7), .A2(n_175), .B1(n_323), .B2(n_328), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_8), .A2(n_160), .B1(n_334), .B2(n_338), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_9), .A2(n_59), .B1(n_318), .B2(n_479), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_10), .A2(n_140), .B1(n_293), .B2(n_318), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_11), .A2(n_193), .B1(n_444), .B2(n_600), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_12), .A2(n_229), .B1(n_444), .B2(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g383 ( .A(n_13), .Y(n_383) );
AO22x1_ASAP7_75t_L g548 ( .A1(n_14), .A2(n_129), .B1(n_549), .B2(n_550), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_15), .A2(n_98), .B1(n_323), .B2(n_527), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_16), .A2(n_81), .B1(n_742), .B2(n_767), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_17), .A2(n_122), .B1(n_348), .B2(n_600), .Y(n_663) );
INVx1_ASAP7_75t_L g488 ( .A(n_18), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_19), .A2(n_247), .B1(n_523), .B2(n_525), .Y(n_553) );
INVx1_ASAP7_75t_L g760 ( .A(n_20), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_21), .A2(n_266), .B1(n_385), .B2(n_574), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_22), .B(n_579), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_23), .A2(n_88), .B1(n_455), .B2(n_479), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_24), .A2(n_180), .B1(n_367), .B2(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_25), .A2(n_159), .B1(n_362), .B2(n_635), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_26), .A2(n_278), .B1(n_348), .B2(n_350), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_27), .A2(n_246), .B1(n_414), .B2(n_420), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_28), .A2(n_71), .B1(n_449), .B2(n_450), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_29), .A2(n_108), .B1(n_367), .B2(n_530), .Y(n_529) );
INVx1_ASAP7_75t_SL g688 ( .A(n_30), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_31), .A2(n_270), .B1(n_454), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_32), .A2(n_174), .B1(n_359), .B2(n_452), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_33), .A2(n_78), .B1(n_730), .B2(n_734), .Y(n_729) );
XOR2x2_ASAP7_75t_L g953 ( .A(n_33), .B(n_954), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_33), .A2(n_994), .B1(n_1026), .B2(n_1028), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_34), .A2(n_73), .B1(n_444), .B2(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g1009 ( .A(n_35), .Y(n_1009) );
INVx1_ASAP7_75t_L g315 ( .A(n_36), .Y(n_315) );
INVxp67_ASAP7_75t_L g378 ( .A(n_36), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_36), .B(n_212), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_37), .A2(n_40), .B1(n_380), .B2(n_430), .C(n_433), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_38), .A2(n_230), .B1(n_549), .B2(n_550), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_39), .A2(n_86), .B1(n_737), .B2(n_749), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_41), .A2(n_158), .B1(n_414), .B2(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g1017 ( .A(n_42), .Y(n_1017) );
INVx1_ASAP7_75t_L g563 ( .A(n_43), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_44), .A2(n_47), .B1(n_523), .B2(n_525), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_45), .A2(n_64), .B1(n_338), .B2(n_445), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_46), .A2(n_223), .B1(n_454), .B2(n_596), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_48), .B(n_300), .Y(n_311) );
INVx1_ASAP7_75t_L g1023 ( .A(n_49), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_50), .A2(n_178), .B1(n_615), .B2(n_616), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_51), .A2(n_116), .B1(n_450), .B2(n_658), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g536 ( .A1(n_52), .A2(n_491), .B(n_537), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_54), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_55), .A2(n_281), .B1(n_746), .B2(n_747), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_56), .A2(n_128), .B1(n_523), .B2(n_1001), .Y(n_1000) );
INVxp67_ASAP7_75t_R g762 ( .A(n_57), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_58), .A2(n_277), .B1(n_444), .B2(n_458), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_60), .A2(n_163), .B1(n_454), .B2(n_455), .Y(n_453) );
INVx2_ASAP7_75t_L g720 ( .A(n_61), .Y(n_720) );
INVx1_ASAP7_75t_L g964 ( .A(n_62), .Y(n_964) );
INVx1_ASAP7_75t_L g732 ( .A(n_63), .Y(n_732) );
AND2x4_ASAP7_75t_L g735 ( .A(n_63), .B(n_720), .Y(n_735) );
INVx1_ASAP7_75t_SL g768 ( .A(n_63), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_65), .A2(n_205), .B1(n_348), .B2(n_458), .Y(n_475) );
INVx1_ASAP7_75t_L g966 ( .A(n_66), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_67), .A2(n_244), .B1(n_974), .B2(n_976), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_68), .A2(n_210), .B1(n_440), .B2(n_441), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_69), .B(n_532), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_70), .A2(n_239), .B1(n_328), .B2(n_481), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_72), .A2(n_573), .B(n_576), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_74), .A2(n_199), .B1(n_742), .B2(n_767), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_75), .A2(n_132), .B1(n_457), .B2(n_458), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_76), .A2(n_217), .B1(n_338), .B2(n_445), .Y(n_673) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_77), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_79), .A2(n_109), .B1(n_525), .B2(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_80), .A2(n_120), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
INVx1_ASAP7_75t_L g686 ( .A(n_81), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_82), .B(n_409), .Y(n_507) );
XOR2x2_ASAP7_75t_L g611 ( .A(n_83), .B(n_612), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_84), .A2(n_102), .B1(n_585), .B2(n_587), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_85), .A2(n_155), .B1(n_449), .B2(n_633), .Y(n_632) );
AO22x2_ASAP7_75t_L g1006 ( .A1(n_87), .A2(n_188), .B1(n_293), .B2(n_1007), .Y(n_1006) );
CKINVDCx16_ASAP7_75t_R g758 ( .A(n_89), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_90), .A2(n_179), .B1(n_737), .B2(n_740), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_91), .A2(n_194), .B1(n_491), .B2(n_492), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_92), .A2(n_218), .B1(n_423), .B2(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g301 ( .A(n_93), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_93), .B(n_211), .Y(n_375) );
AOI33xp33_ASAP7_75t_R g627 ( .A1(n_94), .A2(n_242), .A3(n_336), .B1(n_340), .B2(n_628), .B3(n_1036), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_96), .A2(n_255), .B1(n_369), .B2(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_97), .A2(n_245), .B1(n_559), .B2(n_988), .Y(n_1024) );
AOI21xp5_ASAP7_75t_SL g484 ( .A1(n_99), .A2(n_485), .B(n_487), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_100), .A2(n_150), .B1(n_481), .B2(n_527), .Y(n_547) );
INVx1_ASAP7_75t_L g427 ( .A(n_101), .Y(n_427) );
OAI222xp33_ASAP7_75t_L g446 ( .A1(n_101), .A2(n_447), .B1(n_453), .B2(n_456), .C1(n_1034), .C2(n_1035), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_101), .B(n_456), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_103), .A2(n_110), .B1(n_406), .B2(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g399 ( .A(n_104), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_105), .A2(n_254), .B1(n_479), .B2(n_624), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_106), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_107), .A2(n_209), .B1(n_417), .B2(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g515 ( .A(n_111), .Y(n_515) );
XNOR2x2_ASAP7_75t_L g646 ( .A(n_112), .B(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_113), .A2(n_267), .B1(n_328), .B2(n_457), .Y(n_672) );
INVx1_ASAP7_75t_L g703 ( .A(n_114), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_115), .A2(n_181), .B1(n_730), .B2(n_747), .Y(n_774) );
INVx1_ASAP7_75t_L g790 ( .A(n_117), .Y(n_790) );
INVx1_ASAP7_75t_L g511 ( .A(n_118), .Y(n_511) );
INVx1_ASAP7_75t_L g983 ( .A(n_119), .Y(n_983) );
AOI21xp33_ASAP7_75t_L g509 ( .A1(n_121), .A2(n_403), .B(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_123), .A2(n_269), .B1(n_417), .B2(n_418), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_124), .A2(n_154), .B1(n_338), .B2(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g970 ( .A(n_125), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_126), .A2(n_161), .B1(n_403), .B2(n_404), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_127), .A2(n_166), .B1(n_530), .B2(n_615), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_130), .A2(n_248), .B1(n_338), .B2(n_445), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_131), .A2(n_214), .B1(n_494), .B2(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_133), .A2(n_197), .B1(n_362), .B2(n_656), .Y(n_655) );
AO22x1_ASAP7_75t_L g443 ( .A1(n_134), .A2(n_135), .B1(n_444), .B2(n_445), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_136), .A2(n_198), .B1(n_415), .B2(n_421), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_137), .A2(n_144), .B1(n_454), .B2(n_455), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g977 ( .A1(n_138), .A2(n_236), .B1(n_978), .B2(n_980), .Y(n_977) );
CKINVDCx16_ASAP7_75t_R g394 ( .A(n_139), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_141), .A2(n_157), .B1(n_423), .B2(n_424), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_142), .B(n_359), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_143), .A2(n_186), .B1(n_734), .B2(n_746), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_146), .A2(n_162), .B1(n_380), .B2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_147), .A2(n_261), .B1(n_454), .B2(n_455), .Y(n_662) );
INVx1_ASAP7_75t_L g1018 ( .A(n_148), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_149), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g683 ( .A(n_151), .Y(n_683) );
INVx1_ASAP7_75t_L g1014 ( .A(n_152), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_153), .A2(n_226), .B1(n_367), .B2(n_369), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g956 ( .A1(n_156), .A2(n_238), .B1(n_957), .B2(n_958), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_164), .A2(n_276), .B1(n_334), .B2(n_338), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_165), .A2(n_252), .B1(n_770), .B2(n_771), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_167), .A2(n_204), .B1(n_481), .B2(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g793 ( .A(n_168), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_169), .A2(n_253), .B1(n_359), .B2(n_362), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_170), .A2(n_206), .B1(n_432), .B2(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g791 ( .A(n_171), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_172), .A2(n_280), .B1(n_452), .B2(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g969 ( .A(n_173), .Y(n_969) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_176), .A2(n_380), .B(n_382), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_177), .A2(n_224), .B1(n_338), .B2(n_445), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_182), .A2(n_192), .B1(n_530), .B2(n_557), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_183), .A2(n_570), .B1(n_601), .B2(n_602), .Y(n_569) );
INVx1_ASAP7_75t_L g601 ( .A(n_183), .Y(n_601) );
AOI22x1_ASAP7_75t_L g603 ( .A1(n_183), .A2(n_570), .B1(n_601), .B2(n_602), .Y(n_603) );
INVx1_ASAP7_75t_L g577 ( .A(n_184), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_185), .A2(n_216), .B1(n_367), .B2(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_187), .B(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_189), .B(n_385), .Y(n_684) );
INVx1_ASAP7_75t_L g645 ( .A(n_190), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_191), .A2(n_265), .B1(n_318), .B2(n_479), .Y(n_552) );
OA22x2_ASAP7_75t_L g306 ( .A1(n_195), .A2(n_212), .B1(n_300), .B2(n_304), .Y(n_306) );
INVx1_ASAP7_75t_L g344 ( .A(n_195), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_196), .A2(n_262), .B1(n_385), .B2(n_409), .Y(n_408) );
NAND2xp33_ASAP7_75t_L g354 ( .A(n_200), .B(n_355), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_201), .A2(n_259), .B1(n_328), .B2(n_593), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_202), .A2(n_243), .B1(n_338), .B2(n_549), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_203), .A2(n_220), .B1(n_440), .B2(n_457), .Y(n_692) );
INVx1_ASAP7_75t_L g705 ( .A(n_207), .Y(n_705) );
CKINVDCx6p67_ASAP7_75t_R g756 ( .A(n_208), .Y(n_756) );
INVx1_ASAP7_75t_L g317 ( .A(n_211), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_211), .B(n_342), .Y(n_393) );
OAI21xp33_ASAP7_75t_L g345 ( .A1(n_212), .A2(n_227), .B(n_346), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_213), .A2(n_235), .B1(n_407), .B2(n_411), .Y(n_508) );
XNOR2x1_ASAP7_75t_L g497 ( .A(n_215), .B(n_498), .Y(n_497) );
XNOR2x2_ASAP7_75t_SL g512 ( .A(n_215), .B(n_498), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_219), .A2(n_279), .B1(n_737), .B2(n_749), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_221), .A2(n_995), .B1(n_996), .B2(n_1025), .Y(n_994) );
CKINVDCx5p33_ASAP7_75t_R g995 ( .A(n_221), .Y(n_995) );
OAI21x1_ASAP7_75t_L g543 ( .A1(n_222), .A2(n_544), .B(n_565), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_222), .B(n_547), .Y(n_568) );
INVx1_ASAP7_75t_L g697 ( .A(n_225), .Y(n_697) );
INVx1_ASAP7_75t_L g303 ( .A(n_227), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_227), .B(n_264), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_228), .B(n_411), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_232), .A2(n_258), .B1(n_323), .B2(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g699 ( .A(n_233), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_234), .A2(n_241), .B1(n_559), .B2(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g844 ( .A(n_237), .Y(n_844) );
INVx1_ASAP7_75t_L g708 ( .A(n_240), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_249), .A2(n_260), .B1(n_318), .B2(n_479), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_250), .B(n_355), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_251), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g538 ( .A(n_256), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_257), .A2(n_272), .B1(n_380), .B2(n_677), .Y(n_676) );
AOI22x1_ASAP7_75t_L g493 ( .A1(n_263), .A2(n_273), .B1(n_367), .B2(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_264), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g1020 ( .A(n_268), .Y(n_1020) );
AOI21xp33_ASAP7_75t_L g561 ( .A1(n_271), .A2(n_380), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g739 ( .A(n_274), .Y(n_739) );
HB1xp67_ASAP7_75t_L g1031 ( .A(n_274), .Y(n_1031) );
INVx1_ASAP7_75t_L g1021 ( .A(n_275), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_715), .B(n_723), .Y(n_282) );
XNOR2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_606), .Y(n_283) );
XOR2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_468), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_395), .B1(n_466), .B2(n_467), .Y(n_285) );
INVx1_ASAP7_75t_L g466 ( .A(n_286), .Y(n_466) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
XNOR2x1_ASAP7_75t_L g289 ( .A(n_290), .B(n_394), .Y(n_289) );
NAND4xp75_ASAP7_75t_L g290 ( .A(n_291), .B(n_332), .C(n_353), .D(n_365), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_322), .Y(n_291) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g979 ( .A(n_294), .Y(n_979) );
INVx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_295), .Y(n_454) );
BUFx12f_ASAP7_75t_L g479 ( .A(n_295), .Y(n_479) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_307), .Y(n_295) );
AND2x2_ASAP7_75t_L g319 ( .A(n_296), .B(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g324 ( .A(n_296), .B(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_L g329 ( .A(n_296), .B(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g417 ( .A(n_296), .B(n_325), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_296), .B(n_337), .Y(n_418) );
AND2x4_ASAP7_75t_L g423 ( .A(n_296), .B(n_307), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_296), .B(n_320), .Y(n_424) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_305), .Y(n_296) );
AND2x2_ASAP7_75t_L g361 ( .A(n_297), .B(n_306), .Y(n_361) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g336 ( .A(n_298), .B(n_306), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
NAND2xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g304 ( .A(n_300), .Y(n_304) );
INVx3_ASAP7_75t_L g310 ( .A(n_300), .Y(n_310) );
NAND2xp33_ASAP7_75t_L g316 ( .A(n_300), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g346 ( .A(n_300), .Y(n_346) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_300), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_301), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
OAI21xp5_ASAP7_75t_L g377 ( .A1(n_303), .A2(n_346), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g376 ( .A(n_306), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g368 ( .A(n_307), .B(n_336), .Y(n_368) );
AND2x4_ASAP7_75t_L g381 ( .A(n_307), .B(n_361), .Y(n_381) );
AND2x4_ASAP7_75t_L g403 ( .A(n_307), .B(n_361), .Y(n_403) );
AND2x4_ASAP7_75t_L g406 ( .A(n_307), .B(n_336), .Y(n_406) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_312), .Y(n_307) );
INVx2_ASAP7_75t_L g321 ( .A(n_308), .Y(n_321) );
AND2x4_ASAP7_75t_L g325 ( .A(n_308), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g331 ( .A(n_308), .B(n_327), .Y(n_331) );
AND2x2_ASAP7_75t_L g372 ( .A(n_308), .B(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_310), .B(n_315), .Y(n_314) );
INVxp67_ASAP7_75t_L g342 ( .A(n_310), .Y(n_342) );
NAND3xp33_ASAP7_75t_L g392 ( .A(n_311), .B(n_341), .C(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g320 ( .A(n_312), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g327 ( .A(n_313), .Y(n_327) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
BUFx2_ASAP7_75t_SL g1007 ( .A(n_318), .Y(n_1007) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx5_ASAP7_75t_L g455 ( .A(n_319), .Y(n_455) );
INVx1_ASAP7_75t_L g598 ( .A(n_319), .Y(n_598) );
BUFx3_ASAP7_75t_L g624 ( .A(n_319), .Y(n_624) );
AND2x2_ASAP7_75t_L g357 ( .A(n_320), .B(n_336), .Y(n_357) );
AND2x4_ASAP7_75t_L g360 ( .A(n_320), .B(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g364 ( .A(n_320), .B(n_340), .Y(n_364) );
AND2x4_ASAP7_75t_L g407 ( .A(n_320), .B(n_340), .Y(n_407) );
AND2x2_ASAP7_75t_L g409 ( .A(n_320), .B(n_361), .Y(n_409) );
AND2x2_ASAP7_75t_L g411 ( .A(n_320), .B(n_336), .Y(n_411) );
BUFx12f_ASAP7_75t_L g593 ( .A(n_323), .Y(n_593) );
INVx1_ASAP7_75t_L g975 ( .A(n_323), .Y(n_975) );
BUFx6f_ASAP7_75t_L g1011 ( .A(n_323), .Y(n_1011) );
BUFx12f_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_324), .Y(n_457) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_324), .Y(n_481) );
AND2x2_ASAP7_75t_L g349 ( .A(n_325), .B(n_336), .Y(n_349) );
AND2x4_ASAP7_75t_L g352 ( .A(n_325), .B(n_340), .Y(n_352) );
AND2x4_ASAP7_75t_L g420 ( .A(n_325), .B(n_336), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_325), .B(n_340), .Y(n_421) );
AND2x2_ASAP7_75t_L g524 ( .A(n_325), .B(n_336), .Y(n_524) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_325), .Y(n_628) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_329), .Y(n_440) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_329), .Y(n_527) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_329), .Y(n_626) );
AND2x4_ASAP7_75t_L g339 ( .A(n_330), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g414 ( .A(n_330), .B(n_336), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_330), .B(n_340), .Y(n_415) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g337 ( .A(n_331), .Y(n_337) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_347), .Y(n_332) );
BUFx12f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_335), .Y(n_445) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_335), .Y(n_520) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_335), .Y(n_549) );
BUFx3_ASAP7_75t_L g957 ( .A(n_335), .Y(n_957) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
BUFx3_ASAP7_75t_L g1004 ( .A(n_338), .Y(n_1004) );
BUFx12f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx6_ASAP7_75t_L g442 ( .A(n_339), .Y(n_442) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_345), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx8_ASAP7_75t_L g444 ( .A(n_349), .Y(n_444) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx4_ASAP7_75t_L g458 ( .A(n_351), .Y(n_458) );
INVx4_ASAP7_75t_L g525 ( .A(n_351), .Y(n_525) );
INVx4_ASAP7_75t_L g600 ( .A(n_351), .Y(n_600) );
INVx1_ASAP7_75t_L g961 ( .A(n_351), .Y(n_961) );
INVx8_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_358), .Y(n_353) );
INVx3_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g532 ( .A(n_356), .Y(n_532) );
INVx2_ASAP7_75t_L g681 ( .A(n_356), .Y(n_681) );
INVx2_ASAP7_75t_L g710 ( .A(n_356), .Y(n_710) );
INVx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx3_ASAP7_75t_L g432 ( .A(n_357), .Y(n_432) );
INVx2_ASAP7_75t_L g575 ( .A(n_357), .Y(n_575) );
BUFx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_360), .Y(n_491) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_360), .Y(n_557) );
INVx2_ASAP7_75t_L g583 ( .A(n_360), .Y(n_583) );
BUFx8_ASAP7_75t_SL g656 ( .A(n_360), .Y(n_656) );
INVx2_ASAP7_75t_L g704 ( .A(n_360), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_362), .Y(n_706) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g492 ( .A(n_363), .Y(n_492) );
INVx2_ASAP7_75t_L g616 ( .A(n_363), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_363), .A2(n_965), .B1(n_1020), .B2(n_1021), .Y(n_1019) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_364), .Y(n_452) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_364), .Y(n_530) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_379), .Y(n_365) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g449 ( .A(n_368), .Y(n_449) );
INVx2_ASAP7_75t_L g590 ( .A(n_368), .Y(n_590) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g450 ( .A(n_370), .Y(n_450) );
INVx4_ASAP7_75t_L g494 ( .A(n_370), .Y(n_494) );
OAI21xp33_ASAP7_75t_L g576 ( .A1(n_370), .A2(n_577), .B(n_578), .Y(n_576) );
OAI21xp5_ASAP7_75t_L g682 ( .A1(n_370), .A2(n_683), .B(n_684), .Y(n_682) );
INVx5_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx4f_ASAP7_75t_L g559 ( .A(n_371), .Y(n_559) );
BUFx2_ASAP7_75t_L g618 ( .A(n_371), .Y(n_618) );
BUFx2_ASAP7_75t_L g633 ( .A(n_371), .Y(n_633) );
AND2x4_ASAP7_75t_L g371 ( .A(n_372), .B(n_376), .Y(n_371) );
AND2x2_ASAP7_75t_L g404 ( .A(n_372), .B(n_376), .Y(n_404) );
AND2x4_ASAP7_75t_L g506 ( .A(n_372), .B(n_376), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g388 ( .A(n_374), .Y(n_388) );
INVx4_ASAP7_75t_L g698 ( .A(n_380), .Y(n_698) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g486 ( .A(n_381), .Y(n_486) );
BUFx3_ASAP7_75t_L g535 ( .A(n_381), .Y(n_535) );
BUFx3_ASAP7_75t_L g615 ( .A(n_381), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_386), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_386), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_SL g712 ( .A(n_386), .Y(n_712) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx3_ASAP7_75t_L g436 ( .A(n_387), .Y(n_436) );
AO21x2_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B(n_392), .Y(n_387) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_389), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g467 ( .A(n_395), .Y(n_467) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
XNOR2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_425), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
XNOR2x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_412), .Y(n_400) );
NAND4xp25_ASAP7_75t_L g401 ( .A(n_402), .B(n_405), .C(n_408), .D(n_410), .Y(n_401) );
NAND4xp25_ASAP7_75t_L g412 ( .A(n_413), .B(n_416), .C(n_419), .D(n_422), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_426), .B(n_459), .Y(n_425) );
AOI21x1_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B(n_446), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_437), .Y(n_428) );
BUFx2_ASAP7_75t_L g460 ( .A(n_429), .Y(n_460) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g986 ( .A(n_432), .Y(n_986) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_435), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g658 ( .A(n_435), .Y(n_658) );
INVx4_ASAP7_75t_L g988 ( .A(n_435), .Y(n_988) );
INVx4_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx3_ASAP7_75t_L g580 ( .A(n_436), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_443), .Y(n_437) );
INVxp67_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g464 ( .A(n_439), .B(n_453), .Y(n_464) );
BUFx3_ASAP7_75t_L g1013 ( .A(n_440), .Y(n_1013) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx5_ASAP7_75t_L g550 ( .A(n_442), .Y(n_550) );
INVx2_ASAP7_75t_L g959 ( .A(n_442), .Y(n_959) );
INVx1_ASAP7_75t_L g465 ( .A(n_443), .Y(n_465) );
INVx1_ASAP7_75t_L g463 ( .A(n_447), .Y(n_463) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
NAND4xp75_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .C(n_464), .D(n_465), .Y(n_459) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
AO22x2_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_539), .B1(n_540), .B2(n_605), .Y(n_468) );
INVx2_ASAP7_75t_L g605 ( .A(n_469), .Y(n_605) );
XOR2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_513), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_496), .B2(n_512), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
XNOR2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_495), .Y(n_472) );
NOR3xp33_ASAP7_75t_SL g473 ( .A(n_474), .B(n_477), .C(n_482), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .C(n_490), .D(n_493), .Y(n_482) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_489), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g638 ( .A(n_489), .Y(n_638) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_504), .Y(n_498) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .C(n_502), .D(n_503), .Y(n_499) );
NAND4xp25_ASAP7_75t_L g504 ( .A(n_505), .B(n_507), .C(n_508), .D(n_509), .Y(n_504) );
BUFx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
XNOR2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
NOR4xp75_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .C(n_528), .D(n_533), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_526), .Y(n_521) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx4f_ASAP7_75t_L g643 ( .A(n_524), .Y(n_643) );
BUFx2_ASAP7_75t_L g1001 ( .A(n_525), .Y(n_1001) );
BUFx3_ASAP7_75t_L g976 ( .A(n_527), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx3_ASAP7_75t_L g967 ( .A(n_530), .Y(n_967) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_534), .B(n_536), .Y(n_533) );
INVx2_ASAP7_75t_L g586 ( .A(n_535), .Y(n_586) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_569), .B1(n_603), .B2(n_604), .Y(n_540) );
INVx1_ASAP7_75t_L g604 ( .A(n_541), .Y(n_604) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_554), .Y(n_544) );
NOR3xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .C(n_551), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NOR3xp33_ASAP7_75t_L g567 ( .A(n_548), .B(n_560), .C(n_568), .Y(n_567) );
BUFx3_ASAP7_75t_L g1003 ( .A(n_549), .Y(n_1003) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_551), .B(n_555), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_560), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
INVx2_ASAP7_75t_L g965 ( .A(n_557), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx2_ASAP7_75t_L g602 ( .A(n_570), .Y(n_602) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_591), .Y(n_570) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_581), .C(n_584), .Y(n_571) );
BUFx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_575), .Y(n_651) );
INVx4_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g635 ( .A(n_583), .Y(n_635) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_590), .Y(n_654) );
INVx1_ASAP7_75t_L g701 ( .A(n_590), .Y(n_701) );
NAND4xp25_ASAP7_75t_SL g591 ( .A(n_592), .B(n_594), .C(n_595), .D(n_599), .Y(n_591) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_666), .B1(n_667), .B2(n_713), .Y(n_606) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_646), .B(n_664), .Y(n_608) );
OA21x2_ASAP7_75t_L g714 ( .A1(n_609), .A2(n_646), .B(n_664), .Y(n_714) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g665 ( .A(n_610), .Y(n_665) );
XNOR2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_629), .Y(n_610) );
NOR2x1_ASAP7_75t_L g612 ( .A(n_613), .B(n_621), .Y(n_612) );
NAND4xp25_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .C(n_619), .D(n_620), .Y(n_613) );
NAND4xp25_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .C(n_625), .D(n_627), .Y(n_621) );
BUFx2_ASAP7_75t_L g980 ( .A(n_624), .Y(n_980) );
XOR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_645), .Y(n_629) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_631), .B(n_639), .Y(n_630) );
NAND4xp25_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .C(n_636), .D(n_637), .Y(n_631) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .C(n_642), .D(n_644), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_646), .B(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_659), .Y(n_647) );
NAND4xp25_ASAP7_75t_L g648 ( .A(n_649), .B(n_652), .C(n_655), .D(n_657), .Y(n_648) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g677 ( .A(n_654), .Y(n_677) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_654), .Y(n_971) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .C(n_662), .D(n_663), .Y(n_659) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
XOR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_687), .Y(n_667) );
XOR2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_686), .Y(n_668) );
NOR2x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_675), .Y(n_669) );
NAND4xp25_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .C(n_673), .D(n_674), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .C(n_685), .Y(n_675) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
XNOR2x1_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g843 ( .A1(n_688), .A2(n_755), .B1(n_757), .B2(n_844), .C(n_845), .Y(n_843) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_695), .Y(n_689) );
AND4x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .C(n_693), .D(n_694), .Y(n_690) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_702), .C(n_707), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B1(n_699), .B2(n_700), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g968 ( .A1(n_698), .A2(n_969), .B1(n_970), .B2(n_971), .Y(n_968) );
OAI22xp5_ASAP7_75t_SL g1016 ( .A1(n_698), .A2(n_971), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_702) );
OAI21xp33_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_709), .B(n_711), .Y(n_707) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
BUFx4_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
NAND3xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_721), .C(n_722), .Y(n_717) );
AND2x2_ASAP7_75t_L g990 ( .A(n_718), .B(n_991), .Y(n_990) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_718), .B(n_992), .Y(n_1027) );
AOI21xp5_ASAP7_75t_L g1032 ( .A1(n_718), .A2(n_722), .B(n_768), .Y(n_1032) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AO21x1_ASAP7_75t_L g1029 ( .A1(n_719), .A2(n_1030), .B(n_1032), .Y(n_1029) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g731 ( .A(n_720), .B(n_732), .Y(n_731) );
AND3x4_ASAP7_75t_L g767 ( .A(n_720), .B(n_738), .C(n_768), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g991 ( .A(n_721), .B(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_722), .Y(n_992) );
OAI221xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_949), .B1(n_951), .B2(n_989), .C(n_993), .Y(n_723) );
O2A1O1Ixp33_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_816), .B(n_841), .C(n_846), .Y(n_724) );
OAI211xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_750), .B(n_780), .C(n_799), .Y(n_725) );
INVx1_ASAP7_75t_L g900 ( .A(n_726), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_743), .Y(n_726) );
AND2x2_ASAP7_75t_L g797 ( .A(n_727), .B(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g827 ( .A(n_727), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_727), .B(n_842), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_727), .B(n_842), .Y(n_926) );
NOR3xp33_ASAP7_75t_L g945 ( .A(n_727), .B(n_832), .C(n_946), .Y(n_945) );
INVx3_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OR2x2_ASAP7_75t_L g810 ( .A(n_728), .B(n_743), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_728), .B(n_803), .Y(n_870) );
AND2x2_ASAP7_75t_L g906 ( .A(n_728), .B(n_907), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_728), .B(n_743), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_728), .B(n_835), .Y(n_932) );
AND2x2_ASAP7_75t_L g943 ( .A(n_728), .B(n_744), .Y(n_943) );
AND2x4_ASAP7_75t_L g728 ( .A(n_729), .B(n_736), .Y(n_728) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
AND2x4_ASAP7_75t_L g737 ( .A(n_731), .B(n_738), .Y(n_737) );
AND2x4_ASAP7_75t_L g746 ( .A(n_731), .B(n_733), .Y(n_746) );
AND2x2_ASAP7_75t_L g770 ( .A(n_731), .B(n_733), .Y(n_770) );
AND2x4_ASAP7_75t_L g734 ( .A(n_733), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g747 ( .A(n_733), .B(n_735), .Y(n_747) );
AND2x2_ASAP7_75t_L g771 ( .A(n_733), .B(n_735), .Y(n_771) );
INVx2_ASAP7_75t_L g763 ( .A(n_734), .Y(n_763) );
AND2x4_ASAP7_75t_L g742 ( .A(n_735), .B(n_738), .Y(n_742) );
AND2x4_ASAP7_75t_L g749 ( .A(n_735), .B(n_738), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_735), .B(n_738), .Y(n_757) );
INVx3_ASAP7_75t_L g755 ( .A(n_737), .Y(n_755) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx3_ASAP7_75t_L g824 ( .A(n_743), .Y(n_824) );
AND2x2_ASAP7_75t_L g828 ( .A(n_743), .B(n_753), .Y(n_828) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g835 ( .A(n_744), .B(n_753), .Y(n_835) );
AND2x2_ASAP7_75t_L g865 ( .A(n_744), .B(n_798), .Y(n_865) );
OR2x2_ASAP7_75t_L g875 ( .A(n_744), .B(n_753), .Y(n_875) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_748), .Y(n_744) );
INVx3_ASAP7_75t_L g761 ( .A(n_746), .Y(n_761) );
BUFx2_ASAP7_75t_L g950 ( .A(n_746), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_764), .Y(n_750) );
INVx2_ASAP7_75t_L g853 ( .A(n_751), .Y(n_853) );
O2A1O1Ixp33_ASAP7_75t_SL g910 ( .A1(n_751), .A2(n_782), .B(n_911), .C(n_913), .Y(n_910) );
BUFx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_752), .B(n_801), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_752), .B(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g860 ( .A(n_752), .Y(n_860) );
AND2x2_ASAP7_75t_L g893 ( .A(n_752), .B(n_871), .Y(n_893) );
O2A1O1Ixp33_ASAP7_75t_L g897 ( .A1(n_752), .A2(n_898), .B(n_899), .C(n_900), .Y(n_897) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx3_ASAP7_75t_L g798 ( .A(n_753), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_753), .B(n_787), .Y(n_840) );
OR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_759), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_757), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_759) );
AND2x2_ASAP7_75t_L g786 ( .A(n_764), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g863 ( .A(n_764), .Y(n_863) );
AND2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_772), .Y(n_764) );
CKINVDCx6p67_ASAP7_75t_R g783 ( .A(n_765), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_765), .B(n_777), .Y(n_801) );
INVx1_ASAP7_75t_L g808 ( .A(n_765), .Y(n_808) );
AND2x2_ASAP7_75t_L g820 ( .A(n_765), .B(n_821), .Y(n_820) );
OR2x2_ASAP7_75t_L g890 ( .A(n_765), .B(n_777), .Y(n_890) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_769), .Y(n_765) );
INVx1_ASAP7_75t_L g789 ( .A(n_767), .Y(n_789) );
INVx1_ASAP7_75t_L g796 ( .A(n_770), .Y(n_796) );
INVx1_ASAP7_75t_L g794 ( .A(n_771), .Y(n_794) );
AND2x2_ASAP7_75t_SL g916 ( .A(n_772), .B(n_783), .Y(n_916) );
AND2x2_ASAP7_75t_L g923 ( .A(n_772), .B(n_852), .Y(n_923) );
OR2x2_ASAP7_75t_L g929 ( .A(n_772), .B(n_821), .Y(n_929) );
INVxp33_ASAP7_75t_L g936 ( .A(n_772), .Y(n_936) );
AND2x2_ASAP7_75t_L g772 ( .A(n_773), .B(n_776), .Y(n_772) );
INVx1_ASAP7_75t_L g785 ( .A(n_773), .Y(n_785) );
AND2x2_ASAP7_75t_L g813 ( .A(n_773), .B(n_777), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
AND2x2_ASAP7_75t_L g784 ( .A(n_776), .B(n_785), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_776), .B(n_807), .Y(n_887) );
OAI222xp33_ASAP7_75t_L g920 ( .A1(n_776), .A2(n_904), .B1(n_909), .B2(n_921), .C1(n_922), .C2(n_924), .Y(n_920) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g821 ( .A(n_777), .B(n_785), .Y(n_821) );
AOI322xp5_ASAP7_75t_L g869 ( .A1(n_777), .A2(n_824), .A3(n_826), .B1(n_860), .B2(n_870), .C1(n_871), .C2(n_873), .Y(n_869) );
AND2x4_ASAP7_75t_SL g777 ( .A(n_778), .B(n_779), .Y(n_777) );
OAI21xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_786), .B(n_797), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
AND2x2_ASAP7_75t_L g814 ( .A(n_783), .B(n_815), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_783), .B(n_813), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_783), .B(n_787), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_783), .B(n_829), .Y(n_834) );
AND2x2_ASAP7_75t_L g856 ( .A(n_783), .B(n_785), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_783), .A2(n_862), .B1(n_863), .B2(n_864), .Y(n_861) );
AND2x2_ASAP7_75t_L g881 ( .A(n_783), .B(n_821), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_783), .B(n_859), .Y(n_901) );
AND2x2_ASAP7_75t_L g851 ( .A(n_784), .B(n_852), .Y(n_851) );
AND2x2_ASAP7_75t_L g859 ( .A(n_784), .B(n_787), .Y(n_859) );
INVx1_ASAP7_75t_L g874 ( .A(n_784), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_785), .B(n_807), .Y(n_806) );
AND2x2_ASAP7_75t_L g839 ( .A(n_785), .B(n_807), .Y(n_839) );
INVx1_ASAP7_75t_L g868 ( .A(n_785), .Y(n_868) );
INVx1_ASAP7_75t_L g804 ( .A(n_787), .Y(n_804) );
CKINVDCx6p67_ASAP7_75t_R g815 ( .A(n_787), .Y(n_815) );
AND2x2_ASAP7_75t_L g877 ( .A(n_787), .B(n_798), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_787), .B(n_806), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_787), .B(n_798), .Y(n_941) );
OR2x6_ASAP7_75t_SL g787 ( .A(n_788), .B(n_792), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_795), .B2(n_796), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_798), .B(n_810), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_798), .B(n_827), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_798), .B(n_912), .Y(n_911) );
NOR2xp33_ASAP7_75t_L g947 ( .A(n_798), .B(n_815), .Y(n_947) );
O2A1O1Ixp33_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_802), .B(n_809), .C(n_811), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_805), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_803), .B(n_820), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_803), .B(n_865), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g935 ( .A(n_803), .B(n_936), .Y(n_935) );
INVx3_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_L g852 ( .A(n_807), .B(n_815), .Y(n_852) );
AND2x2_ASAP7_75t_L g858 ( .A(n_807), .B(n_859), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_807), .B(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AOI221xp5_ASAP7_75t_L g892 ( .A1(n_809), .A2(n_842), .B1(n_893), .B2(n_894), .C(n_896), .Y(n_892) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g829 ( .A(n_813), .Y(n_829) );
AND2x2_ASAP7_75t_L g871 ( .A(n_813), .B(n_872), .Y(n_871) );
AND2x2_ASAP7_75t_L g912 ( .A(n_813), .B(n_852), .Y(n_912) );
INVxp67_ASAP7_75t_L g930 ( .A(n_814), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_815), .B(n_824), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_815), .B(n_835), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_815), .B(n_865), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_815), .B(n_881), .Y(n_880) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_815), .B(n_887), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_815), .B(n_875), .Y(n_891) );
OAI221xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_823), .B1(n_825), .B2(n_829), .C(n_830), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_822), .Y(n_818) );
OAI221xp5_ASAP7_75t_L g937 ( .A1(n_819), .A2(n_931), .B1(n_938), .B2(n_942), .C(n_944), .Y(n_937) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
OAI21xp33_ASAP7_75t_L g888 ( .A1(n_820), .A2(n_889), .B(n_891), .Y(n_888) );
INVx1_ASAP7_75t_L g832 ( .A(n_821), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_821), .B(n_877), .Y(n_876) );
OAI321xp33_ASAP7_75t_L g927 ( .A1(n_822), .A2(n_928), .A3(n_930), .B1(n_931), .B2(n_932), .C(n_933), .Y(n_927) );
INVx3_ASAP7_75t_L g837 ( .A(n_824), .Y(n_837) );
INVx1_ASAP7_75t_L g924 ( .A(n_824), .Y(n_924) );
O2A1O1Ixp33_ASAP7_75t_SL g866 ( .A1(n_825), .A2(n_867), .B(n_869), .C(n_878), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_826), .B(n_828), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g914 ( .A(n_826), .B(n_915), .Y(n_914) );
INVx3_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g862 ( .A(n_828), .Y(n_862) );
NAND3xp33_ASAP7_75t_L g933 ( .A(n_828), .B(n_839), .C(n_870), .Y(n_933) );
O2A1O1Ixp33_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_834), .B(n_835), .C(n_836), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
INVx1_ASAP7_75t_L g872 ( .A(n_833), .Y(n_872) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_834), .B(n_851), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_837), .B(n_878), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_837), .B(n_842), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
CKINVDCx16_ASAP7_75t_R g948 ( .A(n_841), .Y(n_948) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
BUFx3_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g878 ( .A(n_843), .Y(n_878) );
NAND5xp2_ASAP7_75t_L g846 ( .A(n_847), .B(n_892), .C(n_905), .D(n_917), .E(n_934), .Y(n_846) );
AOI211xp5_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .B(n_866), .C(n_879), .Y(n_847) );
OAI221xp5_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_853), .B1(n_854), .B2(n_855), .C(n_857), .Y(n_849) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
AOI21xp5_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_860), .B(n_861), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g894 ( .A(n_860), .B(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g904 ( .A(n_865), .Y(n_904) );
INVx1_ASAP7_75t_L g940 ( .A(n_868), .Y(n_940) );
OAI21xp33_ASAP7_75t_SL g873 ( .A1(n_874), .A2(n_875), .B(n_876), .Y(n_873) );
INVx1_ASAP7_75t_L g907 ( .A(n_875), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_877), .B(n_916), .Y(n_915) );
CKINVDCx16_ASAP7_75t_R g898 ( .A(n_878), .Y(n_898) );
NOR2xp33_ASAP7_75t_L g903 ( .A(n_878), .B(n_904), .Y(n_903) );
OAI221xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_882), .B1(n_883), .B2(n_885), .C(n_888), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_881), .B(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g918 ( .A(n_895), .Y(n_918) );
OAI21xp33_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_901), .B(n_902), .Y(n_896) );
AOI211xp5_ASAP7_75t_L g905 ( .A1(n_906), .A2(n_908), .B(n_910), .C(n_914), .Y(n_905) );
A2O1A1Ixp33_ASAP7_75t_L g934 ( .A1(n_906), .A2(n_935), .B(n_937), .C(n_948), .Y(n_934) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g919 ( .A(n_913), .Y(n_919) );
AOI221xp5_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_919), .B1(n_920), .B2(n_925), .C(n_927), .Y(n_917) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVxp67_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_939), .B(n_941), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
CKINVDCx5p33_ASAP7_75t_R g949 ( .A(n_950), .Y(n_949) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
NAND4xp75_ASAP7_75t_L g954 ( .A(n_955), .B(n_962), .C(n_972), .D(n_981), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_956), .B(n_960), .Y(n_955) );
BUFx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
NOR2x1_ASAP7_75t_L g962 ( .A(n_963), .B(n_968), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_964), .A2(n_965), .B1(n_966), .B2(n_967), .Y(n_963) );
AND2x2_ASAP7_75t_L g972 ( .A(n_973), .B(n_977), .Y(n_972) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
BUFx4f_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
OAI21xp33_ASAP7_75t_L g982 ( .A1(n_983), .A2(n_984), .B(n_987), .Y(n_982) );
OAI21xp33_ASAP7_75t_L g1022 ( .A1(n_984), .A2(n_1023), .B(n_1024), .Y(n_1022) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g1025 ( .A(n_996), .Y(n_1025) );
HB1xp67_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
NAND3xp33_ASAP7_75t_L g997 ( .A(n_998), .B(n_1005), .C(n_1015), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1002), .Y(n_999) );
NOR2x1_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1008), .Y(n_1005) );
OAI22x1_ASAP7_75t_SL g1008 ( .A1(n_1009), .A2(n_1010), .B1(n_1012), .B2(n_1014), .Y(n_1008) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
NOR3xp33_ASAP7_75t_SL g1015 ( .A(n_1016), .B(n_1019), .C(n_1022), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
BUFx3_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_1031), .Y(n_1030) );
endmodule