module real_jpeg_32337_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_586;
wire n_405;
wire n_412;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_0),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_0),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_0),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_1),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_1),
.B(n_147),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_1),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_1),
.B(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_1),
.B(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_1),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_2),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_2),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_2),
.B(n_337),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_2),
.B(n_348),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_2),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_2),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_2),
.B(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_2),
.B(n_531),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_3),
.B(n_82),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_3),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_3),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_3),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_3),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_3),
.B(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_SL g366 ( 
.A(n_3),
.B(n_367),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_4),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_5),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_5),
.Y(n_432)
);

NAND2x1_ASAP7_75t_SL g29 ( 
.A(n_6),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_6),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_6),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_6),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_6),
.B(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_6),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_6),
.B(n_178),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_6),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_7),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_7),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_7),
.B(n_416),
.Y(n_415)
);

AND2x4_ASAP7_75t_SL g437 ( 
.A(n_7),
.B(n_438),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_7),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_7),
.B(n_509),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_7),
.B(n_535),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_8),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_8),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_8),
.B(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_SL g347 ( 
.A(n_8),
.B(n_348),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_8),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_8),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_8),
.B(n_256),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_8),
.B(n_498),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_9),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_10),
.Y(n_184)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_11),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_11),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_11),
.Y(n_495)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_12),
.Y(n_119)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_12),
.Y(n_190)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_12),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_13),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_13),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_13),
.B(n_36),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_13),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_13),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_13),
.B(n_188),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_13),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_13),
.B(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_14),
.B(n_40),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_14),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_14),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_14),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_14),
.B(n_166),
.Y(n_165)
);

OAI222xp33_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_21),
.B1(n_133),
.B2(n_134),
.C1(n_588),
.C2(n_589),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_15),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_16),
.B(n_130),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_17),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_17),
.Y(n_180)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_17),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_18),
.B(n_92),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_18),
.B(n_170),
.Y(n_169)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_18),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_18),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_18),
.B(n_149),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_18),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_18),
.B(n_410),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_18),
.B(n_414),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_19),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_19),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_19),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_19),
.B(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_19),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_19),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_19),
.B(n_166),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_129),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_23),
.B(n_129),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_128),
.Y(n_23)
);

NAND2x1p5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_86),
.Y(n_24)
);

OR2x2_ASAP7_75t_SL g128 ( 
.A(n_25),
.B(n_86),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_60),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_44),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.C(n_38),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_28),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_31),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_33),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_32),
.A2(n_33),
.B1(n_38),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_37),
.Y(n_328)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_39),
.A2(n_76),
.B1(n_77),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_39),
.Y(n_123)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_42),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_43),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_43),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_52),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_51),
.Y(n_319)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_66),
.C(n_74),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_61),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_76),
.C(n_81),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_66),
.A2(n_74),
.B1(n_75),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_73),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_73),
.Y(n_254)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_76),
.A2(n_77),
.B1(n_116),
.B2(n_117),
.Y(n_280)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_111),
.C(n_116),
.Y(n_110)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_124),
.C(n_125),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_87),
.B(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_110),
.C(n_120),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_88),
.B(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_98),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_94),
.C(n_98),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_92),
.Y(n_210)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_97),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_106),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_99),
.A2(n_100),
.B1(n_106),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_103),
.B(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_106),
.Y(n_275)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_110),
.B(n_121),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_111),
.B(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g147 ( 
.A(n_115),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_116),
.B(n_201),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_116),
.B(n_201),
.C(n_216),
.Y(n_282)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_119),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_119),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_124),
.B(n_125),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_129),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx12f_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21x1_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_306),
.B(n_583),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_290),
.C(n_301),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_265),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_139),
.B(n_266),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_203),
.C(n_221),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_141),
.A2(n_142),
.B1(n_204),
.B2(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_173),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_158),
.B1(n_171),
.B2(n_172),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_144),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_153),
.C(n_156),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_153),
.C(n_156),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_145),
.B(n_245),
.Y(n_244)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_151),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_146),
.B(n_151),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_148),
.B(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_150),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_150),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_150),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_153),
.A2(n_156),
.B1(n_157),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_153),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_169),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_157),
.B(n_159),
.C(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_167),
.B2(n_168),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_165),
.Y(n_160)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_163),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_163),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_164),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_192),
.C(n_195),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_165),
.B(n_192),
.Y(n_242)
);

INVx8_ASAP7_75t_L g542 ( 
.A(n_166),
.Y(n_542)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_169),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_172),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_173),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_191),
.C(n_199),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_175),
.B(n_391),
.Y(n_390)
);

XNOR2x1_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_185),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_181),
.C(n_186),
.Y(n_206)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_183),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_184),
.Y(n_469)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_189),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_190),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_190),
.Y(n_528)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_191),
.Y(n_391)
);

BUFx4f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_194),
.Y(n_365)
);

XOR2x2_ASAP7_75t_L g241 ( 
.A(n_195),
.B(n_242),
.Y(n_241)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2x2_ASAP7_75t_SL g389 ( 
.A(n_199),
.B(n_390),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_204),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_215),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_206),
.B(n_207),
.C(n_215),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_208),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_212),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_213),
.B(n_284),
.C(n_285),
.Y(n_283)
);

XOR2x1_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_219),
.Y(n_417)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_222),
.B(n_397),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_243),
.C(n_247),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_223),
.A2(n_224),
.B1(n_393),
.B2(n_394),
.Y(n_392)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.C(n_241),
.Y(n_224)
);

XOR2x2_ASAP7_75t_L g354 ( 
.A(n_225),
.B(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_227),
.B(n_241),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.C(n_238),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_228),
.B(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_234),
.A2(n_238),
.B1(n_239),
.B2(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_234),
.Y(n_381)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_244),
.B(n_247),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_259),
.C(n_263),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_248),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.C(n_255),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_249),
.B(n_255),
.Y(n_334)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_252),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_252),
.Y(n_498)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_252),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_253),
.B(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g537 ( 
.A(n_258),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_259),
.B(n_263),
.Y(n_330)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_286),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_278),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_276),
.B2(n_277),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_276),
.C(n_294),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_286),
.C(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_282),
.C(n_283),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_291),
.A2(n_585),
.B(n_586),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_299),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_292),
.B(n_299),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_296),
.C(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

OA21x2_ASAP7_75t_SL g583 ( 
.A1(n_301),
.A2(n_584),
.B(n_587),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_302),
.B(n_304),
.Y(n_587)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_401),
.B(n_580),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_395),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_385),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_310),
.B(n_385),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_354),
.C(n_356),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2x1_ASAP7_75t_L g557 ( 
.A(n_312),
.B(n_354),
.Y(n_557)
);

XOR2x2_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_331),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_329),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_314),
.B(n_329),
.C(n_387),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_322),
.C(n_325),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_315),
.B(n_384),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.C(n_320),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_316),
.A2(n_317),
.B1(n_320),
.B2(n_321),
.Y(n_422)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_318),
.B(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_321),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_322),
.B(n_325),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_324),
.Y(n_377)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_331),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.C(n_340),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_333),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_335),
.A2(n_336),
.B(n_339),
.Y(n_420)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_335),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_340),
.A2(n_568),
.B(n_569),
.Y(n_567)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_341),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_347),
.C(n_351),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_342),
.A2(n_343),
.B1(n_351),
.B2(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx4_ASAP7_75t_SL g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_351),
.Y(n_360)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2x1_ASAP7_75t_L g556 ( 
.A(n_356),
.B(n_557),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_378),
.C(n_382),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_357),
.B(n_561),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.C(n_370),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_358),
.B(n_442),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_361),
.B(n_370),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_366),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_362),
.A2(n_363),
.B1(n_366),
.B2(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_366),
.Y(n_440)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

MAJx2_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.C(n_375),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_371),
.B(n_375),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_372),
.B(n_426),
.Y(n_425)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_374),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_377),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_379),
.A2(n_382),
.B1(n_383),
.B2(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_379),
.Y(n_562)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_388),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_389),
.C(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_392),
.Y(n_400)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_393),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_395),
.A2(n_581),
.B(n_582),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_399),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_396),
.B(n_399),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_555),
.B(n_578),
.Y(n_401)
);

AO21x1_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_458),
.B(n_554),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_443),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_404),
.B(n_443),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_423),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_405),
.B(n_424),
.C(n_574),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_419),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_406),
.B(n_420),
.C(n_421),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_415),
.C(n_418),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_407),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_412),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_408),
.A2(n_409),
.B1(n_412),
.B2(n_413),
.Y(n_450)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_415),
.B(n_418),
.Y(n_448)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_441),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_427),
.C(n_439),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_425),
.B(n_446),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_427),
.B(n_439),
.Y(n_446)
);

MAJx2_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_433),
.C(n_437),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_428),
.A2(n_429),
.B1(n_437),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx8_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_433),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_436),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g480 ( 
.A(n_437),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_441),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_447),
.C(n_449),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_444),
.A2(n_445),
.B1(n_483),
.B2(n_484),
.Y(n_482)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_447),
.B(n_449),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.C(n_454),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_451),
.Y(n_462)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

XOR2x2_ASAP7_75t_SL g461 ( 
.A(n_454),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_457),
.Y(n_454)
);

AO22x1_ASAP7_75t_SL g499 ( 
.A1(n_455),
.A2(n_456),
.B1(n_457),
.B2(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_457),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_485),
.B(n_553),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_482),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_460),
.B(n_482),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_463),
.C(n_478),
.Y(n_460)
);

XNOR2x1_ASAP7_75t_L g501 ( 
.A(n_461),
.B(n_502),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_463),
.B(n_478),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_470),
.C(n_474),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_464),
.A2(n_465),
.B1(n_474),
.B2(n_475),
.Y(n_489)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_470),
.B(n_489),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_472),
.Y(n_470)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_481),
.Y(n_478)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_503),
.B(n_552),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_501),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_SL g552 ( 
.A(n_487),
.B(n_501),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_490),
.C(n_499),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_488),
.B(n_516),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_490),
.A2(n_491),
.B1(n_499),
.B2(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_496),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_492),
.A2(n_493),
.B1(n_496),
.B2(n_497),
.Y(n_507)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_499),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_518),
.B(n_551),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_515),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_505),
.B(n_515),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_508),
.C(n_511),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_506),
.A2(n_507),
.B1(n_548),
.B2(n_549),
.Y(n_547)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_508),
.B(n_511),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_513),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

OA21x2_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_544),
.B(n_550),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_521),
.A2(n_539),
.B(n_543),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_529),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_529),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_524),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_523),
.B(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_530),
.A2(n_533),
.B1(n_534),
.B2(n_538),
.Y(n_529)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_530),
.Y(n_538)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_533),
.B(n_540),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_538),
.Y(n_546)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_536),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_547),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_546),
.B(n_547),
.Y(n_550)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_548),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_556),
.A2(n_558),
.B(n_572),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_556),
.B(n_558),
.C(n_579),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_563),
.C(n_565),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_559),
.A2(n_560),
.B1(n_576),
.B2(n_577),
.Y(n_575)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_564),
.B(n_566),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

XNOR2x1_ASAP7_75t_L g566 ( 
.A(n_567),
.B(n_571),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_570),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_573),
.B(n_575),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_573),
.B(n_575),
.Y(n_579)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);


endmodule