module fake_jpeg_26781_n_174 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_SL g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_29),
.B(n_31),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_15),
.B(n_1),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx6p67_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_13),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_43),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_14),
.B1(n_22),
.B2(n_17),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_19),
.B1(n_29),
.B2(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_53),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_19),
.B1(n_21),
.B2(n_25),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_38),
.B1(n_21),
.B2(n_22),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_18),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_24),
.B1(n_18),
.B2(n_16),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_38),
.B1(n_33),
.B2(n_28),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_69),
.Y(n_83)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_29),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_28),
.Y(n_84)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_70),
.B1(n_45),
.B2(n_54),
.Y(n_71)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_35),
.B1(n_37),
.B2(n_34),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_68),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_36),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_37),
.B1(n_34),
.B2(n_33),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_41),
.B1(n_44),
.B2(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_76),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_40),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_47),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_84),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_85),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_30),
.Y(n_82)
);

OAI21x1_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_32),
.B(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_55),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_60),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_70),
.B1(n_68),
.B2(n_62),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_89),
.A2(n_102),
.B1(n_88),
.B2(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_93),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_46),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_98),
.Y(n_105)
);

OA21x2_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_85),
.B(n_74),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_46),
.B1(n_49),
.B2(n_40),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_17),
.B(n_32),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_83),
.B(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_102),
.B(n_103),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_116),
.B(n_94),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_84),
.C(n_77),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_101),
.C(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_74),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_118),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_71),
.B1(n_73),
.B2(n_18),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_89),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_123),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_103),
.B1(n_100),
.B2(n_88),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_110),
.B1(n_116),
.B2(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_132),
.C(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_116),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_129),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_94),
.C(n_73),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_126),
.B1(n_122),
.B2(n_112),
.C(n_124),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_131),
.B(n_65),
.Y(n_137)
);

OAI21x1_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_23),
.B(n_26),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_128),
.B(n_108),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_32),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_142),
.B(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_137),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_110),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_138),
.B(n_141),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_143),
.B1(n_125),
.B2(n_44),
.Y(n_147)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_120),
.B1(n_113),
.B2(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_145),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g145 ( 
.A(n_135),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_146),
.A2(n_150),
.B1(n_151),
.B2(n_145),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_148),
.C(n_149),
.Y(n_155)
);

AOI31xp33_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_134),
.A3(n_26),
.B(n_23),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_57),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_158),
.B1(n_44),
.B2(n_16),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_148),
.C(n_151),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_157),
.C(n_159),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_57),
.C(n_59),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_10),
.B1(n_12),
.B2(n_11),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_78),
.C(n_44),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_11),
.B(n_10),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_1),
.B(n_2),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_2),
.B(n_4),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_24),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_164),
.B(n_78),
.Y(n_169)
);

OAI221xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_78),
.B1(n_16),
.B2(n_4),
.C(n_5),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_163),
.A2(n_2),
.B(n_3),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_169),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_165),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_173),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_168),
.C(n_24),
.Y(n_173)
);


endmodule