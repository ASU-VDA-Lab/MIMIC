module real_jpeg_515_n_17 (n_108, n_8, n_0, n_111, n_2, n_10, n_9, n_12, n_107, n_6, n_104, n_106, n_11, n_14, n_110, n_112, n_7, n_3, n_5, n_4, n_102, n_105, n_109, n_1, n_16, n_15, n_13, n_103, n_17);

input n_108;
input n_8;
input n_0;
input n_111;
input n_2;
input n_10;
input n_9;
input n_12;
input n_107;
input n_6;
input n_104;
input n_106;
input n_11;
input n_14;
input n_110;
input n_112;
input n_7;
input n_3;
input n_5;
input n_4;
input n_102;
input n_105;
input n_109;
input n_1;
input n_16;
input n_15;
input n_13;
input n_103;

output n_17;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_37),
.C(n_61),
.Y(n_36)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_2),
.A2(n_35),
.B1(n_69),
.B2(n_72),
.Y(n_34)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_3),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_5),
.B(n_29),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_7),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_19)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_8),
.B(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_9),
.A2(n_44),
.B(n_48),
.Y(n_43)
);

AO22x1_ASAP7_75t_L g39 ( 
.A1(n_10),
.A2(n_40),
.B1(n_42),
.B2(n_53),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_39),
.C(n_54),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_12),
.Y(n_83)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_16),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_16),
.Y(n_96)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_26),
.B1(n_99),
.B2(n_100),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_23),
.B(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_24),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_26),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI221xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_34),
.B2(n_75),
.C(n_89),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_30),
.B(n_88),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_41),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_65),
.C(n_66),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_57),
.C(n_58),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_51),
.C(n_52),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_47),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_83),
.Y(n_82)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_84),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_90),
.A3(n_91),
.B1(n_94),
.B2(n_95),
.C1(n_98),
.C2(n_112),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.C(n_81),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_102),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_103),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_104),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_105),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_106),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_107),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_108),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_109),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_110),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_111),
.Y(n_88)
);


endmodule