module fake_jpeg_20027_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

AND2x4_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_49),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_21),
.B1(n_26),
.B2(n_15),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_51),
.B1(n_45),
.B2(n_50),
.Y(n_68)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx2_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_53),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_26),
.B1(n_30),
.B2(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_32),
.B1(n_38),
.B2(n_34),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_58),
.A2(n_78),
.B1(n_63),
.B2(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_77),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_32),
.B1(n_36),
.B2(n_31),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_52),
.B1(n_53),
.B2(n_46),
.Y(n_93)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_31),
.B1(n_27),
.B2(n_30),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_17),
.B1(n_25),
.B2(n_28),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_68),
.Y(n_108)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_27),
.B1(n_29),
.B2(n_25),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_80),
.B1(n_51),
.B2(n_50),
.Y(n_89)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_71),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

AO22x2_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_34),
.B1(n_33),
.B2(n_23),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_52),
.A3(n_16),
.B1(n_20),
.B2(n_19),
.Y(n_107)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_40),
.A2(n_34),
.B1(n_28),
.B2(n_19),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_43),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_85),
.B(n_88),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_40),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_93),
.B1(n_98),
.B2(n_111),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_53),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_100),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_52),
.B1(n_42),
.B2(n_46),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_42),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_42),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_55),
.B1(n_56),
.B2(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_67),
.B(n_18),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_75),
.B1(n_78),
.B2(n_80),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_112),
.A2(n_117),
.B1(n_120),
.B2(n_124),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_126),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_75),
.B(n_60),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_114),
.B(n_139),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_119),
.B1(n_121),
.B2(n_113),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_108),
.A2(n_73),
.B1(n_62),
.B2(n_69),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

AO21x2_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_73),
.B(n_79),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_65),
.B1(n_18),
.B2(n_24),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_57),
.B(n_16),
.C(n_20),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_16),
.B(n_20),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_90),
.B(n_99),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_24),
.B1(n_57),
.B2(n_22),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_129),
.B1(n_130),
.B2(n_137),
.Y(n_141)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_83),
.B1(n_22),
.B2(n_16),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_92),
.B1(n_97),
.B2(n_103),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_22),
.B1(n_16),
.B2(n_5),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_110),
.B1(n_84),
.B2(n_92),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_137)
);

NAND2x1_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_3),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_88),
.C(n_85),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_153),
.C(n_155),
.Y(n_193)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_134),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g173 ( 
.A(n_143),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_146),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_115),
.A2(n_91),
.B1(n_87),
.B2(n_98),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_154),
.B1(n_158),
.B2(n_124),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_87),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_147),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_95),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_150),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_103),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_162),
.B(n_121),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_139),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_97),
.B1(n_92),
.B2(n_106),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_97),
.C(n_106),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_109),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_159),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_137),
.A2(n_92),
.B1(n_105),
.B2(n_90),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_109),
.B1(n_99),
.B2(n_5),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_3),
.Y(n_164)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_109),
.C(n_6),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_166),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_4),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_6),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_167),
.B(n_170),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_119),
.B(n_125),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_198),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

INVxp33_ASAP7_75t_SL g202 ( 
.A(n_175),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_121),
.B(n_119),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_179),
.B(n_171),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_196),
.B1(n_141),
.B2(n_152),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_179),
.A2(n_182),
.B(n_187),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_168),
.A2(n_129),
.B1(n_117),
.B2(n_120),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_185),
.B1(n_189),
.B2(n_190),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_125),
.B(n_119),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_119),
.B1(n_118),
.B2(n_134),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_184),
.A2(n_165),
.B1(n_158),
.B2(n_150),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_168),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

NAND2xp33_ASAP7_75t_R g187 ( 
.A(n_162),
.B(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_151),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_151),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_152),
.Y(n_191)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_151),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_141),
.B1(n_153),
.B2(n_13),
.Y(n_210)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_140),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_195),
.B(n_164),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_204),
.B(n_211),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_207),
.B1(n_185),
.B2(n_200),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_214),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_212),
.B1(n_216),
.B2(n_171),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_148),
.B1(n_157),
.B2(n_144),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_192),
.B1(n_190),
.B2(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_217),
.B(n_220),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_166),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_219),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_12),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_186),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_225),
.A2(n_214),
.B1(n_201),
.B2(n_217),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_183),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_234),
.B1(n_235),
.B2(n_238),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_212),
.B(n_183),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_215),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_198),
.B1(n_176),
.B2(n_180),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_236),
.B1(n_172),
.B2(n_201),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_209),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_205),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_205),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_178),
.B1(n_184),
.B2(n_180),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_240),
.A2(n_210),
.B1(n_203),
.B2(n_216),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_254),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_246),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_240),
.A2(n_203),
.B1(n_182),
.B2(n_194),
.Y(n_243)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_219),
.C(n_177),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_248),
.C(n_191),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_213),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_250),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_227),
.C(n_239),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_194),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_252),
.A2(n_255),
.B1(n_229),
.B2(n_224),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_226),
.B1(n_236),
.B2(n_223),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_258),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_255),
.A2(n_237),
.B1(n_228),
.B2(n_221),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_237),
.B1(n_208),
.B2(n_188),
.Y(n_259)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_261),
.B(n_262),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_191),
.B(n_12),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_242),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_12),
.C(n_13),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_253),
.C(n_244),
.Y(n_273)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_247),
.C(n_246),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_272),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_264),
.Y(n_272)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_273),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_267),
.B(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_276),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_241),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_257),
.Y(n_281)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_281),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_260),
.C(n_265),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_262),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_257),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_284),
.B(n_272),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_290),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_SL g292 ( 
.A(n_288),
.B(n_289),
.C(n_279),
.Y(n_292)
);

NOR2xp67_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_268),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_293),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_288),
.B(n_284),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_291),
.A2(n_285),
.B(n_278),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_283),
.B(n_287),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_295),
.C(n_275),
.Y(n_297)
);

A2O1A1O1Ixp25_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_261),
.B(n_269),
.C(n_266),
.D(n_13),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_298),
.B(n_13),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_266),
.Y(n_300)
);


endmodule