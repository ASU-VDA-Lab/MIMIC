module fake_jpeg_688_n_431 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_431);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_431;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_57),
.B(n_68),
.Y(n_114)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_60),
.Y(n_162)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_17),
.B(n_16),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_17),
.B(n_15),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_84),
.Y(n_127)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_53),
.Y(n_81)
);

INVx5_ASAP7_75t_SL g132 ( 
.A(n_81),
.Y(n_132)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_37),
.B(n_12),
.Y(n_84)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_88),
.Y(n_172)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_91),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_93),
.A2(n_26),
.B(n_53),
.Y(n_170)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_37),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_100),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_98),
.A2(n_25),
.B1(n_44),
.B2(n_47),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_0),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_50),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_35),
.B(n_0),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_11),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_104),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_1),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_23),
.B(n_43),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_111),
.Y(n_169)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_108),
.Y(n_176)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_22),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_109),
.B(n_24),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_120),
.B(n_171),
.C(n_5),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_22),
.B1(n_45),
.B2(n_40),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_122),
.A2(n_135),
.B1(n_141),
.B2(n_151),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_41),
.B1(n_45),
.B2(n_40),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_123),
.A2(n_173),
.B1(n_176),
.B2(n_137),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_65),
.A2(n_40),
.B1(n_45),
.B2(n_48),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_136),
.B(n_139),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_64),
.B(n_51),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_74),
.B1(n_92),
.B2(n_78),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_96),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_164),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_97),
.A2(n_22),
.B1(n_43),
.B2(n_50),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_102),
.A2(n_25),
.B1(n_23),
.B2(n_47),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_155),
.B1(n_168),
.B2(n_174),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_165),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_109),
.A2(n_24),
.B1(n_52),
.B2(n_36),
.Y(n_155)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_69),
.B(n_46),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_60),
.B(n_46),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_178),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_54),
.A2(n_52),
.B1(n_36),
.B2(n_28),
.Y(n_168)
);

OR2x2_ASAP7_75t_SL g210 ( 
.A(n_170),
.B(n_123),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_60),
.B(n_28),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_91),
.A2(n_44),
.B1(n_53),
.B2(n_5),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_85),
.A2(n_103),
.B1(n_110),
.B2(n_77),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_55),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_59),
.B(n_10),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_116),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_181),
.B(n_190),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g275 ( 
.A1(n_182),
.A2(n_191),
.B1(n_204),
.B2(n_209),
.Y(n_275)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_150),
.B(n_3),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_185),
.B(n_201),
.Y(n_266)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_187),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_189),
.A2(n_219),
.B1(n_236),
.B2(n_229),
.Y(n_253)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_191),
.Y(n_277)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_197),
.Y(n_250)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_199),
.Y(n_274)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_114),
.B(n_6),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_7),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_208),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_117),
.B(n_156),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_203),
.B(n_205),
.Y(n_243)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_113),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_130),
.B(n_140),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_146),
.B(n_132),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_206),
.B(n_211),
.Y(n_278)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_134),
.Y(n_207)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_127),
.B(n_167),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_142),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_209),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_210),
.B(n_232),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_132),
.B(n_115),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_212),
.B(n_213),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_121),
.B(n_160),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_147),
.B(n_172),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_214),
.B(n_215),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_119),
.B(n_148),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_152),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_216),
.B(n_218),
.Y(n_269)
);

BUFx12_ASAP7_75t_L g217 ( 
.A(n_142),
.Y(n_217)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_119),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_122),
.A2(n_135),
.B1(n_143),
.B2(n_159),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_131),
.A2(n_124),
.B1(n_152),
.B2(n_128),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_220),
.Y(n_263)
);

AOI32xp33_ASAP7_75t_L g221 ( 
.A1(n_129),
.A2(n_133),
.A3(n_137),
.B1(n_173),
.B2(n_175),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_221),
.B(n_224),
.Y(n_279)
);

OR2x2_ASAP7_75t_SL g222 ( 
.A(n_142),
.B(n_175),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_227),
.Y(n_241)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_138),
.Y(n_223)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_118),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_118),
.A2(n_149),
.B1(n_138),
.B2(n_143),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_145),
.B(n_159),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_230),
.Y(n_265)
);

OR2x2_ASAP7_75t_SL g227 ( 
.A(n_125),
.B(n_158),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_125),
.A2(n_157),
.B(n_180),
.C(n_161),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_218),
.B(n_211),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_180),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_157),
.Y(n_232)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_149),
.Y(n_233)
);

CKINVDCx12_ASAP7_75t_R g260 ( 
.A(n_233),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_161),
.B(n_163),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_235),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_151),
.A2(n_141),
.B1(n_153),
.B2(n_83),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_134),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_238),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_152),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_208),
.C(n_199),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_244),
.B(n_264),
.C(n_217),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_251),
.A2(n_253),
.B1(n_237),
.B2(n_223),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_206),
.B(n_227),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_252),
.A2(n_276),
.B(n_246),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_184),
.A2(n_196),
.B1(n_183),
.B2(n_229),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_255),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_215),
.A2(n_214),
.B1(n_202),
.B2(n_226),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_198),
.A2(n_192),
.B1(n_188),
.B2(n_235),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_198),
.A2(n_230),
.B1(n_200),
.B2(n_216),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_195),
.B(n_198),
.C(n_181),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_222),
.A2(n_186),
.B(n_238),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_187),
.A2(n_197),
.B(n_231),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_281),
.A2(n_263),
.B(n_282),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_194),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_283),
.B(n_295),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_278),
.B(n_231),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_284),
.B(n_303),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_264),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_285),
.B(n_307),
.Y(n_337)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_286),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_287),
.B(n_292),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_249),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_289),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_265),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_290),
.A2(n_248),
.B1(n_240),
.B2(n_260),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_244),
.B(n_217),
.C(n_207),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_253),
.A2(n_233),
.B1(n_252),
.B2(n_251),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_294),
.A2(n_304),
.B1(n_313),
.B2(n_240),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_242),
.B(n_262),
.Y(n_295)
);

A2O1A1O1Ixp25_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_278),
.B(n_279),
.C(n_269),
.D(n_262),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_296),
.A2(n_308),
.B(n_309),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_310),
.Y(n_331)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_298),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_241),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_300),
.B(n_306),
.Y(n_340)
);

XNOR2x1_ASAP7_75t_SL g301 ( 
.A(n_271),
.B(n_241),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_302),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_276),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_266),
.B(n_239),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_241),
.A2(n_256),
.B1(n_245),
.B2(n_272),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_254),
.B(n_275),
.C(n_277),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_250),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_254),
.B(n_280),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_239),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_280),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_245),
.Y(n_311)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_311),
.Y(n_334)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_256),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_246),
.B1(n_263),
.B2(n_275),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_273),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_247),
.Y(n_315)
);

A2O1A1O1Ixp25_ASAP7_75t_L g316 ( 
.A1(n_275),
.A2(n_273),
.B(n_281),
.C(n_247),
.D(n_260),
.Y(n_316)
);

AOI32xp33_ASAP7_75t_L g335 ( 
.A1(n_316),
.A2(n_267),
.A3(n_270),
.B1(n_300),
.B2(n_291),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_317),
.B(n_287),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_314),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_318),
.B(n_329),
.Y(n_349)
);

AO22x1_ASAP7_75t_SL g320 ( 
.A1(n_286),
.A2(n_248),
.B1(n_261),
.B2(n_250),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_299),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_309),
.A2(n_261),
.B(n_267),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_323),
.A2(n_338),
.B(n_288),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_327),
.A2(n_290),
.B1(n_305),
.B2(n_304),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_306),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_316),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_301),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_267),
.B1(n_270),
.B2(n_294),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_336),
.A2(n_298),
.B1(n_311),
.B2(n_315),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_302),
.A2(n_270),
.B(n_308),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_319),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_342),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_337),
.B(n_310),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_331),
.B(n_307),
.Y(n_343)
);

NAND3xp33_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_303),
.C(n_340),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_344),
.A2(n_353),
.B1(n_326),
.B2(n_327),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_339),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_350),
.Y(n_372)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_346),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_329),
.B(n_295),
.Y(n_347)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_347),
.Y(n_375)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_324),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_348),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_330),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_351),
.A2(n_357),
.B(n_360),
.Y(n_367)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_324),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_358),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_321),
.A2(n_283),
.B1(n_313),
.B2(n_312),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_354),
.B(n_325),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_292),
.C(n_285),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_328),
.C(n_317),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_356),
.A2(n_361),
.B1(n_336),
.B2(n_299),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_338),
.A2(n_296),
.B(n_284),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_293),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_340),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_332),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_343),
.B(n_337),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_371),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_377),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_322),
.C(n_341),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_347),
.A2(n_321),
.B1(n_333),
.B2(n_326),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_368),
.A2(n_370),
.B1(n_373),
.B2(n_344),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_360),
.A2(n_322),
.B(n_323),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_369),
.A2(n_357),
.B(n_356),
.Y(n_389)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_376),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_354),
.B(n_328),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_379),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_355),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_382),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_355),
.Y(n_382)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_389),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_350),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_388),
.B(n_392),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_351),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_390),
.B(n_393),
.C(n_377),
.Y(n_396)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_378),
.Y(n_391)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_391),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_366),
.B(n_342),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_372),
.B(n_351),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_349),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_402),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_396),
.B(n_382),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_387),
.A2(n_356),
.B1(n_368),
.B2(n_365),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_369),
.Y(n_410)
);

AOI322xp5_ASAP7_75t_L g401 ( 
.A1(n_386),
.A2(n_349),
.A3(n_365),
.B1(n_378),
.B2(n_375),
.C1(n_345),
.C2(n_358),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_401),
.A2(n_359),
.B(n_374),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_375),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_407),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_405),
.B(n_403),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_381),
.C(n_384),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_380),
.C(n_389),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_408),
.B(n_409),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_374),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_411),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_397),
.Y(n_411)
);

AOI21x1_ASAP7_75t_L g414 ( 
.A1(n_406),
.A2(n_402),
.B(n_396),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_414),
.B(n_403),
.C(n_393),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_410),
.A2(n_400),
.B1(n_394),
.B2(n_399),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_415),
.B(n_416),
.Y(n_422)
);

OA21x2_ASAP7_75t_L g417 ( 
.A1(n_408),
.A2(n_356),
.B(n_400),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_417),
.B(n_367),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_412),
.B(n_407),
.Y(n_419)
);

NOR2x1_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_418),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_420),
.B(n_421),
.C(n_423),
.Y(n_424)
);

AO221x1_ASAP7_75t_L g423 ( 
.A1(n_413),
.A2(n_370),
.B1(n_335),
.B2(n_346),
.C(n_367),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_425),
.A2(n_426),
.B(n_361),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_418),
.C(n_417),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_424),
.B(n_420),
.C(n_380),
.Y(n_427)
);

OAI321xp33_ASAP7_75t_L g429 ( 
.A1(n_427),
.A2(n_428),
.A3(n_348),
.B1(n_352),
.B2(n_332),
.C(n_334),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_429),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_334),
.Y(n_431)
);


endmodule