module fake_jpeg_16003_n_66 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_66);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_66;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_24;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_43;
wire n_37;
wire n_29;
wire n_50;
wire n_32;

INVx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_6),
.B(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_11),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2x1_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_3),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_46),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_7),
.B1(n_10),
.B2(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_39),
.B1(n_34),
.B2(n_37),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_29),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_42),
.B(n_48),
.Y(n_58)
);

NOR4xp25_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_58),
.C(n_54),
.D(n_51),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_59),
.Y(n_62)
);

AOI322xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.A3(n_50),
.B1(n_52),
.B2(n_49),
.C1(n_59),
.C2(n_44),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_36),
.B(n_54),
.Y(n_63)
);

OAI31xp33_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_47),
.A3(n_50),
.B(n_53),
.Y(n_65)
);

XNOR2x2_ASAP7_75t_SL g66 ( 
.A(n_65),
.B(n_47),
.Y(n_66)
);


endmodule