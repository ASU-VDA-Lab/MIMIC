module fake_aes_101_n_16 (n_1, n_2, n_0, n_16);
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
INVx3_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
HB1xp67_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
CKINVDCx5p33_ASAP7_75t_R g5 ( .A(n_4), .Y(n_5) );
INVx2_ASAP7_75t_SL g6 ( .A(n_3), .Y(n_6) );
AND2x4_ASAP7_75t_SL g7 ( .A(n_6), .B(n_3), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
INVxp33_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_7), .B(n_6), .Y(n_10) );
AOI22xp33_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_5), .B1(n_1), .B2(n_0), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_10), .B(n_0), .Y(n_12) );
INVxp33_ASAP7_75t_SL g13 ( .A(n_11), .Y(n_13) );
A2O1A1Ixp33_ASAP7_75t_L g14 ( .A1(n_12), .A2(n_10), .B(n_1), .C(n_2), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
OAI21xp5_ASAP7_75t_L g16 ( .A1(n_15), .A2(n_13), .B(n_1), .Y(n_16) );
endmodule