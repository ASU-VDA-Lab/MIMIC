module fake_aes_1588_n_27 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_27);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_6), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_0), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g16 ( .A(n_12), .B(n_10), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_7), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_9), .Y(n_18) );
A2O1A1Ixp33_ASAP7_75t_L g19 ( .A1(n_14), .A2(n_1), .B(n_2), .C(n_3), .Y(n_19) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_13), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_20), .B(n_15), .Y(n_21) );
AND2x4_ASAP7_75t_L g22 ( .A(n_21), .B(n_20), .Y(n_22) );
OAI31xp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_19), .A3(n_2), .B(n_3), .Y(n_23) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_23), .B(n_22), .Y(n_24) );
NAND3xp33_ASAP7_75t_SL g25 ( .A(n_24), .B(n_23), .C(n_18), .Y(n_25) );
AOI22xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_17), .B1(n_16), .B2(n_4), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_5), .B1(n_8), .B2(n_11), .Y(n_27) );
endmodule