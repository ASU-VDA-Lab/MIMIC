module fake_jpeg_14349_n_199 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_199);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_0),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_88),
.Y(n_98)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_90),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_62),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_57),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_24),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_75),
.B1(n_66),
.B2(n_57),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_74),
.B1(n_56),
.B2(n_58),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_81),
.B1(n_75),
.B2(n_60),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_56),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_81),
.B1(n_60),
.B2(n_77),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_70),
.B1(n_77),
.B2(n_69),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_67),
.B1(n_70),
.B2(n_76),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_80),
.B(n_79),
.C(n_55),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_126),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_120),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_115),
.B1(n_117),
.B2(n_125),
.Y(n_129)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_73),
.B1(n_72),
.B2(n_68),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_127),
.Y(n_140)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_124),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_58),
.B1(n_64),
.B2(n_3),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_123),
.A2(n_4),
.B(n_7),
.Y(n_144)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_64),
.B1(n_2),
.B2(n_3),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_1),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_2),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_106),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_134),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_123),
.B(n_115),
.C(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_136),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_25),
.C(n_50),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_113),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_138),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_26),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_149),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_128),
.A2(n_30),
.B1(n_47),
.B2(n_46),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_31),
.B1(n_45),
.B2(n_44),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_108),
.B(n_9),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_9),
.B(n_10),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_11),
.B(n_12),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_10),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_156),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_155),
.B1(n_163),
.B2(n_14),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_19),
.B1(n_41),
.B2(n_39),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_18),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_160),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_53),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_129),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_17),
.B1(n_36),
.B2(n_35),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_11),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_146),
.C(n_142),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_169),
.B(n_170),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_129),
.B(n_148),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g182 ( 
.A1(n_174),
.A2(n_163),
.B1(n_161),
.B2(n_157),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_143),
.C(n_140),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_165),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_178),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_13),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_174),
.A2(n_155),
.B1(n_151),
.B2(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_182),
.A2(n_186),
.B(n_180),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_183),
.C(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_190),
.C(n_182),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_188),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_187),
.C(n_185),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_193),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_179),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_180),
.B1(n_185),
.B2(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_196),
.B(n_182),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_197),
.B(n_173),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_23),
.Y(n_199)
);


endmodule