module fake_jpeg_17861_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g37 ( 
.A(n_17),
.B(n_8),
.CON(n_37),
.SN(n_37)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_39),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_24),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_55),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_20),
.B1(n_23),
.B2(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_58),
.B1(n_16),
.B2(n_24),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_52),
.Y(n_81)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_54),
.A2(n_28),
.B1(n_33),
.B2(n_27),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_35),
.A2(n_23),
.B1(n_32),
.B2(n_25),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_40),
.B1(n_43),
.B2(n_41),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_93),
.B1(n_71),
.B2(n_63),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_43),
.B1(n_41),
.B2(n_26),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_70),
.A2(n_78),
.B1(n_48),
.B2(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_65),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_60),
.C(n_56),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_73),
.B(n_91),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_86),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_75),
.Y(n_100)
);

NAND2x1_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_43),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_76),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_42),
.C(n_38),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_89),
.C(n_17),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_26),
.B1(n_25),
.B2(n_32),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_39),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_21),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_80),
.B(n_84),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_48),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_32),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_64),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_88),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_33),
.B(n_28),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_0),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_94),
.B1(n_61),
.B2(n_53),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_48),
.B(n_17),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_18),
.B1(n_17),
.B2(n_31),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_97),
.Y(n_133)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_19),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_104),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_19),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_108),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_111),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_69),
.Y(n_108)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_117),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_119),
.B(n_90),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_42),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_122),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_68),
.B(n_31),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_115),
.B(n_84),
.Y(n_126)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_19),
.Y(n_117)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_78),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_60),
.C(n_65),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_121),
.A2(n_72),
.B1(n_68),
.B2(n_74),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_126),
.A2(n_138),
.B(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_68),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_141),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_80),
.B1(n_72),
.B2(n_61),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_136),
.B1(n_106),
.B2(n_113),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_140),
.B1(n_111),
.B2(n_122),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_86),
.B1(n_85),
.B2(n_67),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_89),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_137),
.B(n_146),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_90),
.B(n_76),
.C(n_91),
.D(n_82),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_96),
.A2(n_71),
.B1(n_76),
.B2(n_87),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_31),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_96),
.A2(n_92),
.B(n_31),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_102),
.B(n_19),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_56),
.C(n_82),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_109),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_149),
.A2(n_138),
.B1(n_147),
.B2(n_135),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_150),
.B(n_151),
.Y(n_197)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_168),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_100),
.Y(n_157)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_97),
.B1(n_100),
.B2(n_95),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_159),
.A2(n_164),
.B1(n_165),
.B2(n_173),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_104),
.Y(n_161)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_134),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_133),
.A2(n_85),
.B1(n_95),
.B2(n_108),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_101),
.B1(n_118),
.B2(n_53),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_85),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_171),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_131),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_129),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_144),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_22),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_172),
.C(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_31),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_31),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_127),
.A2(n_133),
.B1(n_136),
.B2(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_118),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_146),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_163),
.B(n_169),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g207 ( 
.A1(n_176),
.A2(n_193),
.B(n_194),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_170),
.C(n_172),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_140),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_180),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_156),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_153),
.Y(n_186)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_173),
.A2(n_123),
.B1(n_148),
.B2(n_145),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_187),
.A2(n_193),
.B1(n_196),
.B2(n_203),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_163),
.Y(n_206)
);

AO21x2_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_147),
.B(n_129),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_165),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_154),
.A2(n_138),
.B1(n_135),
.B2(n_130),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_137),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_203),
.B1(n_193),
.B2(n_181),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_202),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_151),
.A2(n_126),
.B1(n_120),
.B2(n_112),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_217),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_206),
.B(n_211),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_183),
.B(n_189),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_209),
.C(n_215),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_156),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_187),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_190),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_220),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_171),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_174),
.C(n_175),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_183),
.C(n_188),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_193),
.A2(n_168),
.B1(n_155),
.B2(n_98),
.Y(n_221)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_200),
.B1(n_195),
.B2(n_198),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_221),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_188),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_228),
.B(n_88),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_194),
.B(n_180),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_206),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_232),
.C(n_239),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_176),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_22),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_245),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_223),
.B1(n_56),
.B2(n_19),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_200),
.B1(n_192),
.B2(n_189),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_238),
.A2(n_236),
.B1(n_247),
.B2(n_235),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_196),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_182),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_244),
.C(n_247),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_9),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_214),
.B(n_192),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_212),
.B1(n_230),
.B2(n_222),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_88),
.C(n_22),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_219),
.C(n_224),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_251),
.Y(n_273)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_8),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_268),
.Y(n_272)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_205),
.B(n_204),
.C(n_212),
.D(n_226),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_257),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_267),
.B1(n_10),
.B2(n_14),
.Y(n_278)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_265),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_240),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_266),
.Y(n_274)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_239),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_232),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_241),
.C(n_30),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_271),
.C(n_281),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_241),
.C(n_30),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_266),
.Y(n_286)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_7),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_30),
.C(n_1),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_27),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_254),
.C(n_259),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_250),
.C(n_262),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_252),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_284),
.B(n_292),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_271),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_253),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_291),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_257),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_290),
.C(n_293),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_270),
.A2(n_265),
.B(n_7),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_269),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_30),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_297),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_295),
.B(n_275),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_273),
.B(n_6),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_11),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_279),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_277),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_301),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_30),
.C(n_27),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_305),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_11),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_286),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_308),
.Y(n_317)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_6),
.B(n_13),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_2),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_12),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_2),
.C(n_3),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_27),
.Y(n_313)
);

OAI21xp33_ASAP7_75t_L g323 ( 
.A1(n_313),
.A2(n_314),
.B(n_318),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_27),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

O2A1O1Ixp33_ASAP7_75t_SL g319 ( 
.A1(n_315),
.A2(n_316),
.B(n_309),
.C(n_303),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_299),
.B(n_1),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_320),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_3),
.C(n_4),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_324),
.C(n_5),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

AOI21x1_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_325),
.B(n_323),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_3),
.C(n_5),
.Y(n_324)
);

OAI21x1_ASAP7_75t_SL g325 ( 
.A1(n_312),
.A2(n_5),
.B(n_39),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_327),
.B1(n_328),
.B2(n_5),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_329),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_39),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_39),
.Y(n_332)
);


endmodule