module fake_aes_161_n_682 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_682);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_682;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g78 ( .A(n_66), .Y(n_78) );
INVxp67_ASAP7_75t_SL g79 ( .A(n_11), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_35), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_23), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_37), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_28), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_15), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_33), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_9), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_34), .Y(n_87) );
INVxp33_ASAP7_75t_L g88 ( .A(n_59), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_31), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_41), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_20), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_73), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_40), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_76), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_52), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_68), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_4), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_56), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_0), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_30), .Y(n_100) );
NOR2xp67_ASAP7_75t_L g101 ( .A(n_20), .B(n_43), .Y(n_101) );
BUFx2_ASAP7_75t_SL g102 ( .A(n_54), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_67), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_21), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_14), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_61), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_32), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_6), .Y(n_108) );
BUFx2_ASAP7_75t_SL g109 ( .A(n_63), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_36), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_15), .Y(n_111) );
INVxp33_ASAP7_75t_SL g112 ( .A(n_39), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_65), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_8), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_21), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_38), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_26), .Y(n_117) );
INVxp33_ASAP7_75t_L g118 ( .A(n_62), .Y(n_118) );
INVxp33_ASAP7_75t_L g119 ( .A(n_22), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_18), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_5), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_6), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_77), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_2), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_71), .Y(n_125) );
NOR2xp33_ASAP7_75t_R g126 ( .A(n_95), .B(n_29), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_91), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_90), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_97), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_97), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_124), .Y(n_131) );
NOR2xp33_ASAP7_75t_R g132 ( .A(n_96), .B(n_27), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
INVx6_ASAP7_75t_L g134 ( .A(n_111), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_107), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_78), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_111), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_78), .B(n_0), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_113), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_123), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_111), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_80), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_104), .B(n_1), .Y(n_145) );
INVxp67_ASAP7_75t_L g146 ( .A(n_86), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_112), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_81), .Y(n_148) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_81), .A2(n_42), .B(n_74), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_86), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_111), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_100), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_125), .B(n_1), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_83), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_87), .B(n_2), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_105), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_105), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_120), .Y(n_161) );
BUFx8_ASAP7_75t_L g162 ( .A(n_87), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_99), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_89), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_89), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_108), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_137), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_149), .Y(n_168) );
AO22x2_ASAP7_75t_L g169 ( .A1(n_131), .A2(n_106), .B1(n_98), .B2(n_117), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
INVx2_ASAP7_75t_SL g171 ( .A(n_133), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_146), .B(n_82), .Y(n_174) );
INVxp67_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_133), .B(n_122), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_137), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_147), .B(n_88), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
NAND2x1p5_ASAP7_75t_L g181 ( .A(n_153), .B(n_92), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_137), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_151), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_151), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_147), .B(n_118), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g188 ( .A1(n_163), .A2(n_121), .B1(n_108), .B2(n_79), .Y(n_188) );
AND3x1_ASAP7_75t_L g189 ( .A(n_145), .B(n_121), .C(n_92), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
AND2x4_ASAP7_75t_SL g191 ( .A(n_141), .B(n_120), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_153), .B(n_106), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_151), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_162), .B(n_119), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_142), .B(n_103), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_165), .A2(n_120), .B1(n_114), .B2(n_115), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_143), .Y(n_197) );
AOI22x1_ASAP7_75t_L g198 ( .A1(n_165), .A2(n_98), .B1(n_117), .B2(n_116), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_148), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_148), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_157), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_157), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_151), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_164), .Y(n_204) );
NOR3xp33_ASAP7_75t_L g205 ( .A(n_158), .B(n_116), .C(n_93), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_164), .Y(n_206) );
INVx4_ASAP7_75t_L g207 ( .A(n_149), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_144), .B(n_120), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_134), .Y(n_209) );
INVxp67_ASAP7_75t_L g210 ( .A(n_163), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_150), .B(n_110), .Y(n_211) );
NAND3x1_ASAP7_75t_L g212 ( .A(n_155), .B(n_93), .C(n_94), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_134), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_154), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_134), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_156), .B(n_166), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_134), .Y(n_217) );
INVx4_ASAP7_75t_L g218 ( .A(n_149), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_159), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_154), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_160), .B(n_110), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_154), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_129), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_130), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_154), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_162), .B(n_94), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_154), .Y(n_227) );
BUFx2_ASAP7_75t_L g228 ( .A(n_162), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_205), .B(n_138), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_185), .Y(n_230) );
INVxp33_ASAP7_75t_SL g231 ( .A(n_228), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_185), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_180), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_180), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_216), .B(n_126), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_226), .B(n_161), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_197), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_174), .B(n_140), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_197), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_199), .Y(n_240) );
OR2x6_ASAP7_75t_L g241 ( .A(n_228), .B(n_169), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_181), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_199), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_200), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_206), .Y(n_245) );
AND2x6_ASAP7_75t_SL g246 ( .A(n_179), .B(n_127), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_174), .B(n_132), .Y(n_247) );
INVx4_ASAP7_75t_L g248 ( .A(n_216), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_216), .B(n_85), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_216), .B(n_120), .Y(n_250) );
INVx4_ASAP7_75t_L g251 ( .A(n_181), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_171), .B(n_109), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_206), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_206), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_176), .B(n_140), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_176), .B(n_101), .Y(n_256) );
NAND2xp33_ASAP7_75t_R g257 ( .A(n_187), .B(n_139), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_191), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_206), .Y(n_259) );
NOR2xp33_ASAP7_75t_R g260 ( .A(n_210), .B(n_139), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_200), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_181), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_169), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_171), .B(n_109), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_211), .B(n_102), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_208), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_194), .B(n_135), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_176), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_176), .B(n_3), .Y(n_269) );
NOR2xp33_ASAP7_75t_R g270 ( .A(n_175), .B(n_135), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_201), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_211), .B(n_3), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_201), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_211), .B(n_102), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_211), .B(n_128), .Y(n_275) );
AO22x1_ASAP7_75t_L g276 ( .A1(n_168), .A2(n_128), .B1(n_5), .B2(n_7), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_221), .B(n_4), .Y(n_277) );
INVx5_ASAP7_75t_L g278 ( .A(n_225), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_202), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_191), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_202), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_169), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_191), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_169), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_204), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_221), .B(n_10), .Y(n_286) );
NOR3xp33_ASAP7_75t_SL g287 ( .A(n_188), .B(n_10), .C(n_11), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_221), .B(n_12), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_204), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_221), .B(n_12), .Y(n_290) );
CKINVDCx14_ASAP7_75t_R g291 ( .A(n_192), .Y(n_291) );
NOR3xp33_ASAP7_75t_SL g292 ( .A(n_195), .B(n_13), .C(n_14), .Y(n_292) );
INVx4_ASAP7_75t_L g293 ( .A(n_192), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_173), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_252), .A2(n_190), .B(n_168), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_251), .B(n_192), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_294), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_294), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_230), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_251), .B(n_192), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_264), .A2(n_190), .B(n_168), .Y(n_301) );
OR2x6_ASAP7_75t_L g302 ( .A(n_251), .B(n_212), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_233), .Y(n_303) );
NOR2x1_ASAP7_75t_SL g304 ( .A(n_241), .B(n_168), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_242), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_230), .B(n_219), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_242), .Y(n_307) );
AOI222xp33_ASAP7_75t_L g308 ( .A1(n_238), .A2(n_219), .B1(n_224), .B2(n_223), .C1(n_208), .C2(n_196), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_265), .A2(n_190), .B(n_207), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_293), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_231), .B(n_223), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_291), .A2(n_189), .B1(n_212), .B2(n_224), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_233), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_271), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_293), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_274), .A2(n_235), .B(n_249), .Y(n_316) );
NOR2x1_ASAP7_75t_L g317 ( .A(n_275), .B(n_173), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_271), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_232), .B(n_178), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_231), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_248), .B(n_178), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_234), .A2(n_190), .B(n_207), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_232), .B(n_207), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_234), .Y(n_324) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_247), .B(n_198), .C(n_218), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_263), .A2(n_198), .B1(n_218), .B2(n_207), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_255), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_241), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_241), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_262), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_267), .B(n_218), .Y(n_332) );
BUFx4_ASAP7_75t_SL g333 ( .A(n_246), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_241), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_262), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_263), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_237), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_284), .A2(n_218), .B1(n_190), .B2(n_209), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_248), .B(n_190), .Y(n_339) );
NAND2xp33_ASAP7_75t_L g340 ( .A(n_272), .B(n_227), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_293), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_269), .A2(n_209), .B1(n_213), .B2(n_215), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_260), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_272), .A2(n_213), .B1(n_215), .B2(n_217), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_320), .A2(n_280), .B1(n_248), .B2(n_257), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_327), .A2(n_238), .B1(n_255), .B2(n_272), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_343), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_296), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_305), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_322), .A2(n_277), .B(n_290), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_340), .A2(n_269), .B1(n_288), .B2(n_286), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_297), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_314), .Y(n_353) );
AOI21xp33_ASAP7_75t_L g354 ( .A1(n_311), .A2(n_280), .B(n_258), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g355 ( .A1(n_299), .A2(n_270), .B1(n_287), .B2(n_236), .C(n_256), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_314), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_296), .B(n_268), .Y(n_357) );
NAND2xp33_ASAP7_75t_R g358 ( .A(n_320), .B(n_286), .Y(n_358) );
AO31x2_ASAP7_75t_L g359 ( .A1(n_304), .A2(n_239), .A3(n_243), .B(n_244), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g360 ( .A1(n_343), .A2(n_288), .B1(n_286), .B2(n_269), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_319), .B(n_229), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_335), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_297), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_296), .B(n_268), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_323), .A2(n_288), .B1(n_336), .B2(n_319), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_298), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_295), .A2(n_243), .B(n_240), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_298), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_303), .Y(n_369) );
NOR2xp33_ASAP7_75t_SL g370 ( .A(n_328), .B(n_283), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_303), .Y(n_371) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_336), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_340), .A2(n_240), .B(n_237), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_313), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_353), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_352), .B(n_335), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_355), .A2(n_256), .B1(n_323), .B2(n_282), .Y(n_377) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_350), .A2(n_301), .B(n_309), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_360), .A2(n_236), .B1(n_302), .B2(n_332), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_346), .A2(n_236), .B1(n_302), .B2(n_317), .Y(n_380) );
AOI22xp33_ASAP7_75t_SL g381 ( .A1(n_348), .A2(n_328), .B1(n_334), .B2(n_329), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_361), .A2(n_256), .B1(n_276), .B2(n_292), .C(n_306), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_351), .A2(n_334), .B1(n_300), .B2(n_312), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_352), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_351), .A2(n_313), .B1(n_337), .B2(n_324), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_370), .B(n_345), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_348), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_363), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_363), .B(n_324), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_366), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_354), .A2(n_302), .B1(n_300), .B2(n_306), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_362), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_353), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_366), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_356), .Y(n_395) );
OAI21xp5_ASAP7_75t_SL g396 ( .A1(n_365), .A2(n_300), .B(n_308), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_357), .A2(n_302), .B1(n_229), .B2(n_337), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_368), .A2(n_276), .B1(n_316), .B2(n_229), .C(n_239), .Y(n_399) );
OAI211xp5_ASAP7_75t_L g400 ( .A1(n_372), .A2(n_330), .B(n_342), .C(n_305), .Y(n_400) );
OAI21x1_ASAP7_75t_L g401 ( .A1(n_350), .A2(n_326), .B(n_338), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_384), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_384), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_382), .A2(n_357), .B1(n_364), .B2(n_371), .Y(n_404) );
OAI22xp5_ASAP7_75t_SL g405 ( .A1(n_391), .A2(n_347), .B1(n_333), .B2(n_358), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_385), .A2(n_371), .B1(n_369), .B2(n_368), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_376), .Y(n_407) );
NOR2x2_ASAP7_75t_L g408 ( .A(n_375), .B(n_356), .Y(n_408) );
INVx5_ASAP7_75t_SL g409 ( .A(n_376), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_396), .A2(n_374), .B1(n_369), .B2(n_357), .C(n_364), .Y(n_410) );
OR2x6_ASAP7_75t_L g411 ( .A(n_396), .B(n_362), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_376), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_389), .B(n_374), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_388), .B(n_359), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_388), .B(n_357), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_376), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_375), .Y(n_418) );
AO21x2_ASAP7_75t_L g419 ( .A1(n_378), .A2(n_373), .B(n_367), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_382), .A2(n_364), .B1(n_344), .B2(n_266), .C(n_325), .Y(n_420) );
OAI31xp33_ASAP7_75t_L g421 ( .A1(n_400), .A2(n_364), .A3(n_349), .B(n_261), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_389), .B(n_359), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_392), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_390), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_379), .A2(n_310), .B1(n_341), .B2(n_315), .C(n_266), .Y(n_425) );
OAI31xp33_ASAP7_75t_SL g426 ( .A1(n_400), .A2(n_367), .A3(n_318), .B(n_331), .Y(n_426) );
AND2x2_ASAP7_75t_SL g427 ( .A(n_385), .B(n_305), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_386), .A2(n_335), .B1(n_349), .B2(n_307), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_380), .A2(n_310), .B1(n_315), .B2(n_341), .C(n_321), .Y(n_429) );
AO21x2_ASAP7_75t_L g430 ( .A1(n_378), .A2(n_304), .B(n_318), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_393), .Y(n_431) );
OA21x2_ASAP7_75t_L g432 ( .A1(n_378), .A2(n_331), .B(n_261), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_393), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_383), .A2(n_335), .B1(n_349), .B2(n_307), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_377), .A2(n_335), .B1(n_349), .B2(n_273), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_377), .A2(n_341), .B1(n_315), .B2(n_310), .C(n_268), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_390), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_415), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_426), .B(n_399), .C(n_398), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_432), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_422), .B(n_393), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_422), .B(n_395), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_415), .B(n_395), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_433), .B(n_395), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_423), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_430), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_432), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_402), .B(n_394), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_432), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_402), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
OAI21x1_ASAP7_75t_L g452 ( .A1(n_432), .A2(n_401), .B(n_394), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_410), .A2(n_399), .B1(n_389), .B2(n_387), .C(n_383), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_414), .B(n_397), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_414), .B(n_397), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_413), .Y(n_456) );
OAI222xp33_ASAP7_75t_L g457 ( .A1(n_411), .A2(n_381), .B1(n_387), .B2(n_392), .C1(n_307), .C2(n_359), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_403), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_411), .A2(n_381), .B1(n_401), .B2(n_273), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_424), .B(n_359), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_411), .B(n_359), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_413), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_424), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_437), .B(n_401), .Y(n_464) );
CKINVDCx14_ASAP7_75t_R g465 ( .A(n_405), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_437), .B(n_285), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_423), .B(n_289), .Y(n_467) );
AO21x2_ASAP7_75t_L g468 ( .A1(n_435), .A2(n_250), .B(n_281), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_413), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_418), .B(n_289), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_418), .B(n_13), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_418), .Y(n_472) );
INVx3_ASAP7_75t_L g473 ( .A(n_430), .Y(n_473) );
INVx5_ASAP7_75t_L g474 ( .A(n_411), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_431), .B(n_16), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_431), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_406), .B(n_431), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_407), .B(n_16), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_408), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_412), .B(n_244), .Y(n_480) );
AOI221x1_ASAP7_75t_L g481 ( .A1(n_406), .A2(n_434), .B1(n_405), .B2(n_416), .C(n_426), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_417), .B(n_281), .Y(n_482) );
NOR3xp33_ASAP7_75t_SL g483 ( .A(n_425), .B(n_217), .C(n_279), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_419), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_411), .B(n_17), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_404), .B(n_279), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_419), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_409), .B(n_17), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_419), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_454), .B(n_409), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_460), .B(n_430), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_454), .B(n_409), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_445), .Y(n_493) );
BUFx2_ASAP7_75t_L g494 ( .A(n_472), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_444), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_450), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_441), .B(n_409), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_440), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_451), .Y(n_499) );
NAND2xp33_ASAP7_75t_R g500 ( .A(n_483), .B(n_18), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_455), .B(n_409), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_460), .B(n_427), .Y(n_502) );
NOR2xp67_ASAP7_75t_SL g503 ( .A(n_474), .B(n_421), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_451), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_458), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_465), .A2(n_427), .B1(n_434), .B2(n_435), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_438), .B(n_427), .Y(n_507) );
OAI31xp33_ASAP7_75t_SL g508 ( .A1(n_479), .A2(n_421), .A3(n_420), .B(n_436), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_455), .B(n_428), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_457), .A2(n_429), .B(n_339), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_458), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_438), .B(n_19), .Y(n_512) );
AND2x2_ASAP7_75t_SL g513 ( .A(n_461), .B(n_339), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_441), .B(n_19), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_463), .B(n_245), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_444), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_463), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_479), .B(n_245), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_472), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_442), .B(n_24), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_448), .B(n_245), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_448), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_442), .B(n_478), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_472), .B(n_25), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_488), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_443), .B(n_259), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_488), .B(n_44), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_478), .B(n_259), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_440), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_461), .B(n_45), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_443), .B(n_254), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_440), .Y(n_532) );
NAND2xp33_ASAP7_75t_SL g533 ( .A(n_485), .B(n_339), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_471), .B(n_253), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_439), .A2(n_253), .B(n_254), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_485), .B(n_46), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_471), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_475), .B(n_47), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_447), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_475), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_461), .B(n_48), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_466), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_474), .A2(n_278), .B1(n_170), .B2(n_227), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_456), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_439), .A2(n_170), .B(n_227), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_453), .A2(n_461), .B1(n_474), .B2(n_459), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_456), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_453), .B(n_49), .Y(n_548) );
BUFx3_ASAP7_75t_L g549 ( .A(n_493), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_525), .B(n_474), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_522), .B(n_477), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_533), .A2(n_474), .B(n_473), .C(n_446), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_500), .A2(n_474), .B1(n_486), .B2(n_477), .Y(n_553) );
OAI221xp5_ASAP7_75t_SL g554 ( .A1(n_546), .A2(n_486), .B1(n_489), .B2(n_487), .C(n_467), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_519), .B(n_474), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_495), .B(n_489), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_533), .B(n_446), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_506), .A2(n_467), .B1(n_466), .B2(n_480), .Y(n_558) );
OAI21xp33_ASAP7_75t_L g559 ( .A1(n_508), .A2(n_487), .B(n_446), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_496), .Y(n_560) );
AOI33xp33_ASAP7_75t_L g561 ( .A1(n_514), .A2(n_484), .A3(n_447), .B1(n_449), .B2(n_481), .B3(n_469), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_513), .B(n_446), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_516), .B(n_469), .Y(n_563) );
NAND2xp33_ASAP7_75t_SL g564 ( .A(n_503), .B(n_468), .Y(n_564) );
NAND4xp25_ASAP7_75t_L g565 ( .A(n_518), .B(n_481), .C(n_473), .D(n_482), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_502), .B(n_456), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g567 ( .A1(n_512), .A2(n_484), .B1(n_473), .B2(n_482), .C(n_447), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_523), .B(n_469), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_542), .B(n_464), .Y(n_569) );
OAI321xp33_ASAP7_75t_L g570 ( .A1(n_536), .A2(n_541), .A3(n_530), .B1(n_527), .B2(n_548), .C(n_514), .Y(n_570) );
AOI222xp33_ASAP7_75t_L g571 ( .A1(n_512), .A2(n_462), .B1(n_476), .B2(n_449), .C1(n_484), .C2(n_473), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_502), .B(n_476), .Y(n_572) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_503), .A2(n_480), .B1(n_464), .B2(n_449), .C(n_470), .Y(n_573) );
O2A1O1Ixp5_ASAP7_75t_L g574 ( .A1(n_509), .A2(n_476), .B(n_462), .C(n_470), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_513), .B(n_462), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_490), .B(n_468), .Y(n_576) );
AOI22xp33_ASAP7_75t_SL g577 ( .A1(n_530), .A2(n_468), .B1(n_452), .B2(n_53), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_498), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_494), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_497), .A2(n_468), .B1(n_452), .B2(n_55), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g581 ( .A1(n_510), .A2(n_177), .B(n_182), .Y(n_581) );
OAI222xp33_ASAP7_75t_L g582 ( .A1(n_497), .A2(n_492), .B1(n_501), .B2(n_541), .C1(n_494), .C2(n_519), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_521), .B(n_50), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_520), .A2(n_51), .B1(n_57), .B2(n_58), .Y(n_584) );
OAI21xp5_ASAP7_75t_L g585 ( .A1(n_520), .A2(n_535), .B(n_524), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_543), .A2(n_182), .B(n_184), .Y(n_586) );
OAI221xp5_ASAP7_75t_L g587 ( .A1(n_528), .A2(n_182), .B1(n_184), .B2(n_193), .C(n_177), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_L g588 ( .A1(n_515), .A2(n_167), .B(n_184), .C(n_193), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_491), .B(n_60), .Y(n_589) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_524), .B(n_64), .Y(n_590) );
NAND2x1p5_ASAP7_75t_L g591 ( .A(n_526), .B(n_69), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_498), .Y(n_592) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_538), .A2(n_177), .B1(n_203), .B2(n_193), .C(n_167), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_504), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_491), .B(n_70), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_504), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_507), .A2(n_72), .B1(n_75), .B2(n_167), .Y(n_597) );
OAI21xp33_ASAP7_75t_SL g598 ( .A1(n_507), .A2(n_170), .B(n_214), .Y(n_598) );
AND3x2_ASAP7_75t_L g599 ( .A(n_555), .B(n_517), .C(n_505), .Y(n_599) );
NAND4xp75_ASAP7_75t_L g600 ( .A(n_553), .B(n_540), .C(n_537), .D(n_517), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_549), .B(n_505), .Y(n_601) );
NOR3xp33_ASAP7_75t_SL g602 ( .A(n_565), .B(n_570), .C(n_564), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_563), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_551), .B(n_511), .Y(n_604) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_580), .A2(n_526), .B(n_531), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_570), .B(n_499), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_582), .B(n_547), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_556), .B(n_529), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_578), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_560), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_567), .B(n_529), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_592), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_571), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_571), .B(n_532), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_594), .Y(n_615) );
NOR3xp33_ASAP7_75t_SL g616 ( .A(n_558), .B(n_534), .C(n_545), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_596), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_568), .B(n_547), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_569), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_558), .A2(n_544), .B1(n_539), .B2(n_532), .Y(n_620) );
OAI21xp5_ASAP7_75t_SL g621 ( .A1(n_577), .A2(n_544), .B(n_539), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_559), .A2(n_214), .B1(n_203), .B2(n_186), .C(n_183), .Y(n_622) );
NOR4xp25_ASAP7_75t_SL g623 ( .A(n_554), .B(n_214), .C(n_203), .D(n_186), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_566), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_572), .Y(n_625) );
NAND4xp25_ASAP7_75t_SL g626 ( .A(n_561), .B(n_172), .C(n_183), .D(n_220), .Y(n_626) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_591), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_591), .A2(n_590), .B1(n_573), .B2(n_585), .Y(n_628) );
NOR2xp67_ASAP7_75t_SL g629 ( .A(n_589), .B(n_225), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_576), .B(n_172), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_574), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_595), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_L g633 ( .A1(n_602), .A2(n_585), .B(n_555), .C(n_580), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_632), .Y(n_634) );
AOI32xp33_ASAP7_75t_L g635 ( .A1(n_628), .A2(n_550), .A3(n_575), .B1(n_598), .B2(n_562), .Y(n_635) );
INVx8_ASAP7_75t_L g636 ( .A(n_627), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_601), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_613), .B(n_579), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_619), .B(n_583), .Y(n_639) );
OAI21xp33_ASAP7_75t_L g640 ( .A1(n_613), .A2(n_581), .B(n_557), .Y(n_640) );
OAI21xp33_ASAP7_75t_L g641 ( .A1(n_602), .A2(n_581), .B(n_552), .Y(n_641) );
XNOR2x1_ASAP7_75t_L g642 ( .A(n_600), .B(n_590), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_621), .A2(n_584), .B(n_597), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_606), .B(n_588), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g645 ( .A(n_631), .B(n_593), .C(n_587), .Y(n_645) );
NOR2xp67_ASAP7_75t_L g646 ( .A(n_626), .B(n_586), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_601), .B(n_220), .Y(n_647) );
O2A1O1Ixp33_ASAP7_75t_L g648 ( .A1(n_616), .A2(n_222), .B(n_225), .C(n_278), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_614), .B(n_222), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_603), .Y(n_650) );
OA22x2_ASAP7_75t_L g651 ( .A1(n_599), .A2(n_225), .B1(n_278), .B2(n_605), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_607), .B(n_278), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_651), .A2(n_623), .B(n_620), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_633), .A2(n_620), .B1(n_616), .B2(n_627), .Y(n_654) );
OAI221xp5_ASAP7_75t_L g655 ( .A1(n_635), .A2(n_611), .B1(n_604), .B2(n_608), .C(n_617), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_649), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_638), .A2(n_625), .B1(n_624), .B2(n_610), .C(n_615), .Y(n_657) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_634), .Y(n_658) );
NOR2x1_ASAP7_75t_L g659 ( .A(n_642), .B(n_627), .Y(n_659) );
CKINVDCx5p33_ASAP7_75t_R g660 ( .A(n_650), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_641), .B(n_627), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_637), .B(n_599), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_652), .Y(n_663) );
OAI211xp5_ASAP7_75t_L g664 ( .A1(n_640), .A2(n_644), .B(n_643), .C(n_648), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_639), .A2(n_629), .B1(n_630), .B2(n_618), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_645), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_646), .A2(n_622), .B1(n_609), .B2(n_612), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_647), .A2(n_278), .B1(n_636), .B2(n_613), .C(n_638), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_636), .Y(n_669) );
NOR3xp33_ASAP7_75t_L g670 ( .A(n_644), .B(n_641), .C(n_652), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_656), .Y(n_671) );
BUFx10_ASAP7_75t_L g672 ( .A(n_658), .Y(n_672) );
INVx1_ASAP7_75t_SL g673 ( .A(n_660), .Y(n_673) );
OAI221xp5_ASAP7_75t_R g674 ( .A1(n_670), .A2(n_669), .B1(n_667), .B2(n_664), .C(n_665), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_671), .Y(n_675) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_673), .B(n_666), .Y(n_676) );
NAND3xp33_ASAP7_75t_SL g677 ( .A(n_674), .B(n_654), .C(n_655), .Y(n_677) );
OR2x6_ASAP7_75t_L g678 ( .A(n_676), .B(n_672), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_675), .Y(n_679) );
OAI321xp33_ASAP7_75t_L g680 ( .A1(n_678), .A2(n_677), .A3(n_661), .B1(n_668), .B2(n_653), .C(n_672), .Y(n_680) );
OAI211xp5_ASAP7_75t_L g681 ( .A1(n_680), .A2(n_679), .B(n_678), .C(n_659), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_681), .A2(n_662), .B1(n_653), .B2(n_663), .C(n_657), .Y(n_682) );
endmodule