module fake_jpeg_12011_n_583 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_583);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_583;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_61),
.Y(n_166)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_63),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_67),
.Y(n_191)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_69),
.Y(n_194)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_29),
.B(n_17),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_71),
.B(n_77),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_74),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_29),
.B(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_79),
.B(n_88),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_80),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_81),
.Y(n_177)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_83),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_32),
.B(n_15),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_89),
.Y(n_189)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_32),
.B(n_0),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_91),
.B(n_94),
.Y(n_181)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_44),
.Y(n_92)
);

INVx5_ASAP7_75t_SL g195 ( 
.A(n_92),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_93),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_52),
.B(n_0),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_95),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_96),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_97),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_2),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_98),
.B(n_111),
.Y(n_192)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_106),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_108),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_20),
.Y(n_116)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_24),
.Y(n_119)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_39),
.Y(n_120)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_41),
.Y(n_123)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_53),
.B(n_2),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_124),
.B(n_26),
.Y(n_190)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_24),
.Y(n_125)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_126),
.Y(n_199)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_41),
.Y(n_127)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_61),
.A2(n_25),
.B1(n_48),
.B2(n_58),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_130),
.A2(n_152),
.B1(n_172),
.B2(n_38),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_25),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_141),
.B(n_43),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_53),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_145),
.B(n_147),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_56),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_119),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_149),
.B(n_190),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g151 ( 
.A(n_75),
.B(n_31),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_151),
.A2(n_42),
.B(n_44),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_64),
.A2(n_25),
.B1(n_48),
.B2(n_58),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_56),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_153),
.B(n_162),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_60),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_67),
.A2(n_48),
.B1(n_36),
.B2(n_51),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_36),
.C(n_35),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_173),
.A2(n_178),
.B(n_42),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_69),
.A2(n_45),
.B1(n_51),
.B2(n_49),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_174),
.A2(n_184),
.B1(n_187),
.B2(n_45),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_83),
.B(n_35),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_175),
.B(n_44),
.Y(n_254)
);

NAND2x1_ASAP7_75t_L g178 ( 
.A(n_82),
.B(n_42),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_110),
.B(n_60),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_203),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_72),
.A2(n_26),
.B1(n_55),
.B2(n_46),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_73),
.A2(n_26),
.B1(n_55),
.B2(n_46),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_86),
.A2(n_49),
.B(n_47),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g280 ( 
.A(n_193),
.B(n_7),
.C(n_8),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_95),
.B(n_47),
.Y(n_203)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_210),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_211),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_135),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_212),
.Y(n_329)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_154),
.Y(n_213)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_213),
.Y(n_303)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_215),
.Y(n_307)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_217),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_159),
.Y(n_218)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_218),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_219),
.B(n_220),
.Y(n_301)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_222),
.Y(n_306)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_133),
.Y(n_223)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_223),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_224),
.Y(n_310)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_135),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_225),
.Y(n_305)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_226),
.Y(n_322)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_142),
.Y(n_227)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_227),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_178),
.A2(n_43),
.B1(n_26),
.B2(n_116),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_228),
.A2(n_231),
.B1(n_263),
.B2(n_268),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_166),
.Y(n_230)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_230),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_155),
.A2(n_43),
.B1(n_26),
.B2(n_107),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_181),
.B(n_4),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_232),
.B(n_238),
.Y(n_315)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_233),
.Y(n_324)
);

NOR2x1_ASAP7_75t_R g309 ( 
.A(n_234),
.B(n_255),
.Y(n_309)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_235),
.Y(n_325)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_237),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_181),
.B(n_4),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_148),
.B(n_6),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_253),
.Y(n_289)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_240),
.Y(n_335)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

INVx11_ASAP7_75t_L g285 ( 
.A(n_241),
.Y(n_285)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_134),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_242),
.B(n_244),
.Y(n_284)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_200),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_243),
.Y(n_326)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_130),
.A2(n_78),
.B1(n_114),
.B2(n_112),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_245),
.A2(n_251),
.B1(n_260),
.B2(n_231),
.Y(n_327)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_138),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_249),
.Y(n_290)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_247),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

INVx13_ASAP7_75t_L g330 ( 
.A(n_248),
.Y(n_330)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_139),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_192),
.A2(n_96),
.B1(n_109),
.B2(n_104),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_250),
.A2(n_262),
.B1(n_272),
.B2(n_279),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_152),
.A2(n_115),
.B1(n_100),
.B2(n_93),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_128),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_256),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_148),
.B(n_6),
.Y(n_253)
);

AOI21xp33_ASAP7_75t_L g321 ( 
.A1(n_254),
.A2(n_261),
.B(n_270),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_141),
.A2(n_6),
.B(n_7),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_150),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_195),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_258),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_151),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_143),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_259),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_172),
.A2(n_81),
.B1(n_80),
.B2(n_43),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g262 ( 
.A1(n_175),
.A2(n_176),
.B1(n_169),
.B2(n_182),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_166),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_131),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_265),
.Y(n_313)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_144),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_140),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_266),
.B(n_267),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_197),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_196),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_131),
.B(n_7),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_269),
.B(n_273),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_151),
.B(n_43),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_192),
.B(n_7),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_274),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_129),
.A2(n_44),
.B1(n_38),
.B2(n_9),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_171),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_136),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_183),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_276),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_157),
.Y(n_276)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_170),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_278),
.Y(n_291)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_189),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_8),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_219),
.A2(n_132),
.B1(n_208),
.B2(n_177),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_282),
.A2(n_293),
.B1(n_314),
.B2(n_320),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_292),
.B(n_248),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_260),
.A2(n_251),
.B1(n_245),
.B2(n_229),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_221),
.B(n_174),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_294),
.B(n_299),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_216),
.B(n_188),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_185),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_300),
.B(n_225),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_258),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_262),
.A2(n_206),
.B1(n_205),
.B2(n_137),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_319),
.A2(n_323),
.B1(n_334),
.B2(n_241),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_228),
.A2(n_137),
.B1(n_160),
.B2(n_191),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_270),
.A2(n_161),
.B1(n_157),
.B2(n_160),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_327),
.A2(n_332),
.B1(n_276),
.B2(n_218),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_236),
.A2(n_155),
.B1(n_146),
.B2(n_191),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_261),
.B(n_146),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_214),
.C(n_278),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_234),
.A2(n_161),
.B1(n_194),
.B2(n_170),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_311),
.Y(n_336)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_336),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_301),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_337),
.B(n_374),
.C(n_295),
.Y(n_408)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_291),
.Y(n_339)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_339),
.Y(n_385)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_340),
.Y(n_390)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_297),
.Y(n_341)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_341),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_342),
.B(n_353),
.Y(n_388)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_297),
.Y(n_343)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_343),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_300),
.A2(n_255),
.B(n_248),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_344),
.A2(n_358),
.B(n_285),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_345),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_302),
.A2(n_194),
.B1(n_222),
.B2(n_277),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_346),
.A2(n_349),
.B1(n_355),
.B2(n_369),
.Y(n_413)
);

MAJx2_ASAP7_75t_L g407 ( 
.A(n_347),
.B(n_285),
.C(n_330),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_302),
.A2(n_263),
.B1(n_230),
.B2(n_247),
.Y(n_349)
);

BUFx5_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_304),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_351),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_286),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_352),
.Y(n_389)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_304),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_308),
.A2(n_212),
.B(n_274),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_354),
.A2(n_378),
.B(n_283),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_290),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_357),
.Y(n_379)
);

AO22x1_ASAP7_75t_SL g357 ( 
.A1(n_327),
.A2(n_201),
.B1(n_38),
.B2(n_10),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_299),
.B(n_8),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_359),
.B(n_303),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_281),
.B(n_14),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_362),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_315),
.B(n_8),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_361),
.B(n_377),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_310),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_296),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_373),
.Y(n_403)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_305),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_364),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_301),
.A2(n_9),
.B(n_11),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_365),
.B(n_371),
.Y(n_409)
);

BUFx24_ASAP7_75t_SL g366 ( 
.A(n_289),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_366),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_301),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_367),
.A2(n_372),
.B1(n_306),
.B2(n_295),
.Y(n_402)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_305),
.Y(n_368)
);

INVx6_ASAP7_75t_L g392 ( 
.A(n_368),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_294),
.A2(n_316),
.B1(n_281),
.B2(n_288),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_319),
.A2(n_12),
.B1(n_334),
.B2(n_316),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_370),
.A2(n_376),
.B1(n_296),
.B2(n_311),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_309),
.A2(n_12),
.B(n_292),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_293),
.A2(n_282),
.B1(n_320),
.B2(n_314),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_286),
.B(n_313),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_321),
.B(n_325),
.C(n_289),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_375),
.B(n_329),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_309),
.A2(n_325),
.B1(n_284),
.B2(n_326),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_312),
.B(n_287),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_331),
.A2(n_298),
.B(n_326),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_410),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_373),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_382),
.B(n_401),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_384),
.B(n_414),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_338),
.A2(n_328),
.B1(n_335),
.B2(n_324),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_393),
.A2(n_395),
.B1(n_402),
.B2(n_412),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_338),
.A2(n_328),
.B1(n_335),
.B2(n_324),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_344),
.A2(n_318),
.B(n_283),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_397),
.A2(n_384),
.B(n_405),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_348),
.B(n_283),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_400),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_358),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_404),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_376),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_337),
.C(n_347),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_408),
.B(n_351),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_348),
.B(n_306),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_339),
.B(n_306),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_411),
.B(n_362),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_372),
.A2(n_303),
.B1(n_307),
.B2(n_317),
.Y(n_412)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_391),
.Y(n_415)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_415),
.Y(n_467)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_416),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_418),
.B(n_445),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_419),
.A2(n_420),
.B(n_431),
.Y(n_447)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_391),
.Y(n_421)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_421),
.Y(n_475)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_399),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_422),
.B(n_425),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_413),
.A2(n_342),
.B1(n_340),
.B2(n_357),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_423),
.A2(n_438),
.B1(n_388),
.B2(n_402),
.Y(n_466)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_399),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_411),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_426),
.Y(n_450)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_427),
.Y(n_461)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_386),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_429),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_388),
.A2(n_346),
.B1(n_349),
.B2(n_370),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_430),
.A2(n_389),
.B1(n_398),
.B2(n_383),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_397),
.A2(n_354),
.B(n_371),
.Y(n_431)
);

HB1xp67_ASAP7_75t_SL g432 ( 
.A(n_406),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_432),
.A2(n_412),
.B1(n_383),
.B2(n_361),
.Y(n_471)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_433),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_396),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_436),
.Y(n_462)
);

NOR2xp67_ASAP7_75t_SL g437 ( 
.A(n_379),
.B(n_345),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_437),
.B(n_439),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_413),
.A2(n_357),
.B1(n_360),
.B2(n_374),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_404),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_401),
.A2(n_378),
.B(n_365),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_440),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_444),
.C(n_407),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_379),
.A2(n_367),
.B(n_356),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_443),
.B(n_400),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_408),
.B(n_363),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_403),
.B(n_343),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_388),
.A2(n_375),
.B(n_353),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_446),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_434),
.A2(n_390),
.B1(n_385),
.B2(n_382),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_449),
.A2(n_458),
.B1(n_460),
.B2(n_435),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_403),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_453),
.B(n_463),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_417),
.B(n_380),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_455),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_456),
.B(n_457),
.C(n_464),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_444),
.B(n_418),
.C(n_407),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_434),
.A2(n_390),
.B1(n_410),
.B2(n_398),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_409),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_419),
.B(n_389),
.C(n_409),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_466),
.A2(n_428),
.B1(n_430),
.B2(n_426),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_419),
.B(n_409),
.C(n_393),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_470),
.C(n_472),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_440),
.B(n_395),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_471),
.A2(n_431),
.B(n_443),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_420),
.B(n_341),
.C(n_394),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_477),
.A2(n_484),
.B1(n_485),
.B2(n_499),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_472),
.B(n_394),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_478),
.B(n_487),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_479),
.A2(n_486),
.B1(n_491),
.B2(n_493),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_SL g480 ( 
.A(n_464),
.B(n_424),
.C(n_437),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_480),
.B(n_496),
.C(n_481),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_448),
.B(n_438),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_448),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_466),
.A2(n_428),
.B1(n_424),
.B2(n_439),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_450),
.A2(n_441),
.B1(n_416),
.B2(n_433),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_380),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_451),
.Y(n_488)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_488),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_450),
.B(n_441),
.Y(n_489)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_489),
.Y(n_510)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_474),
.Y(n_490)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_490),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_459),
.A2(n_423),
.B1(n_429),
.B2(n_427),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_452),
.B(n_414),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_492),
.B(n_494),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_458),
.A2(n_425),
.B1(n_422),
.B2(n_421),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_474),
.Y(n_494)
);

AND2x2_ASAP7_75t_SL g495 ( 
.A(n_469),
.B(n_446),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_462),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_457),
.B(n_436),
.C(n_415),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_456),
.B(n_387),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_500),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_471),
.A2(n_387),
.B1(n_392),
.B2(n_336),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_473),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_SL g535 ( 
.A(n_503),
.B(n_504),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_497),
.B(n_470),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_483),
.B(n_447),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_505),
.B(n_493),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_447),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_509),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_483),
.B(n_463),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_476),
.Y(n_513)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_513),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_489),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_514),
.B(n_515),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_496),
.B(n_461),
.Y(n_515)
);

MAJx2_ASAP7_75t_L g522 ( 
.A(n_516),
.B(n_518),
.C(n_495),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_482),
.B(n_495),
.C(n_480),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_519),
.B(n_486),
.C(n_491),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_482),
.B(n_449),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_520),
.B(n_465),
.Y(n_536)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_522),
.Y(n_549)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_511),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_524),
.B(n_527),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_525),
.B(n_529),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_502),
.A2(n_479),
.B1(n_494),
.B2(n_490),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_517),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_530),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_501),
.B(n_484),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_512),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_506),
.A2(n_477),
.B1(n_485),
.B2(n_499),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_531),
.A2(n_533),
.B1(n_518),
.B2(n_527),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_532),
.B(n_502),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_520),
.B(n_468),
.C(n_500),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_533),
.B(n_505),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_SL g534 ( 
.A1(n_510),
.A2(n_462),
.B1(n_467),
.B2(n_475),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_534),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_536),
.B(n_516),
.C(n_506),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_539),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_525),
.A2(n_516),
.B(n_519),
.Y(n_540)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_540),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_541),
.B(n_543),
.Y(n_554)
);

INVxp33_ASAP7_75t_L g543 ( 
.A(n_521),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_544),
.B(n_547),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_545),
.B(n_535),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_531),
.A2(n_465),
.B(n_508),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_509),
.C(n_504),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g557 ( 
.A(n_548),
.B(n_550),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_532),
.B(n_503),
.C(n_507),
.Y(n_550)
);

NOR2x1_ASAP7_75t_L g551 ( 
.A(n_549),
.B(n_522),
.Y(n_551)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_551),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_542),
.A2(n_523),
.B1(n_475),
.B2(n_467),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_552),
.B(n_560),
.Y(n_566)
);

NOR2x1_ASAP7_75t_L g553 ( 
.A(n_549),
.B(n_526),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_550),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_555),
.B(n_537),
.Y(n_567)
);

OAI22x1_ASAP7_75t_L g560 ( 
.A1(n_540),
.A2(n_526),
.B1(n_535),
.B2(n_368),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_538),
.A2(n_546),
.B1(n_541),
.B2(n_545),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_561),
.B(n_364),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g562 ( 
.A1(n_558),
.A2(n_543),
.B(n_546),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_562),
.A2(n_564),
.B(n_559),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_554),
.B(n_548),
.C(n_547),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_565),
.B(n_569),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_567),
.B(n_555),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_556),
.B(n_392),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_568),
.B(n_350),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_571),
.A2(n_573),
.B(n_564),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_572),
.B(n_574),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_563),
.A2(n_551),
.B(n_553),
.Y(n_573)
);

AOI21x1_ASAP7_75t_SL g579 ( 
.A1(n_575),
.A2(n_576),
.B(n_560),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_570),
.A2(n_557),
.B(n_566),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_577),
.A2(n_561),
.B(n_556),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_578),
.A2(n_579),
.B(n_336),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g581 ( 
.A1(n_580),
.A2(n_330),
.B(n_317),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_SL g582 ( 
.A1(n_581),
.A2(n_307),
.B(n_322),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_582),
.B(n_322),
.Y(n_583)
);


endmodule