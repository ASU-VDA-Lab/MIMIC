module fake_jpeg_23608_n_265 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_149;
wire n_48;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_33),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_38),
.B(n_18),
.C(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_35),
.B(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_47),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_15),
.B1(n_24),
.B2(n_21),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_62),
.B1(n_66),
.B2(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_63),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_17),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_31),
.B1(n_30),
.B2(n_26),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_22),
.B1(n_28),
.B2(n_19),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_65),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_34),
.A2(n_22),
.B1(n_19),
.B2(n_28),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_72),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_34),
.B1(n_25),
.B2(n_33),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_66),
.B1(n_59),
.B2(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_34),
.B1(n_25),
.B2(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_23),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_25),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_65),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_1),
.B(n_3),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_79),
.B(n_80),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_41),
.B(n_39),
.C(n_37),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_39),
.B1(n_37),
.B2(n_36),
.Y(n_80)
);

AO22x1_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_36),
.B1(n_27),
.B2(n_20),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_86),
.B1(n_52),
.B2(n_54),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_27),
.B1(n_20),
.B2(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_92),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_43),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_51),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_18),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_97),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_98),
.B(n_81),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_102),
.Y(n_113)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_23),
.B(n_30),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_101),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_52),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_100),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_68),
.B(n_69),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_116),
.C(n_120),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_107),
.A2(n_67),
.B1(n_71),
.B2(n_54),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_128),
.B1(n_80),
.B2(n_70),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_71),
.B1(n_80),
.B2(n_52),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_123),
.B1(n_130),
.B2(n_101),
.Y(n_141)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_94),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_51),
.C(n_44),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_80),
.B1(n_65),
.B2(n_64),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_97),
.B1(n_91),
.B2(n_99),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_80),
.B1(n_64),
.B2(n_70),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_44),
.C(n_51),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_92),
.Y(n_146)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_125),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_136),
.B(n_143),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_89),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_138),
.B(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

CKINVDCx11_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_147),
.B1(n_155),
.B2(n_158),
.Y(n_177)
);

CKINVDCx10_ASAP7_75t_R g142 ( 
.A(n_134),
.Y(n_142)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_132),
.B(n_105),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_110),
.Y(n_144)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_149),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_88),
.B1(n_89),
.B2(n_102),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_26),
.Y(n_150)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_20),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_121),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_44),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_156),
.B(n_127),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_70),
.Y(n_154)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_64),
.B1(n_43),
.B2(n_84),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_1),
.Y(n_156)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_175),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_116),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_111),
.C(n_131),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_158),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_156),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_137),
.B(n_133),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_142),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_139),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_179),
.B1(n_126),
.B2(n_151),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_128),
.B1(n_141),
.B2(n_115),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_120),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_167),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_73),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_165),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_196),
.Y(n_208)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

OAI22x1_ASAP7_75t_SL g185 ( 
.A1(n_169),
.A2(n_153),
.B1(n_136),
.B2(n_149),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_187),
.B1(n_199),
.B2(n_87),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_190),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_135),
.B1(n_146),
.B2(n_155),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_178),
.B1(n_170),
.B2(n_160),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_SL g192 ( 
.A(n_168),
.B(n_143),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_192),
.A2(n_195),
.B(n_85),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_126),
.C(n_130),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_194),
.C(n_171),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_136),
.C(n_156),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_198),
.Y(n_216)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_161),
.A2(n_129),
.B1(n_113),
.B2(n_150),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_113),
.B1(n_129),
.B2(n_84),
.Y(n_200)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_187),
.C(n_191),
.Y(n_217)
);

OAI21x1_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_173),
.B(n_166),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_202),
.A2(n_203),
.B(n_209),
.Y(n_227)
);

XOR2x2_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_159),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_179),
.C(n_159),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_184),
.C(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_27),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_178),
.B(n_160),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_163),
.B1(n_129),
.B2(n_84),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_213),
.B1(n_188),
.B2(n_195),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_215),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_214),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_195),
.C(n_199),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_73),
.C(n_31),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_222),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_87),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_223),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_209),
.B(n_203),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_227),
.B(n_229),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_58),
.B1(n_48),
.B2(n_3),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_205),
.B1(n_216),
.B2(n_204),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_58),
.C(n_48),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_226),
.A2(n_228),
.B(n_208),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_58),
.C(n_4),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_236),
.C(n_237),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_215),
.B1(n_207),
.B2(n_3),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_237),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_219),
.A2(n_4),
.B(n_5),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_5),
.C(n_6),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_229),
.Y(n_240)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_224),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_8),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_5),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_7),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_7),
.C(n_8),
.Y(n_247)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_248),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_233),
.A3(n_232),
.B1(n_238),
.B2(n_11),
.C1(n_8),
.C2(n_13),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_253),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_242),
.C(n_243),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_9),
.Y(n_260)
);

AOI21x1_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_245),
.B(n_10),
.Y(n_255)
);

AOI21x1_ASAP7_75t_SL g259 ( 
.A1(n_255),
.A2(n_248),
.B(n_10),
.Y(n_259)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_252),
.B(n_257),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_260),
.C(n_9),
.Y(n_261)
);

AOI321xp33_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_76),
.C(n_95),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g263 ( 
.A(n_261),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_262),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_11),
.Y(n_265)
);


endmodule