module fake_netlist_5_1074_n_1785 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1785);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1785;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_85),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_112),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_83),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_22),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_156),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_29),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_0),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_37),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_3),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_74),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_56),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_19),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_106),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_34),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_68),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_65),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_61),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_34),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_21),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_107),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_101),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_104),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_51),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_23),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_108),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_120),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_134),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_14),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_10),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_143),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_20),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_37),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_151),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_9),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_60),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_94),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_55),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_29),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_149),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_76),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_171),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_3),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_91),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_93),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_66),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_144),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_84),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_57),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_70),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_62),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_9),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_169),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_148),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_14),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_46),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_24),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_97),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_115),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_16),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_79),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_133),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_71),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_127),
.Y(n_251)
);

INVxp33_ASAP7_75t_SL g252 ( 
.A(n_152),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_54),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_10),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_36),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_129),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_27),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_19),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_128),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_36),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_51),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_50),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_73),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_110),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_180),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_4),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_168),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_41),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_82),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_164),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_131),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_53),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_114),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_135),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_96),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_145),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_0),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_15),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_175),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_158),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_123),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_30),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_100),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_27),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_20),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_25),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_47),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_35),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_22),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_24),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_6),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_7),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_7),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_124),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_4),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_42),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_140),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_98),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_99),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_177),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_47),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_23),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_77),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_174),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_78),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_45),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_155),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_11),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_154),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_172),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_26),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_64),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_8),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_21),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_11),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_45),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_67),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_119),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_42),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_153),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_89),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_87),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_1),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_52),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_150),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_25),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_111),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_95),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_146),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_157),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_72),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_105),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_118),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_178),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_92),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_1),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_2),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_35),
.Y(n_338)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_141),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_142),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_33),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_69),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_15),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_8),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_28),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_130),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_58),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_103),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_6),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_33),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_113),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_88),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_122),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_48),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_243),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_208),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_208),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_208),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_208),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_181),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_220),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_206),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_182),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_208),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_315),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_225),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_226),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_223),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_183),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_315),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_315),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_214),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_207),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_227),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_213),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_217),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_331),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_315),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_306),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_285),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_259),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_285),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_234),
.Y(n_385)
);

NAND2xp33_ASAP7_75t_R g386 ( 
.A(n_195),
.B(n_199),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_237),
.B(n_2),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_351),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_235),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_274),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_276),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_222),
.B(n_5),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_249),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_236),
.Y(n_395)
);

NOR2xp67_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_5),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_215),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_240),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_241),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_299),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_256),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_304),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_247),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_353),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_254),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_245),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_246),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_260),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_184),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_321),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_203),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_253),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_184),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_248),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_250),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_251),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_228),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_263),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_265),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_253),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_273),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_261),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_321),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_279),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_280),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_266),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_278),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_228),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_291),
.Y(n_430)
);

INVxp33_ASAP7_75t_SL g431 ( 
.A(n_186),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_281),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_283),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_293),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_295),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_232),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_294),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_300),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_319),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_344),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_253),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_360),
.Y(n_442)
);

NOR2x1_ASAP7_75t_L g443 ( 
.A(n_387),
.B(n_232),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_361),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_356),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_356),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_349),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_367),
.B(n_252),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_357),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_357),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_409),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_358),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_376),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_368),
.B(n_271),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_271),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_359),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_417),
.B(n_320),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_417),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_375),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_364),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_376),
.B(n_343),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_419),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_364),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_385),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_365),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_R g470 ( 
.A(n_404),
.B(n_386),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_365),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_363),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_366),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_366),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_371),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_372),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_372),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_379),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_377),
.B(n_321),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_397),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_397),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_390),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_403),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_370),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_395),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_419),
.A2(n_267),
.B(n_204),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_417),
.B(n_320),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_381),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_R g491 ( 
.A(n_431),
.B(n_185),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_381),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_383),
.B(n_348),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_383),
.Y(n_494)
);

BUFx10_ASAP7_75t_L g495 ( 
.A(n_398),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_403),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_405),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_408),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_399),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_377),
.B(n_325),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_396),
.B(n_237),
.Y(n_502)
);

OA21x2_ASAP7_75t_L g503 ( 
.A1(n_384),
.A2(n_267),
.B(n_204),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_408),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_406),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_393),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_407),
.B(n_415),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_384),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_423),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_373),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_416),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_420),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_427),
.Y(n_515)
);

CKINVDCx8_ASAP7_75t_R g516 ( 
.A(n_410),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_388),
.B(n_193),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_427),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_428),
.Y(n_519)
);

INVx6_ASAP7_75t_L g520 ( 
.A(n_461),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_457),
.B(n_425),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_482),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_471),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_482),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_458),
.B(n_362),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_426),
.Y(n_526)
);

OR2x6_ASAP7_75t_L g527 ( 
.A(n_451),
.B(n_412),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_462),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_488),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_462),
.B(n_432),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_461),
.B(n_200),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_461),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_462),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_458),
.B(n_369),
.Y(n_534)
);

OR2x6_ASAP7_75t_L g535 ( 
.A(n_451),
.B(n_441),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_488),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_462),
.B(n_394),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_483),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_485),
.Y(n_539)
);

BUFx4f_ASAP7_75t_L g540 ( 
.A(n_503),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_446),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_461),
.B(n_489),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_489),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_470),
.B(n_389),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_506),
.B(n_389),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_448),
.B(n_414),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_471),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_456),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_442),
.B(n_418),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_489),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_485),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_496),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_489),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_496),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_444),
.B(n_422),
.Y(n_555)
);

AND2x6_ASAP7_75t_L g556 ( 
.A(n_502),
.B(n_200),
.Y(n_556)
);

AND2x2_ASAP7_75t_SL g557 ( 
.A(n_502),
.B(n_200),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_497),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_502),
.B(n_200),
.Y(n_559)
);

AO22x2_ASAP7_75t_L g560 ( 
.A1(n_480),
.A2(n_401),
.B1(n_378),
.B2(n_355),
.Y(n_560)
);

BUFx10_ASAP7_75t_L g561 ( 
.A(n_463),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_465),
.B(n_413),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_507),
.Y(n_563)
);

AND2x6_ASAP7_75t_L g564 ( 
.A(n_502),
.B(n_200),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_497),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_446),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_456),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_498),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_446),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_447),
.B(n_410),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_456),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_443),
.B(n_270),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_446),
.Y(n_573)
);

BUFx4f_ASAP7_75t_L g574 ( 
.A(n_503),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_460),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_446),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_468),
.B(n_433),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_517),
.B(n_428),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_517),
.B(n_440),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_501),
.B(n_421),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_447),
.B(n_388),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_460),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_491),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_460),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_466),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_443),
.B(n_298),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_469),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_469),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_466),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_498),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_517),
.A2(n_252),
.B1(n_270),
.B2(n_435),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_517),
.B(n_270),
.Y(n_592)
);

XNOR2x2_ASAP7_75t_SL g593 ( 
.A(n_516),
.B(n_219),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_445),
.B(n_305),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_446),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_484),
.B(n_437),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_503),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_499),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_503),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_445),
.B(n_309),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_453),
.B(n_430),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_449),
.B(n_317),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_449),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_466),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_L g605 ( 
.A(n_450),
.B(n_270),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_469),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_454),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_475),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_487),
.B(n_270),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_504),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_450),
.B(n_327),
.Y(n_611)
);

INVxp67_ASAP7_75t_SL g612 ( 
.A(n_452),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_453),
.Y(n_613)
);

AND2x2_ASAP7_75t_SL g614 ( 
.A(n_454),
.B(n_424),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_509),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_452),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_510),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_500),
.B(n_424),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_459),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_510),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_459),
.B(n_330),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_475),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_464),
.B(n_332),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_505),
.B(n_205),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_511),
.B(n_430),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_464),
.B(n_216),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_515),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_513),
.B(n_438),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_515),
.B(n_518),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_518),
.A2(n_440),
.B1(n_439),
.B2(n_435),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_475),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_519),
.B(n_493),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_476),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_509),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_476),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_519),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_467),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_476),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_514),
.B(n_218),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_509),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_477),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_495),
.B(n_221),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_490),
.B(n_439),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_455),
.A2(n_382),
.B1(n_402),
.B2(n_400),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_473),
.B(n_474),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_495),
.B(n_434),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_477),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_474),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_478),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_477),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_L g652 ( 
.A(n_478),
.B(n_339),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_509),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_495),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_479),
.Y(n_655)
);

BUFx8_ASAP7_75t_SL g656 ( 
.A(n_472),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_479),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_486),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_495),
.B(n_391),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_479),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_481),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_481),
.B(n_493),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_481),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_509),
.B(n_494),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_540),
.A2(n_231),
.B(n_230),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_570),
.B(n_516),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_647),
.B(n_525),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_545),
.B(n_185),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_557),
.A2(n_292),
.B1(n_290),
.B2(n_339),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_521),
.B(n_233),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_525),
.B(n_392),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_534),
.B(n_190),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_526),
.B(n_238),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_639),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_534),
.B(n_190),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_562),
.B(n_434),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_537),
.B(n_264),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_629),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_557),
.B(n_550),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_563),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_532),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_586),
.B(n_191),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_639),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_654),
.B(n_191),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_629),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_639),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_599),
.A2(n_339),
.B1(n_275),
.B2(n_318),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_550),
.B(n_297),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_599),
.A2(n_597),
.B1(n_581),
.B2(n_574),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_540),
.A2(n_494),
.B(n_490),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_613),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_612),
.B(n_303),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_SL g693 ( 
.A(n_528),
.B(n_307),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_629),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_560),
.A2(n_194),
.B1(n_196),
.B2(n_198),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_657),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_624),
.B(n_194),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_657),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_658),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_638),
.B(n_310),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_632),
.B(n_196),
.Y(n_701)
);

BUFx5_ASAP7_75t_L g702 ( 
.A(n_543),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_650),
.B(n_312),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_632),
.B(n_322),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_SL g705 ( 
.A(n_561),
.B(n_512),
.Y(n_705)
);

BUFx4f_ASAP7_75t_L g706 ( 
.A(n_614),
.Y(n_706)
);

O2A1O1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_559),
.A2(n_492),
.B(n_328),
.C(n_352),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_657),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_601),
.B(n_258),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_603),
.B(n_329),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_583),
.B(n_198),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_624),
.B(n_201),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_601),
.B(n_187),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_603),
.B(n_334),
.Y(n_714)
);

OAI221xp5_ASAP7_75t_L g715 ( 
.A1(n_591),
.A2(n_335),
.B1(n_229),
.B2(n_354),
.C(n_224),
.Y(n_715)
);

NOR2xp67_ASAP7_75t_L g716 ( 
.A(n_583),
.B(n_549),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_601),
.B(n_258),
.Y(n_717)
);

NOR2xp67_ASAP7_75t_L g718 ( 
.A(n_555),
.B(n_492),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_640),
.B(n_201),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_616),
.B(n_494),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_616),
.B(n_209),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_578),
.B(n_209),
.Y(n_722)
);

OR2x6_ASAP7_75t_L g723 ( 
.A(n_601),
.B(n_325),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_578),
.B(n_210),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_619),
.B(n_210),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_656),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_581),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_580),
.B(n_325),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_585),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_585),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_619),
.B(n_211),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_527),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_578),
.B(n_269),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_553),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_579),
.B(n_269),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_527),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_658),
.Y(n_737)
);

OAI22x1_ASAP7_75t_SL g738 ( 
.A1(n_607),
.A2(n_192),
.B1(n_345),
.B2(n_341),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_579),
.B(n_333),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_579),
.B(n_643),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_542),
.A2(n_347),
.B1(n_346),
.B2(n_342),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_527),
.B(n_258),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_527),
.B(n_282),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_530),
.B(n_340),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_553),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_640),
.B(n_609),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_589),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_R g748 ( 
.A(n_561),
.B(n_340),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_522),
.B(n_342),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_524),
.B(n_346),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_597),
.A2(n_339),
.B1(n_350),
.B2(n_337),
.Y(n_751)
);

BUFx6f_ASAP7_75t_SL g752 ( 
.A(n_561),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_520),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_L g754 ( 
.A(n_531),
.B(n_339),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_538),
.B(n_339),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_539),
.B(n_339),
.Y(n_756)
);

INVx8_ASAP7_75t_L g757 ( 
.A(n_535),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_625),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_551),
.B(n_212),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_625),
.Y(n_760)
);

NOR3x1_ASAP7_75t_L g761 ( 
.A(n_618),
.B(n_544),
.C(n_643),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_520),
.Y(n_762)
);

BUFx6f_ASAP7_75t_SL g763 ( 
.A(n_614),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_552),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_554),
.B(n_239),
.Y(n_765)
);

NOR2xp67_ASAP7_75t_L g766 ( 
.A(n_577),
.B(n_59),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_558),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_531),
.B(n_242),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_560),
.A2(n_287),
.B1(n_244),
.B2(n_255),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_565),
.B(n_257),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_568),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_597),
.A2(n_350),
.B1(n_337),
.B2(n_336),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_590),
.B(n_262),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_520),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_SL g775 ( 
.A(n_596),
.B(n_282),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_598),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_609),
.B(n_272),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_610),
.B(n_277),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_540),
.A2(n_336),
.B1(n_188),
.B2(n_189),
.Y(n_779)
);

AND2x6_ASAP7_75t_SL g780 ( 
.A(n_580),
.B(n_187),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_617),
.B(n_63),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_620),
.B(n_284),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_589),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_535),
.B(n_188),
.Y(n_784)
);

NOR2xp67_ASAP7_75t_L g785 ( 
.A(n_628),
.B(n_137),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_535),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_560),
.A2(n_326),
.B1(n_324),
.B2(n_323),
.Y(n_787)
);

AND2x6_ASAP7_75t_SL g788 ( 
.A(n_580),
.B(n_189),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_627),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_535),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_637),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_580),
.A2(n_623),
.B1(n_621),
.B2(n_611),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_574),
.A2(n_652),
.B1(n_529),
.B2(n_536),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_656),
.Y(n_794)
);

NOR3xp33_ASAP7_75t_L g795 ( 
.A(n_544),
.B(n_316),
.C(n_314),
.Y(n_795)
);

BUFx5_ASAP7_75t_L g796 ( 
.A(n_531),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_644),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_649),
.B(n_528),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_528),
.B(n_313),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_594),
.B(n_311),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_644),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_646),
.Y(n_802)
);

OAI221xp5_ASAP7_75t_L g803 ( 
.A1(n_630),
.A2(n_308),
.B1(n_302),
.B2(n_301),
.C(n_296),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_645),
.B(n_268),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_574),
.A2(n_288),
.B1(n_286),
.B2(n_289),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_600),
.B(n_268),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_589),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_602),
.B(n_202),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_548),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_523),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_533),
.B(n_529),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_572),
.A2(n_618),
.B1(n_662),
.B2(n_531),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_533),
.B(n_197),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_533),
.B(n_197),
.Y(n_814)
);

AND2x6_ASAP7_75t_SL g815 ( 
.A(n_659),
.B(n_192),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_604),
.B(n_12),
.Y(n_816)
);

OAI22xp33_ASAP7_75t_L g817 ( 
.A1(n_626),
.A2(n_12),
.B1(n_13),
.B2(n_17),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_802),
.B(n_673),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_665),
.A2(n_536),
.B(n_529),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_746),
.B(n_604),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_746),
.A2(n_531),
.B1(n_529),
.B2(n_536),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_793),
.A2(n_536),
.B(n_604),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_793),
.A2(n_592),
.B1(n_523),
.B2(n_547),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_811),
.A2(n_653),
.B(n_636),
.Y(n_824)
);

BUFx4f_ASAP7_75t_L g825 ( 
.A(n_680),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_811),
.A2(n_653),
.B(n_636),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_670),
.B(n_547),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_798),
.A2(n_634),
.B(n_653),
.Y(n_828)
);

OAI21x1_ASAP7_75t_L g829 ( 
.A1(n_690),
.A2(n_664),
.B(n_592),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_690),
.A2(n_634),
.B(n_636),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_697),
.A2(n_652),
.B(n_655),
.C(n_660),
.Y(n_831)
);

AOI33xp33_ASAP7_75t_L g832 ( 
.A1(n_772),
.A2(n_593),
.A3(n_661),
.B1(n_651),
.B2(n_648),
.B3(n_642),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_809),
.Y(n_833)
);

NOR2x1_ASAP7_75t_L g834 ( 
.A(n_766),
.B(n_634),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_667),
.A2(n_605),
.B(n_661),
.C(n_651),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_682),
.B(n_556),
.Y(n_836)
);

OAI21xp33_ASAP7_75t_L g837 ( 
.A1(n_751),
.A2(n_605),
.B(n_648),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_689),
.A2(n_663),
.B1(n_642),
.B2(n_548),
.Y(n_838)
);

AOI21x1_ASAP7_75t_L g839 ( 
.A1(n_720),
.A2(n_663),
.B(n_567),
.Y(n_839)
);

NAND2x1p5_ASAP7_75t_L g840 ( 
.A(n_753),
.B(n_762),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_682),
.B(n_556),
.Y(n_841)
);

CKINVDCx14_ASAP7_75t_R g842 ( 
.A(n_726),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_797),
.B(n_556),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_672),
.B(n_556),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_678),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_689),
.A2(n_582),
.B(n_635),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_668),
.B(n_541),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_668),
.B(n_541),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_697),
.A2(n_587),
.B(n_635),
.C(n_633),
.Y(n_849)
);

AOI21x1_ASAP7_75t_L g850 ( 
.A1(n_679),
.A2(n_582),
.B(n_633),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_740),
.A2(n_576),
.B(n_541),
.Y(n_851)
);

OAI21x1_ASAP7_75t_L g852 ( 
.A1(n_729),
.A2(n_606),
.B(n_631),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_672),
.B(n_556),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_691),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_712),
.A2(n_584),
.B(n_622),
.C(n_571),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_711),
.B(n_569),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_712),
.A2(n_719),
.B(n_808),
.C(n_806),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_727),
.B(n_576),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_718),
.B(n_615),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_687),
.A2(n_575),
.B(n_567),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_677),
.A2(n_569),
.B(n_573),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_799),
.A2(n_569),
.B(n_573),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_671),
.B(n_573),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_806),
.B(n_564),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_688),
.A2(n_576),
.B(n_615),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_730),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_774),
.A2(n_615),
.B(n_566),
.Y(n_867)
);

AOI21x1_ASAP7_75t_L g868 ( 
.A1(n_693),
.A2(n_584),
.B(n_571),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_681),
.Y(n_869)
);

AO32x1_ASAP7_75t_L g870 ( 
.A1(n_764),
.A2(n_575),
.A3(n_588),
.B1(n_606),
.B2(n_608),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_774),
.A2(n_615),
.B(n_566),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_808),
.B(n_556),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_719),
.B(n_566),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_676),
.Y(n_874)
);

NOR2x1_ASAP7_75t_L g875 ( 
.A(n_785),
.B(n_608),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_681),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_685),
.B(n_694),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_681),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_767),
.Y(n_879)
);

NAND2x1_ASAP7_75t_L g880 ( 
.A(n_753),
.B(n_762),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_758),
.B(n_564),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_792),
.B(n_813),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_687),
.A2(n_595),
.B1(n_641),
.B2(n_564),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_744),
.A2(n_595),
.B(n_641),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_775),
.B(n_595),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_SL g886 ( 
.A(n_706),
.B(n_564),
.Y(n_886)
);

AO21x1_ASAP7_75t_L g887 ( 
.A1(n_816),
.A2(n_695),
.B(n_769),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_801),
.B(n_564),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_704),
.A2(n_641),
.B(n_531),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_804),
.B(n_13),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_814),
.B(n_641),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_771),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_760),
.B(n_17),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_666),
.A2(n_81),
.B1(n_167),
.B2(n_163),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_776),
.B(n_18),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_747),
.A2(n_80),
.B(n_162),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_789),
.B(n_18),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_783),
.A2(n_75),
.B(n_161),
.Y(n_898)
);

INVx3_ASAP7_75t_SL g899 ( 
.A(n_794),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_791),
.B(n_28),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_699),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_666),
.B(n_86),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_810),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_742),
.Y(n_904)
);

NOR3xp33_ASAP7_75t_L g905 ( 
.A(n_790),
.B(n_31),
.C(n_32),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_681),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_SL g907 ( 
.A(n_706),
.B(n_31),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_807),
.A2(n_90),
.B(n_159),
.Y(n_908)
);

NOR2x1_ASAP7_75t_L g909 ( 
.A(n_716),
.B(n_173),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_674),
.A2(n_147),
.B(n_139),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_692),
.B(n_700),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_675),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_790),
.B(n_38),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_703),
.B(n_39),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_812),
.A2(n_138),
.B1(n_136),
.B2(n_126),
.Y(n_915)
);

AOI21x1_ASAP7_75t_L g916 ( 
.A1(n_755),
.A2(n_125),
.B(n_121),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_745),
.B(n_43),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_734),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_734),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_710),
.B(n_714),
.Y(n_920)
);

AND2x6_ASAP7_75t_L g921 ( 
.A(n_761),
.B(n_781),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_683),
.A2(n_116),
.B(n_109),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_734),
.B(n_44),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_713),
.B(n_44),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_702),
.B(n_102),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_751),
.A2(n_779),
.B(n_772),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_709),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_669),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_669),
.A2(n_779),
.B1(n_762),
.B2(n_753),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_781),
.B(n_49),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_787),
.A2(n_54),
.B(n_756),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_805),
.A2(n_686),
.B(n_696),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_698),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_753),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_708),
.A2(n_707),
.B(n_765),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_784),
.B(n_732),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_715),
.A2(n_795),
.B(n_759),
.C(n_770),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_762),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_702),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_773),
.Y(n_940)
);

O2A1O1Ixp5_ASAP7_75t_L g941 ( 
.A1(n_800),
.A2(n_777),
.B(n_778),
.C(n_782),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_721),
.A2(n_731),
.B(n_725),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_702),
.Y(n_943)
);

INVx4_ASAP7_75t_L g944 ( 
.A(n_757),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_749),
.B(n_750),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_733),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_717),
.B(n_743),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_754),
.A2(n_701),
.B(n_739),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_733),
.B(n_741),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_786),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_684),
.B(n_724),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_722),
.B(n_735),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_736),
.A2(n_728),
.B1(n_757),
.B2(n_723),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_707),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_768),
.A2(n_796),
.B(n_757),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_723),
.A2(n_728),
.B(n_796),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_796),
.A2(n_728),
.B(n_803),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_796),
.A2(n_817),
.B(n_705),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_748),
.B(n_796),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_780),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_737),
.B(n_763),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_796),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_817),
.A2(n_738),
.B(n_748),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_788),
.B(n_815),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_763),
.B(n_752),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_665),
.A2(n_574),
.B(n_540),
.Y(n_966)
);

NAND3xp33_ASAP7_75t_L g967 ( 
.A(n_746),
.B(n_751),
.C(n_667),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_665),
.A2(n_574),
.B(n_540),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_665),
.A2(n_690),
.B(n_574),
.Y(n_969)
);

NAND3xp33_ASAP7_75t_L g970 ( 
.A(n_746),
.B(n_751),
.C(n_667),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_665),
.A2(n_574),
.B(n_540),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_793),
.A2(n_689),
.B1(n_665),
.B2(n_746),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_802),
.B(n_673),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_746),
.A2(n_667),
.B1(n_802),
.B2(n_673),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_802),
.B(n_673),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_746),
.A2(n_665),
.B(n_712),
.C(n_697),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_665),
.A2(n_574),
.B(n_540),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_681),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_793),
.A2(n_689),
.B1(n_665),
.B2(n_746),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_802),
.B(n_673),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_746),
.A2(n_667),
.B1(n_802),
.B2(n_673),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_668),
.B(n_563),
.Y(n_982)
);

OA22x2_ASAP7_75t_L g983 ( 
.A1(n_695),
.A2(n_580),
.B1(n_787),
.B2(n_769),
.Y(n_983)
);

NOR2xp67_ASAP7_75t_L g984 ( 
.A(n_680),
.B(n_654),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_802),
.B(n_673),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_802),
.B(n_673),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_802),
.B(n_673),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_746),
.B(n_654),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_678),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_976),
.A2(n_857),
.B(n_967),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_819),
.A2(n_839),
.B(n_850),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_852),
.A2(n_822),
.B(n_829),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_868),
.A2(n_969),
.B(n_968),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_830),
.A2(n_826),
.B(n_824),
.Y(n_994)
);

AOI21x1_ASAP7_75t_L g995 ( 
.A1(n_966),
.A2(n_977),
.B(n_971),
.Y(n_995)
);

AOI21x1_ASAP7_75t_L g996 ( 
.A1(n_820),
.A2(n_891),
.B(n_882),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_SL g997 ( 
.A1(n_972),
.A2(n_979),
.B(n_926),
.Y(n_997)
);

NOR2xp67_ASAP7_75t_L g998 ( 
.A(n_874),
.B(n_982),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_967),
.A2(n_970),
.B(n_974),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_818),
.B(n_973),
.Y(n_1000)
);

OA21x2_ASAP7_75t_L g1001 ( 
.A1(n_846),
.A2(n_932),
.B(n_855),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_846),
.A2(n_955),
.B(n_932),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_876),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_975),
.B(n_980),
.Y(n_1004)
);

INVx6_ASAP7_75t_L g1005 ( 
.A(n_944),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_854),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_842),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_862),
.A2(n_939),
.B(n_838),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_939),
.A2(n_828),
.B(n_823),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_988),
.A2(n_853),
.B(n_844),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_860),
.A2(n_865),
.B(n_851),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_920),
.A2(n_911),
.B(n_942),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_833),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_985),
.B(n_986),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_847),
.A2(n_848),
.B(n_861),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_860),
.A2(n_884),
.B(n_935),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_987),
.B(n_940),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_981),
.B(n_945),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_873),
.B(n_863),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_834),
.A2(n_821),
.B(n_948),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_854),
.Y(n_1021)
);

NOR2x1_ASAP7_75t_L g1022 ( 
.A(n_984),
.B(n_869),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_827),
.A2(n_859),
.B(n_841),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_892),
.B(n_930),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_876),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_935),
.A2(n_916),
.B(n_943),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_876),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_825),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_970),
.A2(n_926),
.B(n_937),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_836),
.A2(n_883),
.B(n_957),
.Y(n_1030)
);

AOI21x1_ASAP7_75t_L g1031 ( 
.A1(n_875),
.A2(n_864),
.B(n_872),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_929),
.A2(n_949),
.B1(n_952),
.B2(n_951),
.Y(n_1032)
);

AO31x2_ASAP7_75t_L g1033 ( 
.A1(n_887),
.A2(n_831),
.A3(n_849),
.B(n_954),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_928),
.A2(n_931),
.B(n_907),
.C(n_832),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_930),
.A2(n_858),
.B1(n_856),
.B2(n_983),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_845),
.Y(n_1036)
);

OR2x6_ASAP7_75t_L g1037 ( 
.A(n_901),
.B(n_965),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_835),
.A2(n_956),
.B(n_871),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_931),
.B(n_958),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_947),
.B(n_825),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_989),
.B(n_877),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_903),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_877),
.B(n_921),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_888),
.A2(n_904),
.B1(n_919),
.B2(n_978),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_867),
.A2(n_889),
.B(n_923),
.Y(n_1045)
);

OR2x6_ASAP7_75t_L g1046 ( 
.A(n_965),
.B(n_944),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_890),
.B(n_927),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_878),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_961),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_959),
.A2(n_843),
.B(n_925),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_921),
.B(n_914),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_837),
.A2(n_962),
.B(n_880),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_R g1053 ( 
.A(n_899),
.B(n_886),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_921),
.B(n_893),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_921),
.B(n_897),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_895),
.B(n_900),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_933),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_837),
.A2(n_902),
.B(n_886),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_918),
.A2(n_881),
.B(n_840),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_840),
.A2(n_941),
.B(n_934),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_866),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_924),
.B(n_946),
.Y(n_1062)
);

INVxp67_ASAP7_75t_SL g1063 ( 
.A(n_906),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_896),
.A2(n_908),
.B(n_898),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_910),
.A2(n_922),
.B(n_917),
.Y(n_1065)
);

INVx6_ASAP7_75t_L g1066 ( 
.A(n_906),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_961),
.B(n_936),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_909),
.A2(n_915),
.B(n_894),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_913),
.B(n_950),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_906),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_907),
.A2(n_912),
.B(n_963),
.C(n_905),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_953),
.A2(n_870),
.B(n_885),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_870),
.A2(n_938),
.B(n_978),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_938),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_938),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_964),
.B(n_960),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_960),
.A2(n_976),
.B(n_857),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_960),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_818),
.B(n_985),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_879),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_818),
.B(n_985),
.Y(n_1081)
);

AO21x1_ASAP7_75t_L g1082 ( 
.A1(n_972),
.A2(n_979),
.B(n_926),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_966),
.A2(n_793),
.B(n_574),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_818),
.B(n_985),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_854),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_982),
.B(n_671),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_854),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_976),
.B(n_972),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_818),
.B(n_985),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_818),
.B(n_985),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_L g1091 ( 
.A(n_857),
.B(n_982),
.C(n_668),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_854),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_854),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_819),
.A2(n_839),
.B(n_850),
.Y(n_1094)
);

AOI21xp33_ASAP7_75t_L g1095 ( 
.A1(n_982),
.A2(n_857),
.B(n_546),
.Y(n_1095)
);

INVxp67_ASAP7_75t_L g1096 ( 
.A(n_854),
.Y(n_1096)
);

AOI21x1_ASAP7_75t_L g1097 ( 
.A1(n_819),
.A2(n_968),
.B(n_966),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_818),
.B(n_985),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_L g1099 ( 
.A(n_976),
.B(n_972),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_982),
.B(n_671),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_819),
.A2(n_839),
.B(n_850),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_857),
.A2(n_982),
.B1(n_976),
.B2(n_979),
.Y(n_1102)
);

AOI221xp5_ASAP7_75t_SL g1103 ( 
.A1(n_926),
.A2(n_857),
.B1(n_928),
.B2(n_772),
.C(n_779),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_966),
.A2(n_793),
.B(n_574),
.Y(n_1104)
);

O2A1O1Ixp5_ASAP7_75t_L g1105 ( 
.A1(n_857),
.A2(n_976),
.B(n_882),
.C(n_665),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_818),
.B(n_985),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_976),
.A2(n_857),
.B(n_967),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_818),
.B(n_985),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_976),
.A2(n_857),
.B(n_967),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_876),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_966),
.A2(n_793),
.B(n_574),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_SL g1112 ( 
.A(n_857),
.B(n_563),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_842),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_818),
.B(n_985),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_819),
.A2(n_839),
.B(n_850),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_818),
.B(n_985),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_818),
.B(n_985),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_819),
.A2(n_839),
.B(n_850),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_854),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_818),
.B(n_985),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_966),
.A2(n_793),
.B(n_574),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_L g1122 ( 
.A(n_984),
.B(n_869),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_818),
.B(n_985),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_976),
.A2(n_857),
.B(n_967),
.Y(n_1124)
);

AO21x2_ASAP7_75t_L g1125 ( 
.A1(n_976),
.A2(n_969),
.B(n_665),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_966),
.A2(n_793),
.B(n_574),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_854),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_L g1128 ( 
.A(n_874),
.B(n_680),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_976),
.A2(n_979),
.A3(n_972),
.B(n_857),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_966),
.A2(n_793),
.B(n_574),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_819),
.A2(n_839),
.B(n_850),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_818),
.B(n_985),
.Y(n_1132)
);

AOI21x1_ASAP7_75t_L g1133 ( 
.A1(n_819),
.A2(n_968),
.B(n_966),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_966),
.A2(n_793),
.B(n_574),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_966),
.A2(n_793),
.B(n_574),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_819),
.A2(n_839),
.B(n_850),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1095),
.A2(n_1091),
.B(n_1102),
.C(n_1105),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1000),
.A2(n_1120),
.B1(n_1117),
.B2(n_1106),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1012),
.A2(n_1015),
.B(n_1083),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1080),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_1085),
.Y(n_1141)
);

AO22x1_ASAP7_75t_L g1142 ( 
.A1(n_1086),
.A2(n_1100),
.B1(n_1028),
.B2(n_1077),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1004),
.A2(n_1108),
.B1(n_1098),
.B2(n_1079),
.Y(n_1143)
);

BUFx4_ASAP7_75t_SL g1144 ( 
.A(n_1007),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1014),
.A2(n_1084),
.B1(n_1123),
.B2(n_1081),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_1007),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1082),
.A2(n_1099),
.B1(n_1112),
.B2(n_1088),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1089),
.B(n_1090),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1047),
.B(n_1040),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1114),
.B(n_1116),
.Y(n_1150)
);

NOR2xp67_ASAP7_75t_R g1151 ( 
.A(n_1005),
.B(n_1013),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_1046),
.B(n_1037),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_998),
.B(n_1017),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1099),
.A2(n_1103),
.B1(n_1132),
.B2(n_1018),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1069),
.B(n_1092),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1036),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1019),
.B(n_1056),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1092),
.B(n_1087),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1062),
.B(n_1032),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1104),
.A2(n_1121),
.B(n_1135),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1111),
.A2(n_1134),
.B(n_1130),
.Y(n_1161)
);

INVx3_ASAP7_75t_SL g1162 ( 
.A(n_1113),
.Y(n_1162)
);

INVx3_ASAP7_75t_SL g1163 ( 
.A(n_1113),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1024),
.B(n_999),
.Y(n_1164)
);

AND2x6_ASAP7_75t_L g1165 ( 
.A(n_1043),
.B(n_1051),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1126),
.A2(n_1030),
.B(n_1020),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1046),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1105),
.A2(n_997),
.B(n_1029),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1034),
.A2(n_1088),
.B1(n_990),
.B2(n_1107),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_1093),
.Y(n_1170)
);

OA21x2_ASAP7_75t_L g1171 ( 
.A1(n_993),
.A2(n_1026),
.B(n_1002),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1006),
.B(n_1021),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1039),
.A2(n_1023),
.B(n_1058),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1041),
.B(n_1034),
.Y(n_1174)
);

INVx3_ASAP7_75t_SL g1175 ( 
.A(n_1037),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1109),
.A2(n_1124),
.B1(n_1071),
.B2(n_1035),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1096),
.B(n_1119),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1125),
.A2(n_1071),
.B1(n_1054),
.B2(n_1055),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1042),
.B(n_1096),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1046),
.B(n_1037),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1060),
.A2(n_1052),
.A3(n_1050),
.B(n_1044),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1127),
.B(n_1129),
.Y(n_1182)
);

OAI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_1053),
.A2(n_1067),
.B(n_1076),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1049),
.B(n_1122),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1078),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1022),
.B(n_1061),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1002),
.A2(n_994),
.B(n_1009),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1053),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1078),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1128),
.B(n_1057),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1074),
.B(n_1075),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1009),
.A2(n_1011),
.B(n_1008),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1068),
.A2(n_1016),
.B(n_1072),
.C(n_1059),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1070),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_1003),
.Y(n_1195)
);

INVx5_ASAP7_75t_L g1196 ( 
.A(n_1005),
.Y(n_1196)
);

O2A1O1Ixp5_ASAP7_75t_L g1197 ( 
.A1(n_1031),
.A2(n_995),
.B(n_1133),
.C(n_1097),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1001),
.A2(n_1063),
.B1(n_1016),
.B2(n_1072),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1003),
.Y(n_1199)
);

AO21x2_ASAP7_75t_L g1200 ( 
.A1(n_993),
.A2(n_992),
.B(n_991),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1066),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_1066),
.B(n_1048),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1129),
.B(n_1033),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1025),
.Y(n_1204)
);

INVx3_ASAP7_75t_SL g1205 ( 
.A(n_1025),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1027),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1011),
.A2(n_1008),
.B(n_1038),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1038),
.A2(n_1065),
.B(n_1064),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1033),
.B(n_1110),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_996),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_1073),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1010),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1033),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1065),
.B(n_991),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1064),
.A2(n_992),
.B(n_1045),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1094),
.A2(n_1101),
.B1(n_1115),
.B2(n_1118),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1136),
.A2(n_1091),
.B1(n_857),
.B2(n_982),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1118),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1131),
.B(n_1000),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_1046),
.B(n_1037),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1012),
.A2(n_968),
.B(n_966),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1085),
.Y(n_1222)
);

NAND2x1p5_ASAP7_75t_L g1223 ( 
.A(n_1006),
.B(n_854),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1000),
.B(n_1004),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1102),
.A2(n_926),
.B1(n_1004),
.B2(n_1000),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1095),
.B(n_982),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1080),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1092),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1046),
.B(n_944),
.Y(n_1229)
);

CKINVDCx6p67_ASAP7_75t_R g1230 ( 
.A(n_1078),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1085),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1046),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1046),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1012),
.A2(n_968),
.B(n_966),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1085),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1105),
.A2(n_976),
.B(n_997),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1046),
.Y(n_1237)
);

INVx8_ASAP7_75t_L g1238 ( 
.A(n_1046),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1000),
.B(n_1004),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1012),
.A2(n_968),
.B(n_966),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1000),
.B(n_1004),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1086),
.B(n_1100),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1085),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1085),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1086),
.B(n_1100),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1085),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1005),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1000),
.B(n_1004),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1000),
.B(n_1004),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1080),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1105),
.A2(n_976),
.B(n_997),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1046),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1017),
.B(n_737),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1046),
.B(n_1037),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1092),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1046),
.B(n_944),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1005),
.Y(n_1257)
);

AO21x2_ASAP7_75t_L g1258 ( 
.A1(n_1029),
.A2(n_1107),
.B(n_990),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1017),
.B(n_737),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1086),
.B(n_1100),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1085),
.Y(n_1261)
);

BUFx12f_ASAP7_75t_L g1262 ( 
.A(n_1113),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1046),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1000),
.B(n_1004),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_1005),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1102),
.A2(n_926),
.B1(n_1004),
.B2(n_1000),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1046),
.B(n_944),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1000),
.B(n_1004),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1086),
.B(n_1100),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1046),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1085),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1091),
.A2(n_857),
.B1(n_982),
.B2(n_1102),
.Y(n_1272)
);

INVxp67_ASAP7_75t_L g1273 ( 
.A(n_1092),
.Y(n_1273)
);

NOR2xp67_ASAP7_75t_SL g1274 ( 
.A(n_1078),
.B(n_680),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1092),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1229),
.B(n_1256),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1148),
.B(n_1150),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1208),
.A2(n_1215),
.B(n_1207),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1196),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1226),
.A2(n_1272),
.B(n_1159),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1197),
.A2(n_1166),
.B(n_1192),
.Y(n_1281)
);

BUFx12f_ASAP7_75t_L g1282 ( 
.A(n_1262),
.Y(n_1282)
);

BUFx4f_ASAP7_75t_L g1283 ( 
.A(n_1238),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1185),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1224),
.B(n_1239),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1187),
.A2(n_1216),
.B(n_1161),
.Y(n_1286)
);

OAI21xp33_ASAP7_75t_L g1287 ( 
.A1(n_1272),
.A2(n_1248),
.B(n_1241),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1141),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1227),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1160),
.A2(n_1139),
.B(n_1173),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1176),
.A2(n_1169),
.B1(n_1258),
.B2(n_1225),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1170),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1183),
.A2(n_1260),
.B1(n_1242),
.B2(n_1269),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1228),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1236),
.A2(n_1251),
.B(n_1234),
.Y(n_1295)
);

CKINVDCx6p67_ASAP7_75t_R g1296 ( 
.A(n_1162),
.Y(n_1296)
);

OAI21xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1249),
.A2(n_1268),
.B(n_1264),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1196),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1189),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1245),
.A2(n_1153),
.B1(n_1138),
.B2(n_1143),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1146),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1143),
.B(n_1145),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1238),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1202),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1214),
.A2(n_1221),
.B(n_1240),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_1172),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1156),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1229),
.B(n_1256),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1236),
.A2(n_1251),
.B(n_1193),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1176),
.A2(n_1258),
.B1(n_1225),
.B2(n_1266),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1266),
.A2(n_1147),
.B1(n_1168),
.B2(n_1145),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1141),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1250),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1157),
.A2(n_1188),
.B1(n_1253),
.B2(n_1259),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1267),
.B(n_1180),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1158),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1179),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1182),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_1202),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1244),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1168),
.A2(n_1137),
.B(n_1217),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1194),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1155),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1164),
.A2(n_1154),
.B1(n_1174),
.B2(n_1217),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1154),
.B(n_1178),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1199),
.Y(n_1326)
);

BUFx2_ASAP7_75t_SL g1327 ( 
.A(n_1222),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1218),
.A2(n_1198),
.B(n_1219),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1209),
.Y(n_1329)
);

BUFx2_ASAP7_75t_SL g1330 ( 
.A(n_1231),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1171),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1195),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1191),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1181),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1267),
.B(n_1180),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1178),
.A2(n_1165),
.B1(n_1149),
.B2(n_1255),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1191),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1200),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1265),
.B(n_1252),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1200),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1275),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1165),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1213),
.B(n_1203),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1165),
.A2(n_1273),
.B1(n_1177),
.B2(n_1190),
.Y(n_1344)
);

BUFx2_ASAP7_75t_R g1345 ( 
.A(n_1163),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1235),
.B(n_1271),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1223),
.A2(n_1210),
.B1(n_1212),
.B2(n_1261),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1186),
.Y(n_1348)
);

BUFx4f_ASAP7_75t_SL g1349 ( 
.A(n_1230),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1243),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1246),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1165),
.A2(n_1184),
.B1(n_1270),
.B2(n_1232),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1184),
.A2(n_1186),
.B1(n_1270),
.B2(n_1237),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1274),
.B(n_1205),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1151),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_SL g1356 ( 
.A(n_1175),
.B(n_1270),
.Y(n_1356)
);

INVx6_ASAP7_75t_L g1357 ( 
.A(n_1202),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1206),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1167),
.A2(n_1263),
.B1(n_1252),
.B2(n_1237),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1167),
.A2(n_1263),
.B1(n_1237),
.B2(n_1233),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1211),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1206),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1151),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1233),
.Y(n_1364)
);

INVx5_ASAP7_75t_SL g1365 ( 
.A(n_1152),
.Y(n_1365)
);

AOI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1152),
.A2(n_1220),
.B(n_1254),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1144),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1206),
.Y(n_1368)
);

AOI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1152),
.A2(n_1220),
.B(n_1254),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1204),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1220),
.Y(n_1371)
);

BUFx2_ASAP7_75t_R g1372 ( 
.A(n_1247),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1233),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1252),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1254),
.A2(n_1263),
.B1(n_1257),
.B2(n_1201),
.Y(n_1375)
);

OR2x6_ASAP7_75t_L g1376 ( 
.A(n_1142),
.B(n_997),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1226),
.A2(n_1095),
.B1(n_926),
.B2(n_1091),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1140),
.Y(n_1378)
);

BUFx8_ASAP7_75t_L g1379 ( 
.A(n_1188),
.Y(n_1379)
);

BUFx4f_ASAP7_75t_SL g1380 ( 
.A(n_1170),
.Y(n_1380)
);

CKINVDCx11_ASAP7_75t_R g1381 ( 
.A(n_1146),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1272),
.B(n_1077),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1226),
.A2(n_1095),
.B1(n_926),
.B2(n_1091),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1272),
.B(n_1077),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1331),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1278),
.A2(n_1286),
.B(n_1305),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1338),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1280),
.B(n_1302),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_1288),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1338),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1329),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1318),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1340),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_1301),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1361),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1366),
.B(n_1369),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1343),
.B(n_1321),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1325),
.B(n_1382),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1342),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1294),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1294),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1287),
.B(n_1382),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1328),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1316),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1384),
.B(n_1321),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1323),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1290),
.A2(n_1309),
.B(n_1384),
.Y(n_1407)
);

OAI21xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1311),
.A2(n_1291),
.B(n_1377),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1281),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1321),
.Y(n_1410)
);

AOI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1376),
.A2(n_1342),
.B(n_1295),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1291),
.B(n_1310),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1297),
.B(n_1324),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1324),
.B(n_1277),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1334),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1309),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1309),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1295),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1283),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1295),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1310),
.B(n_1311),
.Y(n_1421)
);

AOI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1376),
.A2(n_1363),
.B(n_1355),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1307),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1313),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1377),
.A2(n_1383),
.B(n_1336),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1383),
.B(n_1300),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1376),
.B(n_1336),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1371),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1381),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1376),
.B(n_1326),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1320),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1371),
.Y(n_1432)
);

INVxp33_ASAP7_75t_L g1433 ( 
.A(n_1346),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1365),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1285),
.B(n_1317),
.Y(n_1435)
);

CKINVDCx12_ASAP7_75t_R g1436 ( 
.A(n_1372),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1357),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1322),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1283),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_1301),
.Y(n_1440)
);

AO21x2_ASAP7_75t_L g1441 ( 
.A1(n_1375),
.A2(n_1348),
.B(n_1314),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1344),
.B(n_1347),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1289),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1357),
.Y(n_1444)
);

AO21x2_ASAP7_75t_L g1445 ( 
.A1(n_1293),
.A2(n_1378),
.B(n_1373),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1312),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1365),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1332),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1341),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1365),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1365),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1352),
.B(n_1353),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1304),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1403),
.Y(n_1454)
);

INVxp67_ASAP7_75t_SL g1455 ( 
.A(n_1410),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1430),
.B(n_1303),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1426),
.A2(n_1379),
.B1(n_1335),
.B2(n_1315),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1405),
.B(n_1374),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1400),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1426),
.A2(n_1379),
.B1(n_1335),
.B2(n_1315),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1401),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1421),
.A2(n_1306),
.B1(n_1357),
.B2(n_1359),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1398),
.B(n_1397),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1396),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1407),
.B(n_1368),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1424),
.B(n_1370),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1424),
.B(n_1370),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1427),
.B(n_1276),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_1404),
.Y(n_1469)
);

OAI221xp5_ASAP7_75t_L g1470 ( 
.A1(n_1408),
.A2(n_1356),
.B1(n_1360),
.B2(n_1354),
.C(n_1333),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1430),
.B(n_1364),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1407),
.B(n_1337),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1399),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1407),
.B(n_1351),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1388),
.B(n_1364),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1407),
.B(n_1276),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1417),
.B(n_1350),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1416),
.B(n_1308),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_1394),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1416),
.B(n_1308),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1422),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1385),
.B(n_1308),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1388),
.B(n_1364),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1423),
.B(n_1319),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1391),
.B(n_1319),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1418),
.B(n_1330),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1418),
.B(n_1327),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1391),
.B(n_1362),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1412),
.B(n_1358),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_L g1490 ( 
.A(n_1413),
.B(n_1379),
.C(n_1381),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1418),
.B(n_1420),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1420),
.B(n_1339),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1463),
.B(n_1411),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1490),
.B(n_1414),
.Y(n_1494)
);

NAND3xp33_ASAP7_75t_L g1495 ( 
.A(n_1490),
.B(n_1413),
.C(n_1408),
.Y(n_1495)
);

NAND3xp33_ASAP7_75t_L g1496 ( 
.A(n_1462),
.B(n_1414),
.C(n_1435),
.Y(n_1496)
);

NAND4xp25_ASAP7_75t_L g1497 ( 
.A(n_1470),
.B(n_1435),
.C(n_1402),
.D(n_1421),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1469),
.B(n_1438),
.Y(n_1498)
);

NAND4xp25_ASAP7_75t_SL g1499 ( 
.A(n_1470),
.B(n_1442),
.C(n_1402),
.D(n_1412),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1463),
.B(n_1411),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1458),
.B(n_1476),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1474),
.B(n_1392),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1458),
.B(n_1415),
.Y(n_1503)
);

NAND4xp25_ASAP7_75t_L g1504 ( 
.A(n_1462),
.B(n_1389),
.C(n_1483),
.D(n_1475),
.Y(n_1504)
);

OAI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1457),
.A2(n_1442),
.B1(n_1452),
.B2(n_1292),
.C(n_1367),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1458),
.B(n_1399),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1469),
.B(n_1406),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1456),
.B(n_1437),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1474),
.B(n_1395),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1459),
.B(n_1431),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1459),
.B(n_1448),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1481),
.A2(n_1425),
.B(n_1419),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_L g1513 ( 
.A(n_1461),
.B(n_1449),
.C(n_1446),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1483),
.B(n_1445),
.Y(n_1514)
);

AND2x2_ASAP7_75t_SL g1515 ( 
.A(n_1481),
.B(n_1425),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1479),
.B(n_1433),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1461),
.B(n_1445),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1466),
.B(n_1445),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1476),
.B(n_1387),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1476),
.B(n_1387),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1460),
.A2(n_1436),
.B1(n_1440),
.B2(n_1425),
.Y(n_1521)
);

NAND3xp33_ASAP7_75t_L g1522 ( 
.A(n_1477),
.B(n_1425),
.C(n_1453),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1456),
.A2(n_1441),
.B1(n_1489),
.B2(n_1452),
.Y(n_1523)
);

OAI221xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1486),
.A2(n_1296),
.B1(n_1450),
.B2(n_1451),
.C(n_1428),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1478),
.B(n_1387),
.Y(n_1525)
);

OAI221xp5_ASAP7_75t_L g1526 ( 
.A1(n_1464),
.A2(n_1451),
.B1(n_1450),
.B2(n_1429),
.C(n_1447),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1478),
.B(n_1390),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1466),
.B(n_1467),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1467),
.B(n_1484),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1480),
.B(n_1390),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1484),
.B(n_1445),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_SL g1532 ( 
.A1(n_1468),
.A2(n_1396),
.B(n_1436),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1465),
.B(n_1393),
.Y(n_1533)
);

NOR3xp33_ASAP7_75t_L g1534 ( 
.A(n_1488),
.B(n_1422),
.C(n_1434),
.Y(n_1534)
);

OA21x2_ASAP7_75t_L g1535 ( 
.A1(n_1455),
.A2(n_1386),
.B(n_1409),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1485),
.B(n_1443),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_1456),
.B(n_1444),
.Y(n_1537)
);

OAI221xp5_ASAP7_75t_SL g1538 ( 
.A1(n_1486),
.A2(n_1296),
.B1(n_1432),
.B2(n_1428),
.C(n_1447),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1510),
.B(n_1482),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1501),
.B(n_1464),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1501),
.B(n_1464),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1502),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1493),
.B(n_1465),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1498),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1531),
.B(n_1518),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1493),
.B(n_1465),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1502),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1509),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1500),
.B(n_1472),
.Y(n_1549)
);

AND2x6_ASAP7_75t_SL g1550 ( 
.A(n_1516),
.B(n_1282),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1508),
.B(n_1487),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1537),
.B(n_1471),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1514),
.B(n_1473),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1519),
.B(n_1472),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1533),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1533),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1509),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1519),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1520),
.B(n_1503),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1520),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1529),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1536),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1535),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1525),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1525),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1503),
.B(n_1472),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1528),
.Y(n_1567)
);

INVx4_ASAP7_75t_L g1568 ( 
.A(n_1535),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1506),
.B(n_1492),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1506),
.B(n_1492),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1507),
.Y(n_1571)
);

INVxp67_ASAP7_75t_SL g1572 ( 
.A(n_1513),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1517),
.B(n_1491),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1522),
.B(n_1454),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1549),
.B(n_1515),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1545),
.B(n_1553),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1549),
.B(n_1515),
.Y(n_1577)
);

AND2x4_ASAP7_75t_SL g1578 ( 
.A(n_1552),
.B(n_1534),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1563),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1558),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1572),
.B(n_1513),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1545),
.B(n_1522),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1558),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1543),
.B(n_1515),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1543),
.B(n_1527),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1568),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1571),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1544),
.B(n_1511),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1555),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1556),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1568),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1544),
.B(n_1523),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1557),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1553),
.B(n_1527),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1546),
.B(n_1530),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1557),
.Y(n_1596)
);

INVxp33_ASAP7_75t_L g1597 ( 
.A(n_1539),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1542),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1563),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1554),
.B(n_1566),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1551),
.A2(n_1495),
.B1(n_1499),
.B2(n_1521),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1566),
.B(n_1540),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1547),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1562),
.B(n_1561),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1551),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1564),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_1551),
.Y(n_1607)
);

OAI21xp33_ASAP7_75t_L g1608 ( 
.A1(n_1574),
.A2(n_1495),
.B(n_1497),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1578),
.B(n_1540),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1601),
.A2(n_1494),
.B(n_1496),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1593),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1578),
.B(n_1541),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1607),
.B(n_1574),
.Y(n_1613)
);

NAND3xp33_ASAP7_75t_SL g1614 ( 
.A(n_1601),
.B(n_1496),
.C(n_1505),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1575),
.B(n_1541),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1608),
.B(n_1581),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1578),
.B(n_1560),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1593),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1608),
.B(n_1548),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1598),
.B(n_1567),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1598),
.B(n_1573),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1596),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1579),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1579),
.Y(n_1624)
);

NAND4xp75_ASAP7_75t_L g1625 ( 
.A(n_1592),
.B(n_1439),
.C(n_1419),
.D(n_1550),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1575),
.B(n_1559),
.Y(n_1626)
);

INVxp67_ASAP7_75t_SL g1627 ( 
.A(n_1579),
.Y(n_1627)
);

NOR2xp67_ASAP7_75t_L g1628 ( 
.A(n_1582),
.B(n_1568),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1577),
.B(n_1569),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_SL g1630 ( 
.A(n_1587),
.B(n_1526),
.C(n_1532),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1599),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1596),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1603),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1603),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1577),
.B(n_1559),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1599),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1580),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1580),
.Y(n_1638)
);

INVx2_ASAP7_75t_SL g1639 ( 
.A(n_1607),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1584),
.B(n_1564),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1597),
.B(n_1282),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1599),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1586),
.Y(n_1643)
);

NOR2xp67_ASAP7_75t_L g1644 ( 
.A(n_1582),
.B(n_1532),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1583),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1588),
.B(n_1345),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1584),
.B(n_1569),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1600),
.B(n_1570),
.Y(n_1648)
);

OR2x6_ASAP7_75t_L g1649 ( 
.A(n_1605),
.B(n_1512),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1602),
.B(n_1565),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1637),
.Y(n_1651)
);

NOR2x1p5_ASAP7_75t_L g1652 ( 
.A(n_1614),
.B(n_1504),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1639),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1637),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1638),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1619),
.B(n_1576),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1639),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1639),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_SL g1659 ( 
.A(n_1625),
.B(n_1524),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1619),
.B(n_1576),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1616),
.B(n_1610),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1623),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1638),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1621),
.B(n_1594),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1625),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1645),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1645),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1616),
.B(n_1604),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1610),
.B(n_1602),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1644),
.A2(n_1538),
.B1(n_1521),
.B2(n_1512),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1626),
.B(n_1635),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1623),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1626),
.B(n_1585),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1611),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1626),
.B(n_1635),
.Y(n_1675)
);

NAND3xp33_ASAP7_75t_L g1676 ( 
.A(n_1644),
.B(n_1504),
.C(n_1497),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1617),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1635),
.B(n_1585),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1623),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1614),
.A2(n_1396),
.B1(n_1441),
.B2(n_1471),
.Y(n_1680)
);

AND2x4_ASAP7_75t_SL g1681 ( 
.A(n_1617),
.B(n_1552),
.Y(n_1681)
);

NAND2x1p5_ASAP7_75t_L g1682 ( 
.A(n_1628),
.B(n_1481),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1609),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1609),
.B(n_1595),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1613),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1617),
.Y(n_1686)
);

NOR3xp33_ASAP7_75t_L g1687 ( 
.A(n_1661),
.B(n_1630),
.C(n_1641),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1652),
.A2(n_1630),
.B1(n_1609),
.B2(n_1612),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1657),
.Y(n_1689)
);

A2O1A1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1652),
.A2(n_1646),
.B(n_1628),
.C(n_1613),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1658),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1685),
.Y(n_1692)
);

OAI322xp33_ASAP7_75t_L g1693 ( 
.A1(n_1659),
.A2(n_1634),
.A3(n_1633),
.B1(n_1618),
.B2(n_1622),
.C1(n_1611),
.C2(n_1632),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1656),
.B(n_1621),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1651),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1671),
.B(n_1629),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1685),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1653),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1656),
.B(n_1620),
.Y(n_1699)
);

OAI32xp33_ASAP7_75t_L g1700 ( 
.A1(n_1665),
.A2(n_1612),
.A3(n_1633),
.B1(n_1634),
.B2(n_1620),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1676),
.A2(n_1612),
.B1(n_1649),
.B2(n_1613),
.Y(n_1701)
);

O2A1O1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1676),
.A2(n_1649),
.B(n_1613),
.C(n_1643),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1653),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1677),
.B(n_1629),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1671),
.B(n_1647),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1651),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1675),
.B(n_1647),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1654),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1675),
.B(n_1648),
.Y(n_1709)
);

CKINVDCx14_ASAP7_75t_R g1710 ( 
.A(n_1670),
.Y(n_1710)
);

AOI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1680),
.A2(n_1643),
.B1(n_1618),
.B2(n_1622),
.C(n_1632),
.Y(n_1711)
);

NAND3xp33_ASAP7_75t_L g1712 ( 
.A(n_1668),
.B(n_1643),
.C(n_1649),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1692),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1696),
.B(n_1686),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1705),
.B(n_1683),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1689),
.B(n_1669),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1691),
.B(n_1683),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1707),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1692),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1697),
.B(n_1684),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1687),
.B(n_1684),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1688),
.B(n_1653),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1709),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1687),
.B(n_1673),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1704),
.Y(n_1725)
);

AOI222xp33_ASAP7_75t_L g1726 ( 
.A1(n_1711),
.A2(n_1681),
.B1(n_1678),
.B2(n_1673),
.C1(n_1655),
.C2(n_1663),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_R g1727 ( 
.A(n_1710),
.B(n_1349),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1698),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1690),
.B(n_1678),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1702),
.B(n_1660),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1693),
.A2(n_1660),
.B1(n_1674),
.B2(n_1663),
.C(n_1654),
.Y(n_1731)
);

NAND2x1_ASAP7_75t_L g1732 ( 
.A(n_1701),
.B(n_1649),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1730),
.A2(n_1712),
.B1(n_1681),
.B2(n_1694),
.Y(n_1733)
);

AOI21xp33_ASAP7_75t_SL g1734 ( 
.A1(n_1730),
.A2(n_1729),
.B(n_1721),
.Y(n_1734)
);

AOI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1722),
.A2(n_1690),
.B(n_1700),
.Y(n_1735)
);

AOI211xp5_ASAP7_75t_L g1736 ( 
.A1(n_1722),
.A2(n_1698),
.B(n_1703),
.C(n_1699),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1719),
.Y(n_1737)
);

AOI221x1_ASAP7_75t_L g1738 ( 
.A1(n_1713),
.A2(n_1708),
.B1(n_1706),
.B2(n_1695),
.C(n_1655),
.Y(n_1738)
);

AOI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1724),
.A2(n_1703),
.B1(n_1666),
.B2(n_1667),
.C(n_1674),
.Y(n_1739)
);

AOI211xp5_ASAP7_75t_L g1740 ( 
.A1(n_1727),
.A2(n_1667),
.B(n_1666),
.C(n_1664),
.Y(n_1740)
);

AOI211xp5_ASAP7_75t_L g1741 ( 
.A1(n_1727),
.A2(n_1664),
.B(n_1662),
.C(n_1672),
.Y(n_1741)
);

AOI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1731),
.A2(n_1681),
.B1(n_1662),
.B2(n_1679),
.C(n_1672),
.Y(n_1742)
);

AOI211xp5_ASAP7_75t_SL g1743 ( 
.A1(n_1719),
.A2(n_1380),
.B(n_1679),
.C(n_1672),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1715),
.B(n_1615),
.Y(n_1744)
);

AOI211xp5_ASAP7_75t_SL g1745 ( 
.A1(n_1735),
.A2(n_1728),
.B(n_1717),
.C(n_1725),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1737),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1736),
.B(n_1718),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1742),
.A2(n_1714),
.B1(n_1726),
.B2(n_1723),
.Y(n_1748)
);

NOR3xp33_ASAP7_75t_L g1749 ( 
.A(n_1734),
.B(n_1716),
.C(n_1732),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1738),
.Y(n_1750)
);

NAND3x1_ASAP7_75t_L g1751 ( 
.A(n_1739),
.B(n_1720),
.C(n_1640),
.Y(n_1751)
);

NOR3xp33_ASAP7_75t_L g1752 ( 
.A(n_1740),
.B(n_1679),
.C(n_1662),
.Y(n_1752)
);

NOR3xp33_ASAP7_75t_L g1753 ( 
.A(n_1741),
.B(n_1744),
.C(n_1743),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1733),
.B(n_1682),
.Y(n_1754)
);

NOR2x1_ASAP7_75t_L g1755 ( 
.A(n_1750),
.B(n_1649),
.Y(n_1755)
);

NOR4xp25_ASAP7_75t_L g1756 ( 
.A(n_1747),
.B(n_1642),
.C(n_1631),
.D(n_1636),
.Y(n_1756)
);

NAND5xp2_ASAP7_75t_L g1757 ( 
.A(n_1745),
.B(n_1682),
.C(n_1640),
.D(n_1627),
.E(n_1615),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1746),
.Y(n_1758)
);

NAND3xp33_ASAP7_75t_SL g1759 ( 
.A(n_1749),
.B(n_1753),
.C(n_1748),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1754),
.B(n_1752),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1758),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1759),
.A2(n_1751),
.B1(n_1649),
.B2(n_1682),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1760),
.B(n_1640),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1755),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1756),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1757),
.B(n_1650),
.Y(n_1766)
);

OAI21xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1762),
.A2(n_1631),
.B(n_1624),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_R g1768 ( 
.A1(n_1765),
.A2(n_1642),
.B1(n_1624),
.B2(n_1636),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1763),
.B(n_1627),
.Y(n_1769)
);

AOI221xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1764),
.A2(n_1624),
.B1(n_1642),
.B2(n_1636),
.C(n_1631),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1761),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1769),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1771),
.B(n_1766),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1768),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1773),
.Y(n_1775)
);

AOI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1775),
.A2(n_1774),
.B1(n_1767),
.B2(n_1773),
.C(n_1772),
.Y(n_1776)
);

OA22x2_ASAP7_75t_L g1777 ( 
.A1(n_1776),
.A2(n_1770),
.B1(n_1591),
.B2(n_1586),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1776),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1777),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1778),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1780),
.A2(n_1591),
.B1(n_1284),
.B2(n_1299),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_R g1782 ( 
.A(n_1781),
.B(n_1779),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1782),
.A2(n_1284),
.B1(n_1299),
.B2(n_1650),
.Y(n_1783)
);

AOI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1783),
.A2(n_1589),
.B1(n_1583),
.B2(n_1606),
.C(n_1590),
.Y(n_1784)
);

AOI211xp5_ASAP7_75t_L g1785 ( 
.A1(n_1784),
.A2(n_1279),
.B(n_1298),
.C(n_1428),
.Y(n_1785)
);


endmodule