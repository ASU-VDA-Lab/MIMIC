module fake_jpeg_9110_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_2),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_4),
.B(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_17),
.B(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_4),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_12),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_1),
.B1(n_3),
.B2(n_13),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_14),
.B1(n_10),
.B2(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_18),
.C(n_12),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_27),
.B1(n_20),
.B2(n_19),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_14),
.B1(n_8),
.B2(n_11),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_26),
.B1(n_30),
.B2(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_16),
.C(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_32),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_24),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_38),
.C(n_39),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_16),
.B(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_8),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_16),
.B1(n_34),
.B2(n_15),
.Y(n_42)
);

NOR5xp2_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_43),
.C(n_15),
.D(n_7),
.E(n_3),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_8),
.B(n_15),
.C(n_1),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_43),
.B1(n_41),
.B2(n_3),
.Y(n_45)
);


endmodule