module fake_jpeg_13729_n_568 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_568);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_568;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_6),
.B(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

HAxp5_ASAP7_75t_SL g57 ( 
.A(n_27),
.B(n_0),
.CON(n_57),
.SN(n_57)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_57),
.B(n_106),
.Y(n_150)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_109),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_63),
.Y(n_171)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g132 ( 
.A(n_65),
.Y(n_132)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_9),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_68),
.B(n_80),
.Y(n_144)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_69),
.Y(n_136)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_73),
.Y(n_163)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_29),
.B(n_9),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_77),
.B(n_82),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_29),
.B(n_9),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_33),
.B(n_45),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_81),
.B(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_33),
.B(n_16),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_87),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_23),
.Y(n_95)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_98),
.Y(n_178)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_43),
.B(n_8),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

BUFx4f_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_27),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

CKINVDCx6p67_ASAP7_75t_R g211 ( 
.A(n_113),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_55),
.A2(n_28),
.B1(n_42),
.B2(n_48),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_115),
.A2(n_134),
.B1(n_158),
.B2(n_27),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_41),
.C(n_36),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_122),
.B(n_159),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_45),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_123),
.B(n_142),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_48),
.B1(n_44),
.B2(n_42),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_124),
.A2(n_149),
.B1(n_35),
.B2(n_50),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_54),
.A2(n_28),
.B1(n_44),
.B2(n_48),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_87),
.B(n_43),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_56),
.A2(n_48),
.B1(n_44),
.B2(n_42),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_86),
.B(n_41),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_154),
.B(n_157),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_91),
.B(n_51),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_95),
.A2(n_20),
.B1(n_31),
.B2(n_57),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_71),
.B(n_51),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_79),
.B(n_40),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_167),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_60),
.B(n_40),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_63),
.B(n_32),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_31),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_58),
.B(n_32),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_176),
.Y(n_185)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

BUFx2_ASAP7_75t_SL g210 ( 
.A(n_175),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_75),
.B(n_53),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_103),
.B(n_27),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_177),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_180),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_139),
.A2(n_73),
.B1(n_105),
.B2(n_94),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_181),
.A2(n_196),
.B1(n_203),
.B2(n_213),
.Y(n_290)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_184),
.Y(n_261)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_186),
.Y(n_283)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_189),
.Y(n_281)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_190),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_191),
.B(n_209),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_112),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_192),
.B(n_238),
.Y(n_266)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_135),
.Y(n_193)
);

INVx3_ASAP7_75t_SL g246 ( 
.A(n_193),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_194),
.A2(n_217),
.B1(n_226),
.B2(n_146),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_195),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_89),
.B1(n_88),
.B2(n_78),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_150),
.A2(n_62),
.B1(n_109),
.B2(n_44),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_197),
.A2(n_216),
.B1(n_222),
.B2(n_228),
.Y(n_284)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_198),
.Y(n_292)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_200),
.Y(n_287)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_201),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_202),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_150),
.A2(n_42),
.B1(n_50),
.B2(n_35),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_204),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_144),
.B(n_19),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_205),
.B(n_224),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_208),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_117),
.B(n_53),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_114),
.A2(n_50),
.B1(n_35),
.B2(n_31),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

INVx3_ASAP7_75t_SL g265 ( 
.A(n_214),
.Y(n_265)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_133),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_149),
.A2(n_20),
.B1(n_26),
.B2(n_17),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_140),
.Y(n_218)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_156),
.Y(n_219)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_140),
.Y(n_220)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_221),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_119),
.A2(n_50),
.B1(n_20),
.B2(n_26),
.Y(n_222)
);

NAND2xp33_ASAP7_75t_SL g223 ( 
.A(n_168),
.B(n_65),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_132),
.B(n_136),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_131),
.B(n_19),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_225),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_L g226 ( 
.A1(n_110),
.A2(n_26),
.B1(n_17),
.B2(n_24),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_161),
.A2(n_17),
.B1(n_24),
.B2(n_11),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_141),
.A2(n_24),
.B1(n_11),
.B2(n_12),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_145),
.B(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_229),
.B(n_245),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_127),
.B(n_16),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_230),
.B(n_138),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_179),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_231),
.A2(n_240),
.B1(n_243),
.B2(n_138),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_148),
.Y(n_232)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_116),
.Y(n_234)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_234),
.Y(n_295)
);

OA22x2_ASAP7_75t_SL g235 ( 
.A1(n_179),
.A2(n_132),
.B1(n_162),
.B2(n_135),
.Y(n_235)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_235),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_148),
.Y(n_236)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_236),
.Y(n_300)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_151),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_179),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_110),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_241),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_163),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_130),
.Y(n_241)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_163),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_244),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_128),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_171),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_118),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_136),
.C(n_125),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_247),
.B(n_275),
.C(n_223),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_211),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_250),
.B(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_253),
.Y(n_351)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_183),
.A2(n_132),
.B(n_15),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_254),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_188),
.B(n_174),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_256),
.B(n_302),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_185),
.B(n_166),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_262),
.B(n_286),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_268),
.A2(n_269),
.B1(n_280),
.B2(n_282),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_L g269 ( 
.A1(n_194),
.A2(n_174),
.B1(n_153),
.B2(n_118),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_211),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_212),
.B(n_155),
.Y(n_275)
);

OAI32xp33_ASAP7_75t_L g276 ( 
.A1(n_187),
.A2(n_153),
.A3(n_128),
.B1(n_146),
.B2(n_155),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_276),
.B(n_288),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_202),
.A2(n_126),
.B1(n_164),
.B2(n_143),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_196),
.A2(n_126),
.B1(n_164),
.B2(n_143),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_204),
.B(n_137),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_203),
.B(n_213),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_289),
.B(n_4),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_296),
.A2(n_193),
.B1(n_235),
.B2(n_137),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_211),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_303),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_181),
.B(n_1),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_211),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_231),
.B(n_243),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_304),
.B(n_303),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_305),
.A2(n_307),
.B1(n_308),
.B2(n_319),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_284),
.A2(n_235),
.B1(n_242),
.B2(n_220),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_284),
.A2(n_201),
.B1(n_198),
.B2(n_233),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_226),
.B1(n_208),
.B2(n_219),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_310),
.A2(n_329),
.B1(n_334),
.B2(n_350),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_312),
.B(n_339),
.Y(n_385)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_313),
.Y(n_358)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_259),
.Y(n_314)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_314),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_258),
.A2(n_180),
.B(n_189),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_315),
.A2(n_317),
.B(n_321),
.Y(n_375)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_259),
.Y(n_316)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_316),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_258),
.A2(n_186),
.B(n_225),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_290),
.A2(n_236),
.B1(n_232),
.B2(n_218),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_184),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_320),
.B(n_333),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_298),
.A2(n_182),
.B(n_221),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_SL g322 ( 
.A1(n_298),
.A2(n_137),
.B(n_210),
.C(n_195),
.Y(n_322)
);

AO22x1_ASAP7_75t_SL g355 ( 
.A1(n_322),
.A2(n_274),
.B1(n_301),
.B2(n_263),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_256),
.C(n_247),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_325),
.C(n_312),
.Y(n_359)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_259),
.Y(n_324)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_324),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_267),
.B(n_249),
.C(n_289),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_266),
.A2(n_239),
.B(n_13),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_326),
.A2(n_328),
.B(n_338),
.Y(n_383)
);

OAI22x1_ASAP7_75t_SL g327 ( 
.A1(n_290),
.A2(n_214),
.B1(n_207),
.B2(n_8),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_327),
.A2(n_346),
.B1(n_347),
.B2(n_349),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_296),
.A2(n_15),
.B(n_8),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_269),
.A2(n_8),
.B1(n_13),
.B2(n_4),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_292),
.Y(n_330)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_271),
.B(n_13),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_302),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_277),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_345),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_272),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_337),
.B(n_257),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_262),
.A2(n_4),
.B(n_6),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_287),
.Y(n_340)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_340),
.Y(n_396)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_287),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_341),
.Y(n_360)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_264),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_276),
.A2(n_4),
.B(n_6),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_343),
.A2(n_263),
.B(n_301),
.Y(n_378)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_287),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_344),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_248),
.A2(n_264),
.B1(n_246),
.B2(n_299),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_248),
.A2(n_246),
.B1(n_273),
.B2(n_252),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_295),
.B(n_293),
.C(n_291),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_348),
.B(n_313),
.C(n_340),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_246),
.A2(n_285),
.B1(n_252),
.B2(n_300),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_295),
.A2(n_279),
.B1(n_255),
.B2(n_291),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_293),
.B(n_255),
.Y(n_352)
);

NAND3xp33_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_354),
.C(n_292),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_278),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_353),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_279),
.B(n_274),
.Y(n_354)
);

OA22x2_ASAP7_75t_L g403 ( 
.A1(n_355),
.A2(n_309),
.B1(n_310),
.B2(n_322),
.Y(n_403)
);

AOI32xp33_ASAP7_75t_L g356 ( 
.A1(n_331),
.A2(n_300),
.A3(n_285),
.B1(n_260),
.B2(n_283),
.Y(n_356)
);

AOI21xp33_ASAP7_75t_L g397 ( 
.A1(n_356),
.A2(n_388),
.B(n_365),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_359),
.B(n_392),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_257),
.C(n_297),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_386),
.C(n_392),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_297),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_363),
.B(n_378),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_364),
.B(n_372),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_351),
.A2(n_283),
.B(n_260),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_365),
.A2(n_338),
.B(n_326),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_368),
.B(n_389),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_350),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_335),
.A2(n_265),
.B1(n_251),
.B2(n_261),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_373),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_307),
.A2(n_265),
.B1(n_278),
.B2(n_281),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_379),
.A2(n_341),
.B1(n_344),
.B2(n_329),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_306),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_314),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_281),
.Y(n_381)
);

XNOR2x1_ASAP7_75t_L g431 ( 
.A(n_381),
.B(n_395),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_308),
.A2(n_261),
.B1(n_251),
.B2(n_265),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_384),
.A2(n_349),
.B1(n_316),
.B2(n_324),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_339),
.B(n_331),
.C(n_348),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_318),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_393),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_336),
.B(n_337),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_311),
.A2(n_343),
.B1(n_309),
.B2(n_321),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_390),
.A2(n_327),
.B1(n_319),
.B2(n_347),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_315),
.A2(n_351),
.B(n_317),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_391),
.A2(n_375),
.B(n_393),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_332),
.B(n_333),
.Y(n_392)
);

A2O1A1Ixp33_ASAP7_75t_L g393 ( 
.A1(n_335),
.A2(n_328),
.B(n_322),
.C(n_305),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_346),
.Y(n_394)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_394),
.Y(n_401)
);

BUFx12f_ASAP7_75t_SL g453 ( 
.A(n_397),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_359),
.B(n_385),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_404),
.C(n_422),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_402),
.A2(n_377),
.B1(n_373),
.B2(n_376),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_403),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_362),
.B(n_381),
.C(n_385),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_405),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_406),
.A2(n_417),
.B(n_419),
.Y(n_433)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_361),
.Y(n_407)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_407),
.Y(n_450)
);

NOR2x1p5_ASAP7_75t_SL g408 ( 
.A(n_370),
.B(n_322),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_430),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_410),
.B(n_360),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_411),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_412),
.A2(n_416),
.B1(n_424),
.B2(n_401),
.Y(n_458)
);

INVx13_ASAP7_75t_L g413 ( 
.A(n_374),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_413),
.Y(n_439)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_361),
.Y(n_414)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_414),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_390),
.A2(n_322),
.B1(n_342),
.B2(n_353),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_415),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_370),
.A2(n_334),
.B1(n_353),
.B2(n_330),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_375),
.A2(n_391),
.B(n_383),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_378),
.A2(n_394),
.B(n_383),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_421),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_386),
.C(n_357),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_357),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_429),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_372),
.A2(n_377),
.B1(n_379),
.B2(n_363),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_369),
.Y(n_425)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_425),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_427),
.C(n_371),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_367),
.B(n_380),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_369),
.Y(n_428)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_428),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_382),
.Y(n_429)
);

INVx8_ASAP7_75t_L g430 ( 
.A(n_366),
.Y(n_430)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_436),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_360),
.Y(n_440)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_440),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_409),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_400),
.B(n_371),
.C(n_396),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_442),
.B(n_444),
.C(n_452),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_396),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_443),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_382),
.C(n_358),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_358),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_432),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_355),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_448),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_418),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_462),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_355),
.C(n_387),
.Y(n_452)
);

INVxp33_ASAP7_75t_SL g482 ( 
.A(n_454),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_402),
.A2(n_374),
.B1(n_387),
.B2(n_401),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_457),
.A2(n_458),
.B1(n_421),
.B2(n_399),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_398),
.B(n_426),
.C(n_422),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_463),
.C(n_399),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_407),
.B(n_428),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_398),
.B(n_427),
.C(n_432),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_464),
.B(n_468),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_465),
.B(n_469),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_441),
.B(n_417),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_434),
.B(n_420),
.Y(n_469)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_439),
.Y(n_471)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_471),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_451),
.B(n_420),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_473),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_433),
.A2(n_449),
.B(n_419),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_463),
.B(n_425),
.Y(n_475)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_475),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_476),
.A2(n_446),
.B1(n_445),
.B2(n_403),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_479),
.C(n_483),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_434),
.B(n_460),
.C(n_444),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_442),
.B(n_406),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_486),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_447),
.B(n_414),
.C(n_403),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_436),
.B(n_430),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_487),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_433),
.A2(n_408),
.B(n_416),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_473),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_440),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_453),
.B(n_408),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_458),
.B(n_412),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_488),
.B(n_489),
.C(n_457),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_403),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_488),
.Y(n_492)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_492),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_494),
.B(n_455),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_482),
.A2(n_446),
.B1(n_435),
.B2(n_448),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_495),
.A2(n_501),
.B1(n_505),
.B2(n_476),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_437),
.C(n_454),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_507),
.C(n_510),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_467),
.A2(n_446),
.B1(n_435),
.B2(n_437),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_481),
.B(n_453),
.Y(n_502)
);

NAND3xp33_ASAP7_75t_L g514 ( 
.A(n_502),
.B(n_465),
.C(n_477),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_503),
.A2(n_494),
.B1(n_496),
.B2(n_497),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_485),
.A2(n_456),
.B1(n_453),
.B2(n_443),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_470),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_506),
.A2(n_509),
.B1(n_438),
.B2(n_405),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_474),
.B(n_439),
.C(n_462),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_508),
.A2(n_466),
.B(n_483),
.Y(n_512)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_478),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_474),
.B(n_439),
.C(n_461),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_512),
.A2(n_518),
.B(n_490),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_503),
.A2(n_478),
.B1(n_489),
.B2(n_487),
.Y(n_513)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_513),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_514),
.B(n_515),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_510),
.B(n_469),
.C(n_486),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_468),
.C(n_480),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_516),
.B(n_517),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_508),
.A2(n_464),
.B(n_471),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_491),
.B(n_450),
.C(n_455),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_519),
.B(n_520),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_505),
.B(n_450),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_523),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_499),
.B(n_493),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_522),
.B(n_498),
.Y(n_535)
);

OA21x2_ASAP7_75t_L g523 ( 
.A1(n_501),
.A2(n_459),
.B(n_461),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_504),
.B(n_459),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_524),
.B(n_525),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_495),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_529),
.A2(n_541),
.B(n_512),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_530),
.B(n_535),
.Y(n_546)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_519),
.B(n_491),
.Y(n_531)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_531),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_511),
.B(n_498),
.C(n_504),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_538),
.B(n_539),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_511),
.B(n_500),
.C(n_438),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_515),
.B(n_500),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_540),
.B(n_516),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_518),
.A2(n_413),
.B(n_524),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_532),
.B(n_533),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_542),
.B(n_544),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_545),
.B(n_549),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_538),
.B(n_527),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_547),
.B(n_548),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_539),
.B(n_530),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_536),
.A2(n_523),
.B1(n_526),
.B2(n_513),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_527),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_550),
.B(n_528),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_551),
.A2(n_529),
.B(n_520),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_555),
.A2(n_557),
.B(n_549),
.Y(n_561)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_556),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_543),
.A2(n_517),
.B(n_523),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_554),
.A2(n_553),
.B(n_545),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_558),
.A2(n_560),
.B(n_561),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_552),
.B(n_546),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_559),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_562),
.B(n_528),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_564),
.A2(n_563),
.B(n_521),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_565),
.A2(n_523),
.B(n_537),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_566),
.B(n_537),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_567),
.B(n_413),
.Y(n_568)
);


endmodule