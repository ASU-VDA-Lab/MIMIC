module fake_jpeg_23513_n_300 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_33),
.B(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_13),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_20),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_42),
.A2(n_50),
.B(n_22),
.C(n_27),
.Y(n_81)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_46),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_16),
.B1(n_18),
.B2(n_14),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_16),
.B1(n_14),
.B2(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_23),
.B(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_15),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_60),
.B(n_58),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_26),
.B(n_25),
.C(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_72),
.B1(n_19),
.B2(n_38),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_26),
.B1(n_28),
.B2(n_37),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_35),
.B1(n_34),
.B2(n_16),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_13),
.Y(n_103)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_71),
.Y(n_84)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_26),
.B1(n_28),
.B2(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_73),
.Y(n_98)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_36),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_58),
.C(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_56),
.B(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_21),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_68),
.B(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_83),
.B(n_91),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_92),
.B(n_94),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_42),
.B(n_39),
.C(n_37),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_42),
.B(n_24),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_97),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_96),
.A2(n_104),
.B1(n_70),
.B2(n_35),
.Y(n_119)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_100),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_71),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_66),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_33),
.B1(n_19),
.B2(n_21),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_46),
.C(n_53),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_107),
.C(n_66),
.Y(n_130)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_125),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_63),
.Y(n_107)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_63),
.A3(n_75),
.B1(n_61),
.B2(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_103),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_94),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_116),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_78),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_61),
.B1(n_63),
.B2(n_34),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_75),
.B1(n_76),
.B2(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_120),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_128),
.B1(n_85),
.B2(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_60),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_122),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_83),
.A2(n_35),
.B1(n_44),
.B2(n_51),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_44),
.B1(n_65),
.B2(n_87),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_79),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_124),
.B(n_126),
.Y(n_141)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_145),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_134),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_103),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_106),
.B1(n_114),
.B2(n_113),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_127),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_143),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_0),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_148),
.B(n_114),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_118),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_111),
.B1(n_107),
.B2(n_123),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_147),
.B1(n_152),
.B2(n_153),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_65),
.B1(n_101),
.B2(n_87),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_116),
.B1(n_107),
.B2(n_120),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_109),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_150),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_37),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_107),
.A2(n_41),
.B1(n_57),
.B2(n_47),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_107),
.A2(n_97),
.B1(n_99),
.B2(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_156),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_122),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_162),
.Y(n_184)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_124),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_171),
.B(n_177),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_152),
.B1(n_133),
.B2(n_115),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_131),
.B(n_123),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_116),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_172),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_178),
.B1(n_117),
.B2(n_119),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_125),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_115),
.B(n_117),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_37),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_196),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_129),
.B1(n_149),
.B2(n_133),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_183),
.A2(n_197),
.B1(n_172),
.B2(n_161),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_187),
.B1(n_202),
.B2(n_159),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_168),
.A2(n_133),
.B1(n_119),
.B2(n_115),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_110),
.B(n_142),
.C(n_112),
.Y(n_191)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_142),
.C(n_134),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_182),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_110),
.C(n_52),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_198),
.C(n_201),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_176),
.B(n_39),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_128),
.B1(n_106),
.B2(n_90),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_39),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_169),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_158),
.A2(n_128),
.B1(n_73),
.B2(n_67),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_189),
.B1(n_188),
.B2(n_198),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_195),
.A2(n_160),
.B1(n_173),
.B2(n_156),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_SL g229 ( 
.A1(n_206),
.A2(n_211),
.B(n_213),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_214),
.B1(n_222),
.B2(n_187),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_162),
.B1(n_179),
.B2(n_154),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_166),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_218),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_164),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_193),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_219),
.A2(n_181),
.B(n_199),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_170),
.C(n_167),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_221),
.C(n_223),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_170),
.C(n_155),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_17),
.B1(n_15),
.B2(n_29),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_52),
.C(n_55),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_228),
.B1(n_230),
.B2(n_55),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_188),
.C(n_203),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_241),
.C(n_238),
.Y(n_249)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_194),
.B1(n_201),
.B2(n_202),
.Y(n_230)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_235),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_219),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_183),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_238),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_214),
.B(n_203),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_216),
.B(n_181),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_205),
.C(n_223),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_199),
.C(n_52),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_205),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_245),
.Y(n_261)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_239),
.A2(n_215),
.B(n_212),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_211),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_251),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_229),
.A2(n_102),
.B1(n_73),
.B2(n_67),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_248),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_252),
.C(n_254),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_102),
.C(n_52),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_52),
.C(n_49),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_255),
.A2(n_256),
.B1(n_3),
.B2(n_4),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_SL g256 ( 
.A1(n_228),
.A2(n_224),
.B(n_230),
.C(n_237),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_247),
.A2(n_234),
.B1(n_236),
.B2(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_231),
.C(n_39),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_263),
.C(n_265),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_263),
.B1(n_269),
.B2(n_265),
.Y(n_274)
);

XOR2x2_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_12),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_262),
.A2(n_256),
.B(n_4),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_0),
.C(n_2),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_0),
.C(n_3),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_12),
.B1(n_22),
.B2(n_5),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_266),
.B(n_7),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_12),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_269),
.B1(n_3),
.B2(n_6),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_253),
.B(n_256),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_259),
.B(n_268),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_254),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_271),
.B(n_272),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_276),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_3),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_277),
.B(n_280),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_6),
.C(n_7),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.C(n_7),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_6),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_273),
.B(n_275),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_7),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_8),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_8),
.C(n_9),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_286),
.A2(n_273),
.B(n_278),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_290),
.C(n_291),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_287),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_289),
.A2(n_292),
.B(n_283),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_283),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_293),
.C(n_10),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_296),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_9),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_298),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_9),
.B1(n_10),
.B2(n_295),
.Y(n_300)
);


endmodule