module real_jpeg_5080_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_1),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_1),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_1),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_1),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_2),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_2),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_2),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_2),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_2),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_2),
.B(n_234),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_3),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_4),
.B(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_5),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_5),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_5),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_5),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_5),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_5),
.B(n_250),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_5),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_5),
.B(n_230),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_6),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_6),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_6),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_6),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_6),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_6),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_6),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_7),
.B(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_7),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_7),
.B(n_81),
.Y(n_156)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_9),
.Y(n_139)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_9),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_9),
.Y(n_268)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_10),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_10),
.B(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_11),
.Y(n_171)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_13),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_14),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_14),
.B(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_14),
.B(n_71),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_14),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_14),
.B(n_81),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_14),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_15),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_15),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_15),
.B(n_83),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_15),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_15),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_15),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_15),
.B(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_16),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_17),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_17),
.B(n_167),
.Y(n_166)
);

XNOR2x2_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_195),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_194),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_146),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_22),
.B(n_146),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_100),
.C(n_132),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_23),
.B(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_62),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_24),
.B(n_63),
.C(n_78),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_42),
.C(n_51),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_25),
.B(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_26),
.B(n_36),
.C(n_40),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_29),
.Y(n_175)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_29),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_39),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_39),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_42),
.B(n_51),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_43),
.B(n_47),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_50),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.C(n_58),
.Y(n_51)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_52),
.B(n_54),
.CI(n_58),
.CON(n_205),
.SN(n_205)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_57),
.Y(n_231)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_57),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_60),
.Y(n_168)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_61),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_78),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_64),
.B(n_70),
.C(n_74),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_68),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_68),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_87),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_80),
.B(n_82),
.C(n_87),
.Y(n_153)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.C(n_97),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_97),
.Y(n_131)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_100),
.B(n_132),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_122),
.C(n_129),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_101),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_115),
.C(n_119),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_102),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_109),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_103),
.A2(n_104),
.B1(n_109),
.B2(n_110),
.Y(n_226)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_108),
.Y(n_266)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_114),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_115),
.B(n_119),
.Y(n_240)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_122),
.A2(n_129),
.B1(n_130),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B(n_128),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_124),
.Y(n_128)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_128),
.B(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_133),
.C(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_143),
.B2(n_145),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_138),
.C(n_140),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_164),
.B1(n_192),
.B2(n_193),
.Y(n_148)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_163),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_162),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_176),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_165),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.CI(n_172),
.CON(n_165),
.SN(n_165)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_188),
.B2(n_189),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_184),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI21x1_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_319),
.B(n_323),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_241),
.B(n_318),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_221),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_198),
.B(n_221),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_220),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_199),
.B(n_204),
.C(n_218),
.Y(n_322)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_218),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.C(n_217),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_223),
.Y(n_222)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_205),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_207),
.B1(n_217),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.C(n_215),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_208),
.A2(n_209),
.B1(n_215),
.B2(n_216),
.Y(n_311)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_210),
.B(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_217),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.C(n_239),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_222),
.B(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_225),
.B(n_239),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.C(n_232),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_226),
.B(n_227),
.Y(n_304)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_232),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_237),
.Y(n_283)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21x1_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_313),
.B(n_317),
.Y(n_241)
);

OA21x2_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_298),
.B(n_312),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_280),
.B(n_297),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_269),
.B(n_279),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_252),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_252),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_249),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_261),
.B2(n_262),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_256),
.C(n_261),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_267),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_274),
.B(n_278),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_272),
.Y(n_278)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_296),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_296),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_284),
.C(n_300),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_290),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_293),
.C(n_295),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

INVx11_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_291),
.Y(n_295)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_301),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_308),
.C(n_309),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_315),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_322),
.Y(n_323)
);


endmodule