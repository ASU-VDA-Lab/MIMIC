module fake_netlist_1_6240_n_935 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_935);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_935;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_383;
wire n_288;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_704;
wire n_611;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_245;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_898;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_912;
wire n_924;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_406;
wire n_395;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g231 ( .A(n_195), .Y(n_231) );
INVxp67_ASAP7_75t_SL g232 ( .A(n_156), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_214), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_112), .Y(n_234) );
INVxp67_ASAP7_75t_SL g235 ( .A(n_99), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_11), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_134), .Y(n_237) );
INVxp67_ASAP7_75t_SL g238 ( .A(n_167), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_76), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_43), .Y(n_240) );
NOR2xp67_ASAP7_75t_L g241 ( .A(n_115), .B(n_181), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_202), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_213), .Y(n_243) );
BUFx3_ASAP7_75t_L g244 ( .A(n_142), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_121), .Y(n_245) );
CKINVDCx16_ASAP7_75t_R g246 ( .A(n_66), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_135), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_185), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_179), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_219), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_43), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_192), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_108), .Y(n_253) );
INVxp67_ASAP7_75t_SL g254 ( .A(n_31), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_67), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_85), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_164), .Y(n_257) );
INVxp67_ASAP7_75t_SL g258 ( .A(n_133), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_70), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_147), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_83), .Y(n_261) );
CKINVDCx16_ASAP7_75t_R g262 ( .A(n_130), .Y(n_262) );
BUFx2_ASAP7_75t_SL g263 ( .A(n_17), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_143), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g265 ( .A(n_92), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_180), .Y(n_266) );
NOR2xp67_ASAP7_75t_L g267 ( .A(n_73), .B(n_136), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_145), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_90), .B(n_132), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_198), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_101), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_26), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_207), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_160), .Y(n_274) );
INVxp33_ASAP7_75t_SL g275 ( .A(n_140), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_120), .Y(n_276) );
INVxp67_ASAP7_75t_SL g277 ( .A(n_47), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_6), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_153), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_19), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_75), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_109), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_201), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_81), .Y(n_284) );
BUFx10_ASAP7_75t_L g285 ( .A(n_186), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_223), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_91), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_212), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g289 ( .A(n_124), .Y(n_289) );
CKINVDCx14_ASAP7_75t_R g290 ( .A(n_196), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_161), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_127), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_65), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_218), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_197), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_204), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_78), .Y(n_297) );
INVxp67_ASAP7_75t_SL g298 ( .A(n_148), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_98), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_191), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_23), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_13), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_193), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_159), .Y(n_304) );
INVxp67_ASAP7_75t_SL g305 ( .A(n_82), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_72), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_32), .Y(n_307) );
INVxp33_ASAP7_75t_L g308 ( .A(n_118), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_56), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_209), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_221), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_228), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_3), .Y(n_313) );
INVxp33_ASAP7_75t_L g314 ( .A(n_162), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_187), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_35), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_158), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_21), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_30), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_188), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_17), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_217), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_80), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_199), .Y(n_324) );
NOR2xp67_ASAP7_75t_L g325 ( .A(n_70), .B(n_144), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_206), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_44), .Y(n_327) );
BUFx10_ASAP7_75t_L g328 ( .A(n_22), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_0), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_2), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_205), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_79), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_116), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_203), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_71), .Y(n_335) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_229), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_165), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_166), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_29), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_169), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_149), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_15), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_138), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_163), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_208), .Y(n_345) );
INVxp33_ASAP7_75t_L g346 ( .A(n_102), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_42), .Y(n_347) );
INVxp67_ASAP7_75t_L g348 ( .A(n_260), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_237), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_237), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_264), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_260), .B(n_1), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_244), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_237), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_285), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_285), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_271), .B(n_1), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_264), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_237), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_313), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_246), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_237), .Y(n_362) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_306), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_306), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_255), .B(n_2), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_271), .B(n_3), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_285), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_308), .B(n_4), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_313), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_306), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_306), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_306), .Y(n_372) );
OA21x2_ASAP7_75t_L g373 ( .A1(n_261), .A2(n_77), .B(n_74), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_261), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_280), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_329), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_329), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_262), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_330), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_327), .Y(n_380) );
AND3x2_ASAP7_75t_L g381 ( .A(n_343), .B(n_7), .C(n_8), .Y(n_381) );
NAND2x1_ASAP7_75t_L g382 ( .A(n_255), .B(n_7), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_266), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_244), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_355), .B(n_308), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_357), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_357), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_348), .B(n_236), .Y(n_388) );
AND2x6_ASAP7_75t_L g389 ( .A(n_352), .B(n_300), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_353), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_348), .B(n_236), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_357), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_355), .B(n_314), .Y(n_393) );
INVx6_ASAP7_75t_L g394 ( .A(n_357), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_350), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_357), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_355), .B(n_346), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_350), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_366), .B(n_266), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_350), .Y(n_400) );
OR2x2_ASAP7_75t_SL g401 ( .A(n_380), .B(n_265), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_366), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_368), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_355), .B(n_356), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_352), .A2(n_275), .B1(n_319), .B2(n_280), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_356), .B(n_346), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_356), .B(n_319), .Y(n_407) );
OR2x6_ASAP7_75t_L g408 ( .A(n_352), .B(n_263), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_350), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_356), .B(n_268), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_378), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_378), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_356), .B(n_268), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_367), .B(n_283), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_366), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_367), .B(n_272), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_361), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_350), .Y(n_418) );
OAI22x1_ASAP7_75t_L g419 ( .A1(n_375), .A2(n_339), .B1(n_321), .B2(n_277), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_366), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_366), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_368), .Y(n_422) );
AO22x2_ASAP7_75t_L g423 ( .A1(n_352), .A2(n_263), .B1(n_293), .B2(n_254), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_353), .Y(n_424) );
BUFx3_ASAP7_75t_L g425 ( .A(n_384), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_351), .B(n_284), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_368), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_408), .B(n_381), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_423), .A2(n_405), .B1(n_408), .B2(n_403), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_403), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_416), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_422), .B(n_233), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_411), .B(n_365), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_394), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_390), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_385), .B(n_351), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_385), .B(n_358), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_407), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_406), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
BUFx4f_ASAP7_75t_L g441 ( .A(n_389), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_423), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_423), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_427), .B(n_358), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_394), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_394), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_402), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_393), .A2(n_289), .B1(n_312), .B2(n_234), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_393), .B(n_382), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_388), .B(n_233), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_397), .B(n_382), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_388), .B(n_381), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_391), .B(n_243), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_412), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_399), .A2(n_387), .B(n_386), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_402), .Y(n_456) );
INVx4_ASAP7_75t_L g457 ( .A(n_389), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_424), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_421), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_421), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_392), .B(n_275), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_419), .B(n_328), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_396), .B(n_249), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_425), .Y(n_464) );
INVx5_ASAP7_75t_L g465 ( .A(n_389), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_415), .B(n_270), .Y(n_466) );
INVx4_ASAP7_75t_L g467 ( .A(n_389), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_420), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_404), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_399), .B(n_270), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_410), .B(n_281), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_410), .A2(n_332), .B1(n_340), .B2(n_312), .Y(n_472) );
INVxp67_ASAP7_75t_L g473 ( .A(n_426), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_413), .B(n_332), .Y(n_474) );
INVx6_ASAP7_75t_L g475 ( .A(n_425), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_413), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_414), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_417), .Y(n_478) );
NAND2x1p5_ASAP7_75t_L g479 ( .A(n_426), .B(n_293), .Y(n_479) );
BUFx3_ASAP7_75t_L g480 ( .A(n_401), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_395), .B(n_281), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_395), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_398), .B(n_344), .Y(n_483) );
OAI22xp5_ASAP7_75t_SL g484 ( .A1(n_398), .A2(n_302), .B1(n_251), .B2(n_259), .Y(n_484) );
INVx2_ASAP7_75t_SL g485 ( .A(n_398), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_400), .B(n_328), .Y(n_486) );
INVx4_ASAP7_75t_L g487 ( .A(n_400), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_409), .B(n_304), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_409), .A2(n_316), .B1(n_272), .B2(n_290), .Y(n_489) );
OR2x6_ASAP7_75t_L g490 ( .A(n_418), .B(n_240), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_418), .B(n_360), .Y(n_491) );
OR2x2_ASAP7_75t_SL g492 ( .A(n_418), .B(n_373), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_390), .Y(n_493) );
BUFx3_ASAP7_75t_L g494 ( .A(n_416), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_422), .B(n_323), .Y(n_495) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_394), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_422), .B(n_323), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_403), .Y(n_498) );
INVx6_ASAP7_75t_L g499 ( .A(n_416), .Y(n_499) );
BUFx12f_ASAP7_75t_L g500 ( .A(n_417), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_403), .B(n_331), .Y(n_501) );
BUFx4f_ASAP7_75t_L g502 ( .A(n_408), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_423), .Y(n_503) );
BUFx3_ASAP7_75t_L g504 ( .A(n_500), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_503), .A2(n_443), .B1(n_442), .B2(n_429), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_473), .A2(n_383), .B1(n_374), .B2(n_278), .Y(n_506) );
NOR2xp67_ASAP7_75t_L g507 ( .A(n_465), .B(n_269), .Y(n_507) );
O2A1O1Ixp5_ASAP7_75t_L g508 ( .A1(n_449), .A2(n_235), .B(n_238), .C(n_232), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_436), .A2(n_373), .B(n_298), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_439), .B(n_374), .Y(n_510) );
NOR2xp33_ASAP7_75t_SL g511 ( .A(n_457), .B(n_335), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_502), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_436), .A2(n_373), .B(n_305), .Y(n_513) );
INVx3_ASAP7_75t_L g514 ( .A(n_446), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_437), .A2(n_373), .B(n_336), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_428), .B(n_301), .Y(n_516) );
BUFx4f_ASAP7_75t_L g517 ( .A(n_428), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_473), .A2(n_383), .B1(n_374), .B2(n_309), .Y(n_518) );
BUFx2_ASAP7_75t_L g519 ( .A(n_483), .Y(n_519) );
BUFx2_ASAP7_75t_L g520 ( .A(n_483), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_437), .A2(n_373), .B(n_258), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_449), .A2(n_239), .B(n_231), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_438), .B(n_318), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_451), .A2(n_245), .B(n_242), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_430), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_498), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_474), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_496), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_496), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_469), .B(n_383), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_445), .Y(n_531) );
BUFx12f_ASAP7_75t_L g532 ( .A(n_478), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_451), .A2(n_248), .B(n_247), .Y(n_533) );
NOR2xp67_ASAP7_75t_L g534 ( .A(n_465), .B(n_84), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_440), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_499), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_501), .B(n_335), .Y(n_537) );
INVx5_ASAP7_75t_L g538 ( .A(n_490), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_457), .Y(n_539) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_467), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_476), .B(n_342), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_477), .B(n_347), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_452), .Y(n_543) );
BUFx4f_ASAP7_75t_L g544 ( .A(n_499), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_455), .A2(n_252), .B(n_250), .Y(n_545) );
BUFx2_ASAP7_75t_L g546 ( .A(n_472), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_447), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_455), .A2(n_325), .B(n_376), .C(n_369), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_444), .A2(n_377), .B(n_379), .C(n_376), .Y(n_549) );
INVx6_ASAP7_75t_L g550 ( .A(n_494), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_491), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_467), .B(n_253), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_461), .A2(n_257), .B(n_256), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_456), .Y(n_554) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_490), .Y(n_555) );
INVx8_ASAP7_75t_L g556 ( .A(n_465), .Y(n_556) );
INVx2_ASAP7_75t_SL g557 ( .A(n_479), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_459), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_468), .A2(n_274), .B(n_276), .C(n_273), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_460), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_435), .Y(n_561) );
OAI22xp5_ASAP7_75t_SL g562 ( .A1(n_480), .A2(n_282), .B1(n_286), .B2(n_279), .Y(n_562) );
BUFx2_ASAP7_75t_L g563 ( .A(n_448), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_463), .A2(n_288), .B(n_287), .Y(n_564) );
BUFx12f_ASAP7_75t_L g565 ( .A(n_462), .Y(n_565) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_490), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_450), .B(n_291), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_479), .B(n_292), .Y(n_568) );
NOR2xp67_ASAP7_75t_L g569 ( .A(n_466), .B(n_86), .Y(n_569) );
BUFx2_ASAP7_75t_L g570 ( .A(n_484), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_495), .B(n_307), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_466), .Y(n_572) );
INVx2_ASAP7_75t_SL g573 ( .A(n_453), .Y(n_573) );
INVx4_ASAP7_75t_L g574 ( .A(n_441), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_486), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_475), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_458), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_497), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_432), .B(n_294), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_471), .B(n_295), .Y(n_580) );
O2A1O1Ixp33_ASAP7_75t_L g581 ( .A1(n_471), .A2(n_296), .B(n_299), .C(n_297), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_470), .B(n_303), .Y(n_582) );
INVx3_ASAP7_75t_L g583 ( .A(n_475), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_493), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_481), .Y(n_585) );
OR2x6_ASAP7_75t_L g586 ( .A(n_481), .B(n_241), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_488), .Y(n_587) );
INVx3_ASAP7_75t_L g588 ( .A(n_487), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_492), .A2(n_311), .B1(n_315), .B2(n_310), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_489), .B(n_322), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_464), .B(n_9), .Y(n_591) );
OR2x6_ASAP7_75t_L g592 ( .A(n_485), .B(n_267), .Y(n_592) );
AO32x1_ASAP7_75t_L g593 ( .A1(n_482), .A2(n_349), .A3(n_364), .B1(n_371), .B2(n_370), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_434), .Y(n_594) );
BUFx2_ASAP7_75t_L g595 ( .A(n_454), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_439), .B(n_326), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_503), .A2(n_334), .B1(n_337), .B2(n_333), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_439), .B(n_338), .Y(n_598) );
INVx4_ASAP7_75t_L g599 ( .A(n_502), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_434), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_433), .B(n_341), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_439), .B(n_345), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_431), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_439), .B(n_284), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_439), .B(n_317), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_436), .A2(n_320), .B(n_317), .Y(n_606) );
AO21x2_ASAP7_75t_L g607 ( .A1(n_548), .A2(n_324), .B(n_320), .Y(n_607) );
OAI21x1_ASAP7_75t_L g608 ( .A1(n_509), .A2(n_364), .B(n_349), .Y(n_608) );
AO31x2_ASAP7_75t_L g609 ( .A1(n_589), .A2(n_370), .A3(n_371), .B(n_364), .Y(n_609) );
OAI21x1_ASAP7_75t_L g610 ( .A1(n_513), .A2(n_371), .B(n_370), .Y(n_610) );
OAI21x1_ASAP7_75t_L g611 ( .A1(n_515), .A2(n_521), .B(n_534), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_525), .Y(n_612) );
OAI21xp5_ASAP7_75t_L g613 ( .A1(n_572), .A2(n_384), .B(n_354), .Y(n_613) );
OAI21x1_ASAP7_75t_L g614 ( .A1(n_530), .A2(n_384), .B(n_354), .Y(n_614) );
OAI21x1_ASAP7_75t_SL g615 ( .A1(n_557), .A2(n_10), .B(n_11), .Y(n_615) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_589), .A2(n_581), .B(n_586), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_585), .A2(n_508), .B(n_545), .Y(n_617) );
AO21x2_ASAP7_75t_L g618 ( .A1(n_569), .A2(n_384), .B(n_354), .Y(n_618) );
OAI21x1_ASAP7_75t_L g619 ( .A1(n_530), .A2(n_354), .B(n_350), .Y(n_619) );
INVx3_ASAP7_75t_SL g620 ( .A(n_599), .Y(n_620) );
BUFx2_ASAP7_75t_L g621 ( .A(n_595), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_526), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_578), .B(n_10), .Y(n_623) );
INVx2_ASAP7_75t_SL g624 ( .A(n_517), .Y(n_624) );
OA21x2_ASAP7_75t_L g625 ( .A1(n_606), .A2(n_354), .B(n_350), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_563), .A2(n_372), .B1(n_363), .B2(n_362), .Y(n_626) );
INVxp67_ASAP7_75t_L g627 ( .A(n_555), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_538), .B(n_372), .Y(n_628) );
NOR2xp67_ASAP7_75t_L g629 ( .A(n_532), .B(n_12), .Y(n_629) );
CKINVDCx6p67_ASAP7_75t_R g630 ( .A(n_504), .Y(n_630) );
BUFx3_ASAP7_75t_L g631 ( .A(n_550), .Y(n_631) );
OAI21x1_ASAP7_75t_L g632 ( .A1(n_510), .A2(n_362), .B(n_359), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_564), .A2(n_362), .B(n_359), .Y(n_633) );
OAI21x1_ASAP7_75t_L g634 ( .A1(n_510), .A2(n_362), .B(n_359), .Y(n_634) );
NAND2x1p5_ASAP7_75t_L g635 ( .A(n_538), .B(n_363), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_551), .Y(n_636) );
OAI21x1_ASAP7_75t_L g637 ( .A1(n_506), .A2(n_372), .B(n_363), .Y(n_637) );
OAI21x1_ASAP7_75t_L g638 ( .A1(n_518), .A2(n_507), .B(n_604), .Y(n_638) );
NAND2x1_ASAP7_75t_L g639 ( .A(n_555), .B(n_363), .Y(n_639) );
OAI21x1_ASAP7_75t_L g640 ( .A1(n_518), .A2(n_372), .B(n_363), .Y(n_640) );
BUFx8_ASAP7_75t_SL g641 ( .A(n_565), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_603), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_505), .A2(n_372), .B1(n_15), .B2(n_16), .Y(n_643) );
OAI21x1_ASAP7_75t_L g644 ( .A1(n_507), .A2(n_88), .B(n_87), .Y(n_644) );
OAI21x1_ASAP7_75t_L g645 ( .A1(n_604), .A2(n_93), .B(n_89), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_523), .B(n_14), .Y(n_646) );
OA21x2_ASAP7_75t_L g647 ( .A1(n_522), .A2(n_95), .B(n_94), .Y(n_647) );
OAI21x1_ASAP7_75t_L g648 ( .A1(n_605), .A2(n_97), .B(n_96), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_547), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_597), .A2(n_16), .B1(n_18), .B2(n_20), .Y(n_650) );
OAI21x1_ASAP7_75t_L g651 ( .A1(n_524), .A2(n_103), .B(n_100), .Y(n_651) );
OAI21x1_ASAP7_75t_L g652 ( .A1(n_533), .A2(n_105), .B(n_104), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_527), .B(n_18), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_596), .B(n_20), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_596), .B(n_24), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_554), .Y(n_656) );
OR2x6_ASAP7_75t_L g657 ( .A(n_566), .B(n_25), .Y(n_657) );
OAI21x1_ASAP7_75t_L g658 ( .A1(n_588), .A2(n_107), .B(n_106), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_512), .B(n_543), .Y(n_659) );
OAI21x1_ASAP7_75t_L g660 ( .A1(n_588), .A2(n_111), .B(n_110), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_566), .B(n_113), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_593), .A2(n_117), .B(n_114), .Y(n_662) );
OAI21x1_ASAP7_75t_L g663 ( .A1(n_514), .A2(n_122), .B(n_119), .Y(n_663) );
AO21x2_ASAP7_75t_L g664 ( .A1(n_549), .A2(n_125), .B(n_123), .Y(n_664) );
BUFx10_ASAP7_75t_L g665 ( .A(n_516), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_575), .B(n_27), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_560), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_598), .B(n_27), .Y(n_668) );
INVx1_ASAP7_75t_SL g669 ( .A(n_535), .Y(n_669) );
OAI21x1_ASAP7_75t_SL g670 ( .A1(n_568), .A2(n_28), .B(n_29), .Y(n_670) );
OAI21x1_ASAP7_75t_L g671 ( .A1(n_514), .A2(n_128), .B(n_126), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_601), .B(n_28), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_598), .B(n_33), .Y(n_673) );
BUFx12f_ASAP7_75t_L g674 ( .A(n_516), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_573), .B(n_34), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_553), .B(n_36), .Y(n_676) );
AO32x2_ASAP7_75t_L g677 ( .A1(n_562), .A2(n_36), .A3(n_37), .B1(n_38), .B2(n_39), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_558), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_597), .A2(n_39), .B1(n_40), .B2(n_41), .Y(n_679) );
INVxp67_ASAP7_75t_L g680 ( .A(n_519), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_520), .A2(n_511), .B1(n_567), .B2(n_537), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_561), .Y(n_682) );
OAI21x1_ASAP7_75t_L g683 ( .A1(n_528), .A2(n_150), .B(n_227), .Y(n_683) );
OAI21x1_ASAP7_75t_L g684 ( .A1(n_594), .A2(n_151), .B(n_226), .Y(n_684) );
AND2x4_ASAP7_75t_L g685 ( .A(n_574), .B(n_41), .Y(n_685) );
O2A1O1Ixp33_ASAP7_75t_SL g686 ( .A1(n_587), .A2(n_146), .B(n_225), .C(n_224), .Y(n_686) );
INVxp67_ASAP7_75t_SL g687 ( .A(n_568), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_541), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_541), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_SL g690 ( .A1(n_587), .A2(n_152), .B(n_222), .C(n_220), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_544), .B(n_45), .Y(n_691) );
AND2x4_ASAP7_75t_L g692 ( .A(n_574), .B(n_46), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_577), .Y(n_693) );
AO31x2_ASAP7_75t_L g694 ( .A1(n_559), .A2(n_46), .A3(n_47), .B(n_48), .Y(n_694) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_539), .Y(n_695) );
AO31x2_ASAP7_75t_L g696 ( .A1(n_582), .A2(n_49), .A3(n_50), .B(n_51), .Y(n_696) );
OR2x6_ASAP7_75t_L g697 ( .A(n_556), .B(n_52), .Y(n_697) );
AO21x2_ASAP7_75t_L g698 ( .A1(n_582), .A2(n_155), .B(n_216), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_602), .A2(n_52), .B(n_53), .Y(n_699) );
OA21x2_ASAP7_75t_L g700 ( .A1(n_542), .A2(n_154), .B(n_215), .Y(n_700) );
OAI21xp5_ASAP7_75t_L g701 ( .A1(n_580), .A2(n_54), .B(n_55), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_SL g702 ( .A1(n_590), .A2(n_157), .B(n_211), .C(n_210), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_536), .B(n_57), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_539), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_571), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_531), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_584), .Y(n_707) );
NOR2xp67_ASAP7_75t_L g708 ( .A(n_579), .B(n_58), .Y(n_708) );
BUFx4_ASAP7_75t_SL g709 ( .A(n_592), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_591), .Y(n_710) );
BUFx4f_ASAP7_75t_L g711 ( .A(n_630), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_687), .A2(n_593), .B(n_552), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_612), .Y(n_713) );
INVx1_ASAP7_75t_SL g714 ( .A(n_669), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_622), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_689), .A2(n_576), .B1(n_583), .B2(n_600), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_667), .Y(n_717) );
BUFx2_ASAP7_75t_L g718 ( .A(n_621), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_617), .A2(n_529), .B(n_540), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_707), .Y(n_720) );
OA21x2_ASAP7_75t_L g721 ( .A1(n_638), .A2(n_168), .B(n_230), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_649), .Y(n_722) );
BUFx2_ASAP7_75t_L g723 ( .A(n_697), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_646), .B(n_59), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_656), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_678), .Y(n_726) );
AO31x2_ASAP7_75t_L g727 ( .A1(n_662), .A2(n_60), .A3(n_61), .B(n_62), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_657), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_616), .A2(n_68), .B1(n_69), .B2(n_129), .Y(n_729) );
OAI22xp33_ASAP7_75t_L g730 ( .A1(n_697), .A2(n_68), .B1(n_69), .B2(n_131), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_642), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_666), .Y(n_732) );
AOI22xp33_ASAP7_75t_SL g733 ( .A1(n_697), .A2(n_666), .B1(n_675), .B2(n_679), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_623), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_657), .A2(n_137), .B1(n_139), .B2(n_141), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_654), .A2(n_170), .B1(n_171), .B2(n_172), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_655), .A2(n_173), .B1(n_174), .B2(n_175), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_672), .B(n_176), .Y(n_738) );
OAI21xp5_ASAP7_75t_L g739 ( .A1(n_617), .A2(n_177), .B(n_178), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_653), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_740) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_675), .A2(n_189), .B1(n_190), .B2(n_194), .Y(n_741) );
INVx6_ASAP7_75t_L g742 ( .A(n_674), .Y(n_742) );
INVx3_ASAP7_75t_L g743 ( .A(n_635), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_624), .B(n_200), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_633), .A2(n_610), .B(n_608), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_613), .A2(n_619), .B(n_632), .Y(n_746) );
OA21x2_ASAP7_75t_L g747 ( .A1(n_640), .A2(n_614), .B(n_634), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_685), .A2(n_692), .B1(n_710), .B2(n_650), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_641), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_668), .A2(n_673), .B1(n_643), .B2(n_681), .Y(n_750) );
AOI211xp5_ASAP7_75t_L g751 ( .A1(n_629), .A2(n_699), .B(n_701), .C(n_620), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_665), .B(n_680), .Y(n_752) );
OAI22xp33_ASAP7_75t_L g753 ( .A1(n_673), .A2(n_701), .B1(n_680), .B2(n_676), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_682), .Y(n_754) );
BUFx12f_ASAP7_75t_L g755 ( .A(n_631), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_708), .A2(n_705), .B1(n_703), .B2(n_676), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_693), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_691), .A2(n_706), .B1(n_659), .B2(n_670), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_618), .A2(n_625), .B(n_702), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_702), .A2(n_690), .B(n_686), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_636), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_627), .A2(n_626), .B1(n_635), .B2(n_695), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_607), .A2(n_615), .B1(n_627), .B2(n_695), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_704), .A2(n_628), .B1(n_664), .B2(n_661), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_696), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_696), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_694), .B(n_704), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_700), .A2(n_647), .B1(n_709), .B2(n_639), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_664), .A2(n_698), .B1(n_647), .B2(n_700), .Y(n_769) );
OR2x6_ASAP7_75t_L g770 ( .A(n_644), .B(n_658), .Y(n_770) );
OAI211xp5_ASAP7_75t_SL g771 ( .A1(n_686), .A2(n_690), .B(n_677), .C(n_694), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_694), .B(n_696), .Y(n_772) );
AOI222xp33_ASAP7_75t_L g773 ( .A1(n_677), .A2(n_694), .B1(n_696), .B2(n_652), .C1(n_651), .C2(n_660), .Y(n_773) );
AOI221xp5_ASAP7_75t_L g774 ( .A1(n_698), .A2(n_677), .B1(n_609), .B2(n_645), .C(n_648), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_677), .Y(n_775) );
INVx6_ASAP7_75t_L g776 ( .A(n_663), .Y(n_776) );
OAI22xp5_ASAP7_75t_SL g777 ( .A1(n_609), .A2(n_671), .B1(n_683), .B2(n_684), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_612), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_687), .A2(n_657), .B1(n_689), .B2(n_688), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_688), .A2(n_570), .B1(n_563), .B2(n_546), .Y(n_780) );
OA21x2_ASAP7_75t_L g781 ( .A1(n_611), .A2(n_638), .B(n_637), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_688), .B(n_689), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_717), .B(n_754), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_765), .Y(n_784) );
BUFx2_ASAP7_75t_L g785 ( .A(n_779), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_733), .B(n_734), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_766), .Y(n_787) );
AND2x2_ASAP7_75t_SL g788 ( .A(n_723), .B(n_748), .Y(n_788) );
INVxp67_ASAP7_75t_L g789 ( .A(n_779), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_772), .Y(n_790) );
OR2x2_ASAP7_75t_L g791 ( .A(n_782), .B(n_714), .Y(n_791) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_714), .Y(n_792) );
INVx3_ASAP7_75t_L g793 ( .A(n_743), .Y(n_793) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_718), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_767), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_757), .B(n_715), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_713), .B(n_722), .Y(n_797) );
OR2x2_ASAP7_75t_L g798 ( .A(n_775), .B(n_780), .Y(n_798) );
INVxp67_ASAP7_75t_L g799 ( .A(n_744), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_727), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_725), .B(n_726), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_727), .Y(n_802) );
BUFx2_ASAP7_75t_L g803 ( .A(n_781), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_727), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_731), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_778), .B(n_720), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_761), .B(n_728), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_728), .B(n_732), .Y(n_808) );
AND2x2_ASAP7_75t_SL g809 ( .A(n_721), .B(n_758), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_773), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_753), .B(n_750), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_750), .B(n_756), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_724), .B(n_751), .Y(n_813) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_752), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_747), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_773), .Y(n_816) );
AND2x4_ASAP7_75t_L g817 ( .A(n_719), .B(n_770), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_735), .B(n_729), .Y(n_818) );
AND2x4_ASAP7_75t_L g819 ( .A(n_770), .B(n_739), .Y(n_819) );
OR2x6_ASAP7_75t_L g820 ( .A(n_762), .B(n_768), .Y(n_820) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_711), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_763), .B(n_716), .Y(n_822) );
INVx3_ASAP7_75t_L g823 ( .A(n_776), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_741), .B(n_737), .Y(n_824) );
OR2x6_ASAP7_75t_L g825 ( .A(n_762), .B(n_760), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_736), .B(n_738), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_774), .B(n_764), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_777), .Y(n_828) );
OR2x2_ASAP7_75t_L g829 ( .A(n_730), .B(n_712), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_771), .Y(n_830) );
INVx4_ASAP7_75t_L g831 ( .A(n_711), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_769), .B(n_745), .Y(n_832) );
BUFx3_ASAP7_75t_L g833 ( .A(n_755), .Y(n_833) );
INVx3_ASAP7_75t_SL g834 ( .A(n_742), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_784), .Y(n_835) );
OR2x2_ASAP7_75t_L g836 ( .A(n_810), .B(n_746), .Y(n_836) );
INVxp67_ASAP7_75t_SL g837 ( .A(n_799), .Y(n_837) );
OR2x2_ASAP7_75t_L g838 ( .A(n_810), .B(n_759), .Y(n_838) );
OR2x2_ASAP7_75t_L g839 ( .A(n_816), .B(n_791), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_815), .Y(n_840) );
AND2x4_ASAP7_75t_L g841 ( .A(n_817), .B(n_740), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_828), .B(n_749), .Y(n_842) );
BUFx2_ASAP7_75t_L g843 ( .A(n_820), .Y(n_843) );
OR2x2_ASAP7_75t_L g844 ( .A(n_798), .B(n_812), .Y(n_844) );
INVx1_ASAP7_75t_SL g845 ( .A(n_792), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_815), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_797), .B(n_801), .Y(n_847) );
INVxp67_ASAP7_75t_L g848 ( .A(n_794), .Y(n_848) );
INVxp67_ASAP7_75t_SL g849 ( .A(n_807), .Y(n_849) );
INVx2_ASAP7_75t_SL g850 ( .A(n_793), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_828), .B(n_830), .Y(n_851) );
INVx3_ASAP7_75t_L g852 ( .A(n_823), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_834), .B(n_831), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_787), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_831), .B(n_814), .Y(n_855) );
BUFx3_ASAP7_75t_L g856 ( .A(n_793), .Y(n_856) );
INVx4_ASAP7_75t_L g857 ( .A(n_820), .Y(n_857) );
OR2x2_ASAP7_75t_L g858 ( .A(n_798), .B(n_795), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_806), .B(n_790), .Y(n_859) );
INVx3_ASAP7_75t_L g860 ( .A(n_823), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_795), .B(n_796), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_796), .B(n_786), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_788), .A2(n_818), .B1(n_813), .B2(n_824), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_786), .B(n_805), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_805), .B(n_827), .Y(n_865) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_833), .B(n_821), .Y(n_866) );
OR2x2_ASAP7_75t_L g867 ( .A(n_785), .B(n_811), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_800), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_783), .B(n_785), .Y(n_869) );
OR2x2_ASAP7_75t_L g870 ( .A(n_839), .B(n_789), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_869), .B(n_804), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_869), .B(n_804), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_840), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_862), .B(n_802), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_862), .B(n_800), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_864), .B(n_802), .Y(n_876) );
OR2x2_ASAP7_75t_L g877 ( .A(n_867), .B(n_829), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_864), .B(n_817), .Y(n_878) );
OR2x2_ASAP7_75t_L g879 ( .A(n_867), .B(n_829), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_859), .B(n_808), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_835), .Y(n_881) );
AND2x2_ASAP7_75t_L g882 ( .A(n_859), .B(n_817), .Y(n_882) );
CKINVDCx14_ASAP7_75t_R g883 ( .A(n_866), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_846), .Y(n_884) );
OR2x2_ASAP7_75t_L g885 ( .A(n_858), .B(n_849), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_865), .B(n_817), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g887 ( .A(n_842), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_865), .B(n_819), .Y(n_888) );
OR2x2_ASAP7_75t_L g889 ( .A(n_858), .B(n_832), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_854), .Y(n_890) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_845), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_861), .B(n_803), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_847), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_836), .B(n_825), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_836), .B(n_825), .Y(n_895) );
INVxp67_ASAP7_75t_L g896 ( .A(n_891), .Y(n_896) );
AOI31xp33_ASAP7_75t_L g897 ( .A1(n_883), .A2(n_853), .A3(n_863), .B(n_855), .Y(n_897) );
OR2x2_ASAP7_75t_L g898 ( .A(n_885), .B(n_844), .Y(n_898) );
OR2x2_ASAP7_75t_L g899 ( .A(n_877), .B(n_838), .Y(n_899) );
OR2x2_ASAP7_75t_L g900 ( .A(n_879), .B(n_843), .Y(n_900) );
OR2x2_ASAP7_75t_L g901 ( .A(n_879), .B(n_843), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_881), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_893), .B(n_851), .Y(n_903) );
OR2x2_ASAP7_75t_L g904 ( .A(n_880), .B(n_848), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_873), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_874), .B(n_857), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_890), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_884), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_875), .B(n_837), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_899), .B(n_876), .Y(n_910) );
AOI21xp33_ASAP7_75t_L g911 ( .A1(n_897), .A2(n_896), .B(n_887), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_899), .B(n_871), .Y(n_912) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_904), .B(n_870), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_902), .Y(n_914) );
NOR3xp33_ASAP7_75t_SL g915 ( .A(n_903), .B(n_832), .C(n_868), .Y(n_915) );
NAND4xp25_ASAP7_75t_SL g916 ( .A(n_906), .B(n_882), .C(n_888), .D(n_878), .Y(n_916) );
O2A1O1Ixp33_ASAP7_75t_L g917 ( .A1(n_911), .A2(n_898), .B(n_909), .C(n_907), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_916), .A2(n_895), .B1(n_894), .B2(n_913), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_914), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_919), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_918), .A2(n_915), .B1(n_912), .B2(n_910), .Y(n_921) );
O2A1O1Ixp33_ASAP7_75t_L g922 ( .A1(n_917), .A2(n_826), .B(n_900), .C(n_901), .Y(n_922) );
O2A1O1Ixp33_ASAP7_75t_L g923 ( .A1(n_921), .A2(n_850), .B(n_822), .C(n_889), .Y(n_923) );
OAI221xp5_ASAP7_75t_SL g924 ( .A1(n_922), .A2(n_889), .B1(n_886), .B2(n_872), .C(n_892), .Y(n_924) );
OR2x2_ASAP7_75t_L g925 ( .A(n_924), .B(n_920), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_923), .B(n_908), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_926), .Y(n_927) );
INVx2_ASAP7_75t_L g928 ( .A(n_925), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_928), .A2(n_841), .B1(n_905), .B2(n_809), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_927), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_930), .Y(n_931) );
OAI22xp5_ASAP7_75t_SL g932 ( .A1(n_931), .A2(n_929), .B1(n_809), .B2(n_856), .Y(n_932) );
AOI21xp5_ASAP7_75t_L g933 ( .A1(n_932), .A2(n_783), .B(n_850), .Y(n_933) );
INVxp67_ASAP7_75t_L g934 ( .A(n_933), .Y(n_934) );
AOI21xp5_ASAP7_75t_L g935 ( .A1(n_934), .A2(n_852), .B(n_860), .Y(n_935) );
endmodule