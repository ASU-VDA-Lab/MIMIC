module fake_jpeg_26587_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx5_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_11),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_10),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_30),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_18),
.B1(n_15),
.B2(n_14),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_29),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_16),
.B1(n_13),
.B2(n_12),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_11),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_23),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_23),
.B(n_2),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_39),
.B(n_0),
.Y(n_46)
);

CKINVDCx12_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_32),
.B(n_8),
.C(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_6),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_33),
.C(n_35),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_33),
.Y(n_47)
);

OAI221xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_42),
.C(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_50),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_40),
.B1(n_22),
.B2(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_53),
.Y(n_55)
);

NOR2xp67_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_40),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_55),
.C(n_7),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_3),
.B(n_0),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_2),
.Y(n_60)
);


endmodule