module fake_jpeg_16792_n_217 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_217);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NAND2x1_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_0),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_28),
.A2(n_17),
.B(n_24),
.C(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_37),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

HAxp5_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_26),
.CON(n_38),
.SN(n_38)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_47),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_21),
.B1(n_27),
.B2(n_20),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_42),
.B1(n_52),
.B2(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_25),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_49),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_30),
.A2(n_14),
.B1(n_17),
.B2(n_20),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_20),
.B1(n_15),
.B2(n_22),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_66),
.Y(n_79)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_70),
.Y(n_81)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_69),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_22),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_34),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_9),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_49),
.A3(n_42),
.B1(n_39),
.B2(n_52),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_22),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_49),
.B(n_47),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_77),
.B(n_85),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_45),
.B1(n_48),
.B2(n_43),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_86),
.B1(n_67),
.B2(n_60),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_1),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_88),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_54),
.C(n_31),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_62),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_34),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_102),
.B(n_105),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_100),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_76),
.Y(n_119)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_101),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_1),
.B(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_55),
.B1(n_68),
.B2(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_76),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_102),
.A2(n_94),
.B(n_82),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_112),
.B(n_119),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_86),
.B(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_111),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_81),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_123),
.C(n_100),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_77),
.B(n_89),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_120),
.B(n_121),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_77),
.B(n_72),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_88),
.B(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_87),
.C(n_76),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_76),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_55),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_97),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_122),
.A2(n_91),
.B1(n_96),
.B2(n_107),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_137),
.B1(n_140),
.B2(n_123),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_119),
.A2(n_92),
.B1(n_105),
.B2(n_103),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_111),
.B(n_108),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_138),
.C(n_118),
.Y(n_144)
);

AO22x2_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_101),
.B1(n_106),
.B2(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_134),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_57),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_106),
.B1(n_57),
.B2(n_37),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_15),
.Y(n_141)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_6),
.C(n_2),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_11),
.C(n_2),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_152),
.C(n_154),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_130),
.C(n_142),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_158),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_118),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_129),
.B(n_128),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_149),
.A2(n_131),
.B1(n_132),
.B2(n_139),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_161),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_127),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_166),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_132),
.B1(n_158),
.B2(n_153),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_169),
.B1(n_170),
.B2(n_159),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_115),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_165),
.B(n_167),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_139),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_131),
.B1(n_152),
.B2(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_109),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_144),
.C(n_155),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_177),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_129),
.C(n_154),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_180),
.B(n_178),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_121),
.C(n_117),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_173),
.C(n_168),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_179),
.B(n_181),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_140),
.C(n_145),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_161),
.C(n_170),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_184),
.Y(n_190)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_7),
.C(n_3),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_192),
.B(n_195),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_160),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_4),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_202),
.B(n_10),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_5),
.B(n_6),
.Y(n_199)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_7),
.B(n_8),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_201),
.A2(n_195),
.B(n_190),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_8),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_194),
.B(n_8),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_207),
.B(n_201),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_200),
.B1(n_198),
.B2(n_191),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_208),
.Y(n_209)
);

AOI31xp67_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_211),
.A3(n_11),
.B(n_13),
.Y(n_214)
);

AO21x1_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_10),
.B(n_11),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_213),
.A2(n_214),
.B(n_212),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_215),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_208),
.Y(n_217)
);


endmodule