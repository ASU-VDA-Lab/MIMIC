module fake_jpeg_9720_n_259 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_259);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_259;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_6),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_45),
.Y(n_53)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_27),
.B1(n_20),
.B2(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_40),
.B(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_0),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_43),
.C(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_17),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_2),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_2),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_52),
.Y(n_80)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_57),
.B(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_44),
.B(n_27),
.Y(n_76)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_46),
.B1(n_39),
.B2(n_44),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_38),
.B(n_24),
.C(n_21),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_76),
.A2(n_25),
.B(n_22),
.Y(n_115)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_82),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_44),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_25),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_36),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_36),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_27),
.B1(n_21),
.B2(n_22),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_92),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_60),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_49),
.A2(n_37),
.B1(n_36),
.B2(n_38),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_47),
.B1(n_37),
.B2(n_70),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_37),
.B1(n_47),
.B2(n_51),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_95),
.A2(n_116),
.B1(n_71),
.B2(n_79),
.Y(n_142)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_48),
.A3(n_51),
.B1(n_65),
.B2(n_55),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_103),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_65),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_113),
.C(n_73),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_47),
.B1(n_67),
.B2(n_69),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_105),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_69),
.B1(n_61),
.B2(n_38),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_62),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_54),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_110),
.B(n_93),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_25),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_57),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_25),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_20),
.B(n_77),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_69),
.B1(n_38),
.B2(n_56),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_92),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_118),
.A2(n_93),
.B(n_85),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_76),
.B1(n_95),
.B2(n_115),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_142),
.B1(n_118),
.B2(n_99),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_122),
.B(n_134),
.Y(n_151)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_127),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_84),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_81),
.C(n_73),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_31),
.Y(n_165)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_72),
.B(n_78),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_138),
.B(n_143),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_89),
.B1(n_72),
.B2(n_83),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_112),
.B1(n_105),
.B2(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_137),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_139),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_83),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_147),
.B1(n_159),
.B2(n_136),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_100),
.B1(n_77),
.B2(n_71),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_114),
.B1(n_109),
.B2(n_110),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_153),
.B(n_155),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_162),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_110),
.B1(n_109),
.B2(n_96),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_98),
.B(n_107),
.C(n_31),
.D(n_23),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_90),
.Y(n_156)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_71),
.B1(n_18),
.B2(n_34),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_90),
.Y(n_162)
);

NOR2x1_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_33),
.Y(n_163)
);

NAND2x1_ASAP7_75t_SL g184 ( 
.A(n_163),
.B(n_23),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_164),
.A2(n_29),
.B1(n_19),
.B2(n_18),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_124),
.C(n_128),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_31),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_166),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_3),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_134),
.B(n_131),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_169),
.A2(n_173),
.B1(n_174),
.B2(n_189),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_171),
.B(n_145),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_180),
.C(n_187),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_137),
.B1(n_135),
.B2(n_130),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_127),
.B1(n_123),
.B2(n_32),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_31),
.Y(n_177)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_29),
.C(n_19),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_181),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_3),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_152),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_185),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_161),
.B1(n_164),
.B2(n_167),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_23),
.C(n_4),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_151),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_188),
.A2(n_144),
.B(n_166),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_23),
.B1(n_5),
.B2(n_6),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_162),
.C(n_165),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_170),
.C(n_178),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_194),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_171),
.A2(n_146),
.B(n_167),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_205),
.B(n_189),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_146),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_187),
.B(n_9),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_155),
.C(n_153),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_183),
.B1(n_176),
.B2(n_182),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_208),
.B1(n_184),
.B2(n_180),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_174),
.Y(n_212)
);

AO22x1_ASAP7_75t_SL g205 ( 
.A1(n_190),
.A2(n_148),
.B1(n_5),
.B2(n_6),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_173),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_221),
.C(n_193),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g211 ( 
.A(n_197),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_222),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_202),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_183),
.B(n_182),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_220),
.B(n_205),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_204),
.A2(n_181),
.B1(n_184),
.B2(n_186),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_217),
.A2(n_218),
.B1(n_194),
.B2(n_201),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_206),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_179),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

AO22x1_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_205),
.B1(n_203),
.B2(n_196),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_SL g237 ( 
.A1(n_223),
.A2(n_218),
.B(n_209),
.C(n_213),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_228),
.B1(n_7),
.B2(n_9),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_233),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_192),
.C(n_191),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_230),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_213),
.C(n_216),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_231),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_192),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_212),
.Y(n_234)
);

A2O1A1O1Ixp25_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_227),
.B(n_233),
.C(n_229),
.D(n_223),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_237),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_230),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_7),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_241),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_9),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_244),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_245),
.B(n_13),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_246),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_16),
.B(n_249),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_236),
.B(n_237),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_235),
.C(n_242),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_253),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_254),
.A2(n_255),
.B(n_16),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_248),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_16),
.B(n_255),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_257),
.Y(n_259)
);


endmodule