module fake_ariane_1857_n_1245 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1245);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1245;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_187;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_232;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_200;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_238;
wire n_365;
wire n_1013;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_461;
wire n_1121;
wire n_209;
wire n_490;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_555;
wire n_804;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_179;
wire n_1178;
wire n_1026;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_564;
wire n_205;
wire n_1029;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_233;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_888;
wire n_845;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_642;
wire n_211;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_197;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_272;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_181;
wire n_617;
wire n_543;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_243;
wire n_185;
wire n_1204;
wire n_994;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_385;
wire n_917;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_174;
wire n_275;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_250;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_84),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_16),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_86),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_160),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_128),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_15),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_113),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_136),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_125),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_163),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_153),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_9),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_8),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_91),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_138),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_60),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_137),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_76),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_69),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_127),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_146),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_61),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_66),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_107),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_12),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_135),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_6),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_29),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_157),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_151),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_42),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_126),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_134),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_18),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_149),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_22),
.Y(n_206)
);

BUFx8_ASAP7_75t_SL g207 ( 
.A(n_54),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_121),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_89),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_122),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_156),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_147),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_3),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_8),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_130),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_46),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_58),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_108),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_123),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_49),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_164),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_77),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_103),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_43),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_4),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_80),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_85),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_16),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_150),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_34),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_23),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_55),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_57),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_73),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_133),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_4),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_14),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_131),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_129),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_21),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_42),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_96),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_115),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_140),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_59),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_35),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_98),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_71),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_148),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_82),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_14),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_124),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_62),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_152),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_26),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_97),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_93),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_114),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_83),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_90),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_56),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_38),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_13),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_99),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_144),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_145),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_47),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_36),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_143),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_26),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_34),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_6),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_81),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_23),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_36),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_95),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_32),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_72),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_67),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_22),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_112),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_19),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_40),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_207),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_223),
.B(n_0),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_193),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_239),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_284),
.Y(n_292)
);

INVxp33_ASAP7_75t_SL g293 ( 
.A(n_267),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_239),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_167),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_167),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_284),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_171),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_168),
.B(n_0),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_167),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_207),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_167),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_167),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_166),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_196),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_167),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_179),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_167),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_238),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_238),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_238),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_176),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_238),
.Y(n_313)
);

INVxp33_ASAP7_75t_SL g314 ( 
.A(n_180),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_179),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_245),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_238),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_257),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_238),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g320 ( 
.A(n_181),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_218),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_238),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_172),
.B(n_1),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_199),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_257),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_245),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_204),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_283),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_283),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_206),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_243),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_248),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_283),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_195),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_173),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_213),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_203),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_209),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_208),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_222),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_R g343 ( 
.A(n_165),
.B(n_169),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_224),
.Y(n_344)
);

BUFx6f_ASAP7_75t_SL g345 ( 
.A(n_218),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_214),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_228),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_235),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_235),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_265),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_265),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_226),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_229),
.B(n_231),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_237),
.B(n_1),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_246),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_227),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_230),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_250),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_251),
.B(n_2),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g360 ( 
.A(n_232),
.B(n_2),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_233),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_L g362 ( 
.A(n_242),
.B(n_253),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_201),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_277),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_254),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_261),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_262),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_264),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_270),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_272),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_277),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_268),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_273),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_269),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_279),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_275),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_337),
.B(n_339),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_304),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_295),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_296),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_300),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_304),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_312),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_300),
.Y(n_384)
);

OAI21x1_ASAP7_75t_L g385 ( 
.A1(n_303),
.A2(n_201),
.B(n_281),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_304),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_321),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_321),
.B(n_185),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_348),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_302),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_306),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_308),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_215),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_349),
.B(n_363),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_340),
.B(n_187),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_309),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_348),
.B(n_166),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_292),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_303),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_310),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_304),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_311),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_304),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_313),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_317),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_319),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_338),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_353),
.B(n_221),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_370),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_342),
.B(n_170),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_344),
.B(n_166),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_365),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_365),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_347),
.B(n_174),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_376),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_355),
.B(n_166),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_358),
.B(n_175),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_366),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_372),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_324),
.Y(n_425)
);

NAND2xp33_ASAP7_75t_SL g426 ( 
.A(n_292),
.B(n_285),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_327),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_290),
.B(n_177),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_359),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_331),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_333),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_305),
.B(n_178),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_334),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_287),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_289),
.B(n_182),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_299),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_323),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_332),
.B(n_183),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_293),
.B(n_184),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_293),
.A2(n_280),
.B1(n_278),
.B2(n_271),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_354),
.A2(n_258),
.B(n_188),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_330),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_288),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_329),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_297),
.B(n_186),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_345),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_395),
.B(n_297),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_407),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_437),
.A2(n_320),
.B1(n_314),
.B2(n_346),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_381),
.Y(n_451)
);

CKINVDCx6p67_ASAP7_75t_R g452 ( 
.A(n_444),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_436),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_395),
.B(n_298),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_407),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_384),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_384),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_379),
.B(n_328),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_407),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_400),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_429),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_400),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_379),
.B(n_328),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_400),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_405),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_314),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_399),
.B(n_301),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_410),
.A2(n_439),
.B1(n_437),
.B2(n_443),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_405),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_445),
.B(n_335),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_383),
.B(n_291),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_445),
.B(n_335),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_380),
.B(n_258),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_389),
.B(n_320),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_383),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_395),
.B(n_373),
.Y(n_479)
);

OAI22xp33_ASAP7_75t_L g480 ( 
.A1(n_410),
.A2(n_437),
.B1(n_443),
.B2(n_442),
.Y(n_480)
);

AND2x2_ASAP7_75t_SL g481 ( 
.A(n_436),
.B(n_315),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_380),
.B(n_258),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_442),
.B(n_425),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_407),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_406),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_406),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_436),
.A2(n_346),
.B1(n_360),
.B2(n_345),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_409),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_445),
.B(n_356),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_436),
.A2(n_345),
.B1(n_356),
.B2(n_368),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_409),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_390),
.B(n_258),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_409),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_407),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_390),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_440),
.B(n_357),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_387),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_436),
.A2(n_361),
.B1(n_357),
.B2(n_368),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_391),
.Y(n_502)
);

INVx6_ASAP7_75t_L g503 ( 
.A(n_398),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_429),
.B(n_258),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_399),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_391),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_392),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_389),
.B(n_361),
.Y(n_508)
);

NAND3xp33_ASAP7_75t_L g509 ( 
.A(n_436),
.B(n_352),
.C(n_336),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_378),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_392),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_378),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_396),
.B(n_258),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_436),
.A2(n_362),
.B1(n_375),
.B2(n_258),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_396),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_440),
.B(n_343),
.Y(n_516)
);

NAND3xp33_ASAP7_75t_SL g517 ( 
.A(n_432),
.B(n_301),
.C(n_286),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_471),
.B(n_419),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_471),
.B(n_419),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_511),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_450),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_480),
.B(n_419),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_480),
.B(n_501),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_469),
.B(n_429),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_500),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_455),
.B(n_326),
.Y(n_526)
);

AO221x1_ASAP7_75t_L g527 ( 
.A1(n_505),
.A2(n_399),
.B1(n_408),
.B2(n_429),
.C(n_307),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_501),
.B(n_429),
.Y(n_528)
);

NOR2x1p5_ASAP7_75t_L g529 ( 
.A(n_452),
.B(n_307),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_450),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_509),
.A2(n_435),
.B1(n_429),
.B2(n_428),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_461),
.B(n_429),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_500),
.Y(n_533)
);

NAND3xp33_ASAP7_75t_L g534 ( 
.A(n_449),
.B(n_408),
.C(n_397),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_484),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_464),
.B(n_397),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_484),
.B(n_389),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_477),
.B(n_428),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_464),
.B(n_411),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_450),
.Y(n_540)
);

NOR2xp67_ASAP7_75t_SL g541 ( 
.A(n_492),
.B(n_411),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_511),
.Y(n_542)
);

NAND3xp33_ASAP7_75t_L g543 ( 
.A(n_505),
.B(n_432),
.C(n_426),
.Y(n_543)
);

INVx8_ASAP7_75t_L g544 ( 
.A(n_504),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_461),
.B(n_428),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_455),
.B(n_444),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_498),
.A2(n_415),
.B1(n_417),
.B2(n_420),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_498),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_479),
.B(n_442),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_498),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_L g551 ( 
.A(n_478),
.B(n_446),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_464),
.B(n_401),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_502),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_465),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_466),
.B(n_428),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_466),
.B(n_428),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_465),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_479),
.B(n_438),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_465),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_467),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_464),
.B(n_401),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_502),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_509),
.B(n_453),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_453),
.B(n_438),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_453),
.B(n_438),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_493),
.B(n_403),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_458),
.B(n_403),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_467),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_447),
.B(n_387),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_458),
.B(n_438),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_467),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_458),
.B(n_438),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_502),
.Y(n_573)
);

A2O1A1Ixp33_ASAP7_75t_L g574 ( 
.A1(n_506),
.A2(n_441),
.B(n_515),
.C(n_507),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_516),
.A2(n_435),
.B1(n_416),
.B2(n_412),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_447),
.B(n_435),
.Y(n_576)
);

NOR2xp67_ASAP7_75t_SL g577 ( 
.A(n_473),
.B(n_425),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_474),
.Y(n_578)
);

NOR2x1p5_ASAP7_75t_L g579 ( 
.A(n_452),
.B(n_316),
.Y(n_579)
);

BUFx8_ASAP7_75t_L g580 ( 
.A(n_452),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_474),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_497),
.A2(n_416),
.B(n_412),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_490),
.B(n_506),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_506),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_507),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_490),
.B(n_422),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_507),
.B(n_422),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_515),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_458),
.B(n_481),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_458),
.B(n_431),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_515),
.Y(n_591)
);

OAI221xp5_ASAP7_75t_L g592 ( 
.A1(n_499),
.A2(n_434),
.B1(n_422),
.B2(n_430),
.C(n_424),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_481),
.B(n_341),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_468),
.Y(n_594)
);

O2A1O1Ixp33_ASAP7_75t_L g595 ( 
.A1(n_468),
.A2(n_425),
.B(n_430),
.C(n_423),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_472),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_487),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_472),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_514),
.B(n_426),
.C(n_316),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_487),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_487),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_475),
.B(n_364),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_485),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_514),
.B(n_387),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_481),
.A2(n_388),
.B1(n_424),
.B2(n_421),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_489),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_470),
.B(n_341),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_503),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_503),
.B(n_394),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_485),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_517),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_503),
.B(n_394),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_458),
.B(n_431),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_488),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_503),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_488),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_582),
.A2(n_532),
.B(n_535),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_529),
.Y(n_618)
);

BUFx4f_ASAP7_75t_L g619 ( 
.A(n_569),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_524),
.B(n_425),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_520),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_615),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_524),
.B(n_425),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_556),
.B(n_377),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_556),
.B(n_377),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_538),
.B(n_609),
.Y(n_626)
);

BUFx12f_ASAP7_75t_L g627 ( 
.A(n_580),
.Y(n_627)
);

AOI21xp33_ASAP7_75t_L g628 ( 
.A1(n_522),
.A2(n_496),
.B(n_494),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_532),
.A2(n_441),
.B(n_494),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_609),
.B(n_612),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_552),
.A2(n_497),
.B(n_462),
.Y(n_631)
);

AO21x1_ASAP7_75t_L g632 ( 
.A1(n_523),
.A2(n_483),
.B(n_476),
.Y(n_632)
);

AND3x1_ASAP7_75t_L g633 ( 
.A(n_546),
.B(n_576),
.C(n_558),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_612),
.B(n_377),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_542),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_545),
.B(n_503),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_616),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_594),
.Y(n_638)
);

OAI21xp33_ASAP7_75t_L g639 ( 
.A1(n_555),
.A2(n_517),
.B(n_423),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_552),
.A2(n_497),
.B(n_462),
.Y(n_640)
);

NOR3xp33_ASAP7_75t_L g641 ( 
.A(n_534),
.B(n_421),
.C(n_434),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_549),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_526),
.B(n_291),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_559),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_543),
.B(n_608),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_561),
.A2(n_462),
.B(n_448),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_561),
.A2(n_462),
.B(n_448),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_564),
.A2(n_482),
.B(n_448),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_559),
.Y(n_649)
);

CKINVDCx10_ASAP7_75t_R g650 ( 
.A(n_578),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_523),
.B(n_448),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_544),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_565),
.A2(n_441),
.B(n_496),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_L g654 ( 
.A1(n_574),
.A2(n_491),
.B(n_489),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_574),
.A2(n_491),
.B(n_489),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_518),
.B(n_500),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_595),
.A2(n_491),
.B(n_483),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_567),
.A2(n_486),
.B(n_482),
.Y(n_658)
);

AOI21x1_ASAP7_75t_L g659 ( 
.A1(n_589),
.A2(n_495),
.B(n_476),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_519),
.B(n_388),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_575),
.B(n_388),
.Y(n_661)
);

O2A1O1Ixp5_ASAP7_75t_L g662 ( 
.A1(n_577),
.A2(n_482),
.B(n_486),
.C(n_513),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_531),
.B(n_388),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_567),
.A2(n_486),
.B(n_482),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_536),
.A2(n_513),
.B(n_495),
.C(n_486),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_537),
.B(n_388),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_593),
.B(n_446),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_580),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_525),
.Y(n_669)
);

OAI21xp33_ASAP7_75t_L g670 ( 
.A1(n_536),
.A2(n_393),
.B(n_413),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_569),
.B(n_413),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_581),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_596),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_615),
.B(n_456),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_539),
.B(n_451),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_560),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_548),
.A2(n_454),
.B(n_451),
.Y(n_677)
);

O2A1O1Ixp5_ASAP7_75t_L g678 ( 
.A1(n_528),
.A2(n_510),
.B(n_459),
.C(n_454),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_598),
.A2(n_456),
.B1(n_460),
.B2(n_463),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_590),
.A2(n_456),
.B(n_510),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_539),
.B(n_457),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_570),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_590),
.A2(n_613),
.B(n_563),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_602),
.B(n_294),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_605),
.B(n_413),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_607),
.B(n_294),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_611),
.B(n_550),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_613),
.A2(n_510),
.B(n_459),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_553),
.A2(n_460),
.B(n_457),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_579),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_603),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_563),
.A2(n_510),
.B(n_463),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_562),
.A2(n_504),
.B(n_385),
.Y(n_693)
);

O2A1O1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_570),
.A2(n_427),
.B(n_393),
.C(n_414),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_599),
.A2(n_415),
.B1(n_417),
.B2(n_414),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_572),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_610),
.A2(n_614),
.B1(n_572),
.B2(n_573),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_584),
.B(n_418),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_551),
.B(n_427),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_585),
.B(n_418),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_587),
.A2(n_427),
.B(n_420),
.C(n_418),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_588),
.A2(n_591),
.B(n_544),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_586),
.B(n_597),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_525),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_528),
.A2(n_398),
.B(n_417),
.C(n_415),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_597),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_583),
.A2(n_431),
.B1(n_433),
.B2(n_318),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_592),
.B(n_431),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_541),
.Y(n_709)
);

O2A1O1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_566),
.A2(n_398),
.B(n_404),
.C(n_402),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_566),
.A2(n_398),
.B(n_404),
.C(n_402),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_533),
.B(n_398),
.Y(n_712)
);

O2A1O1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_600),
.A2(n_402),
.B(n_404),
.C(n_351),
.Y(n_713)
);

OAI321xp33_ASAP7_75t_L g714 ( 
.A1(n_604),
.A2(n_433),
.A3(n_431),
.B1(n_325),
.B2(n_350),
.C(n_351),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_R g715 ( 
.A(n_672),
.B(n_690),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_654),
.A2(n_385),
.B(n_600),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_644),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_644),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_686),
.B(n_318),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_652),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_643),
.B(n_325),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_630),
.A2(n_544),
.B1(n_547),
.B2(n_533),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_619),
.B(n_589),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_621),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_642),
.B(n_601),
.Y(n_725)
);

OAI22x1_ASAP7_75t_L g726 ( 
.A1(n_684),
.A2(n_371),
.B1(n_350),
.B2(n_527),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_619),
.B(n_601),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_626),
.A2(n_639),
.B(n_645),
.C(n_625),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_633),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_624),
.A2(n_547),
.B1(n_606),
.B2(n_560),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_635),
.Y(n_731)
);

OAI21xp33_ASAP7_75t_L g732 ( 
.A1(n_634),
.A2(n_371),
.B(n_606),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_660),
.B(n_637),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_704),
.A2(n_645),
.B1(n_696),
.B2(n_682),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_617),
.A2(n_571),
.B(n_530),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_620),
.A2(n_568),
.B(n_540),
.Y(n_736)
);

A2O1A1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_675),
.A2(n_557),
.B(n_554),
.C(n_521),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_709),
.B(n_431),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_675),
.A2(n_385),
.B(n_433),
.C(n_431),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_623),
.A2(n_512),
.B(n_190),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_649),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_682),
.A2(n_504),
.B1(n_433),
.B2(n_236),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_629),
.A2(n_512),
.B(n_191),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_649),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_636),
.A2(n_433),
.B1(n_189),
.B2(n_225),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_638),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_676),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_655),
.A2(n_512),
.B(n_433),
.Y(n_748)
);

BUFx8_ASAP7_75t_L g749 ( 
.A(n_627),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_673),
.B(n_691),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_SL g751 ( 
.A1(n_627),
.A2(n_192),
.B1(n_194),
.B2(n_197),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_687),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_656),
.B(n_504),
.Y(n_753)
);

OAI21xp33_ASAP7_75t_SL g754 ( 
.A1(n_666),
.A2(n_504),
.B(n_5),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_667),
.B(n_433),
.Y(n_755)
);

BUFx8_ASAP7_75t_L g756 ( 
.A(n_668),
.Y(n_756)
);

BUFx12f_ASAP7_75t_L g757 ( 
.A(n_618),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_709),
.A2(n_504),
.B1(n_244),
.B2(n_241),
.Y(n_758)
);

OAI21xp5_ASAP7_75t_L g759 ( 
.A1(n_651),
.A2(n_504),
.B(n_512),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_697),
.A2(n_3),
.B(n_5),
.C(n_7),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_671),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_702),
.A2(n_512),
.B(n_247),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_701),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_669),
.B(n_198),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_676),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_706),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_653),
.A2(n_512),
.B(n_249),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_681),
.A2(n_504),
.B(n_240),
.C(n_234),
.Y(n_768)
);

OA21x2_ASAP7_75t_L g769 ( 
.A1(n_693),
.A2(n_252),
.B(n_202),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_669),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_R g771 ( 
.A(n_650),
.B(n_200),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_699),
.B(n_714),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_641),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_651),
.A2(n_11),
.B(n_13),
.C(n_15),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_652),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_622),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_683),
.A2(n_512),
.B(n_255),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_712),
.Y(n_778)
);

BUFx12f_ASAP7_75t_L g779 ( 
.A(n_618),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_659),
.A2(n_116),
.B(n_161),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_622),
.B(n_205),
.Y(n_781)
);

BUFx10_ASAP7_75t_L g782 ( 
.A(n_721),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_728),
.A2(n_708),
.B(n_679),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_748),
.A2(n_708),
.B(n_657),
.Y(n_784)
);

NOR2xp67_ASAP7_75t_L g785 ( 
.A(n_752),
.B(n_757),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_719),
.B(n_641),
.Y(n_786)
);

BUFx4f_ASAP7_75t_L g787 ( 
.A(n_779),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_733),
.B(n_681),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_724),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_729),
.B(n_712),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_733),
.B(n_685),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_778),
.Y(n_792)
);

BUFx10_ASAP7_75t_L g793 ( 
.A(n_770),
.Y(n_793)
);

AOI221x1_ASAP7_75t_L g794 ( 
.A1(n_726),
.A2(n_707),
.B1(n_661),
.B2(n_628),
.C(n_670),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_770),
.Y(n_795)
);

NAND3x1_ASAP7_75t_L g796 ( 
.A(n_734),
.B(n_663),
.C(n_700),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_SL g797 ( 
.A1(n_781),
.A2(n_674),
.B(n_665),
.C(n_698),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_749),
.Y(n_798)
);

AOI221xp5_ASAP7_75t_SL g799 ( 
.A1(n_760),
.A2(n_694),
.B1(n_648),
.B2(n_692),
.C(n_647),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_750),
.A2(n_677),
.B1(n_689),
.B2(n_695),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_748),
.A2(n_688),
.B(n_680),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_731),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_746),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_720),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_739),
.A2(n_662),
.B(n_632),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_L g806 ( 
.A(n_770),
.B(n_646),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_750),
.B(n_695),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_773),
.B(n_658),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_766),
.Y(n_809)
);

OAI21x1_ASAP7_75t_L g810 ( 
.A1(n_716),
.A2(n_678),
.B(n_703),
.Y(n_810)
);

NAND2x1_ASAP7_75t_L g811 ( 
.A(n_720),
.B(n_664),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_717),
.Y(n_812)
);

AOI31xp67_ASAP7_75t_L g813 ( 
.A1(n_753),
.A2(n_674),
.A3(n_711),
.B(n_710),
.Y(n_813)
);

INVx5_ASAP7_75t_L g814 ( 
.A(n_775),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_718),
.Y(n_815)
);

AO31x2_ASAP7_75t_L g816 ( 
.A1(n_730),
.A2(n_640),
.A3(n_631),
.B(n_705),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_735),
.A2(n_713),
.B(n_386),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_763),
.A2(n_256),
.B(n_211),
.C(n_212),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_753),
.A2(n_259),
.B(n_216),
.Y(n_819)
);

AO31x2_ASAP7_75t_L g820 ( 
.A1(n_730),
.A2(n_386),
.A3(n_382),
.B(n_378),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_722),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_722),
.A2(n_386),
.B(n_382),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_741),
.Y(n_823)
);

OAI21x1_ASAP7_75t_L g824 ( 
.A1(n_780),
.A2(n_386),
.B(n_382),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_755),
.A2(n_260),
.B(n_217),
.C(n_219),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_774),
.A2(n_266),
.B(n_263),
.C(n_220),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_732),
.A2(n_210),
.B1(n_382),
.B2(n_378),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_744),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_725),
.B(n_17),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_725),
.B(n_20),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_715),
.A2(n_751),
.B1(n_723),
.B2(n_727),
.Y(n_831)
);

OAI221xp5_ASAP7_75t_L g832 ( 
.A1(n_761),
.A2(n_386),
.B1(n_382),
.B2(n_378),
.C(n_25),
.Y(n_832)
);

NOR2x1_ASAP7_75t_SL g833 ( 
.A(n_738),
.B(n_764),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_736),
.A2(n_386),
.B(n_382),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_743),
.A2(n_386),
.B(n_382),
.Y(n_835)
);

OR2x6_ASAP7_75t_L g836 ( 
.A(n_723),
.B(n_775),
.Y(n_836)
);

OA21x2_ASAP7_75t_L g837 ( 
.A1(n_759),
.A2(n_378),
.B(n_102),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_776),
.B(n_378),
.Y(n_838)
);

OA21x2_ASAP7_75t_L g839 ( 
.A1(n_759),
.A2(n_101),
.B(n_158),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_789),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_812),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_786),
.A2(n_756),
.B1(n_772),
.B2(n_749),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_790),
.A2(n_756),
.B1(n_758),
.B2(n_742),
.Y(n_843)
);

INVx6_ASAP7_75t_L g844 ( 
.A(n_793),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_795),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_815),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_787),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_821),
.A2(n_769),
.B1(n_747),
.B2(n_765),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_798),
.Y(n_849)
);

BUFx8_ASAP7_75t_SL g850 ( 
.A(n_787),
.Y(n_850)
);

CKINVDCx11_ASAP7_75t_R g851 ( 
.A(n_782),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_802),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_823),
.Y(n_853)
);

INVx6_ASAP7_75t_L g854 ( 
.A(n_793),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_782),
.Y(n_855)
);

CKINVDCx14_ASAP7_75t_R g856 ( 
.A(n_830),
.Y(n_856)
);

CKINVDCx11_ASAP7_75t_R g857 ( 
.A(n_803),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_821),
.A2(n_832),
.B1(n_791),
.B2(n_788),
.Y(n_858)
);

INVx5_ASAP7_75t_L g859 ( 
.A(n_836),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_792),
.Y(n_860)
);

OAI22x1_ASAP7_75t_L g861 ( 
.A1(n_831),
.A2(n_809),
.B1(n_788),
.B2(n_829),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_828),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_836),
.Y(n_863)
);

BUFx2_ASAP7_75t_R g864 ( 
.A(n_791),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_832),
.A2(n_769),
.B1(n_745),
.B2(n_754),
.Y(n_865)
);

BUFx8_ASAP7_75t_SL g866 ( 
.A(n_836),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_807),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_827),
.A2(n_745),
.B1(n_771),
.B2(n_776),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_785),
.B(n_737),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_796),
.B(n_20),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_814),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_800),
.A2(n_740),
.B1(n_767),
.B2(n_777),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_800),
.A2(n_768),
.B1(n_762),
.B2(n_25),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_808),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_SL g875 ( 
.A1(n_833),
.A2(n_21),
.B1(n_24),
.B2(n_27),
.Y(n_875)
);

INVx6_ASAP7_75t_L g876 ( 
.A(n_814),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_820),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_814),
.Y(n_878)
);

CKINVDCx11_ASAP7_75t_R g879 ( 
.A(n_806),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_814),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_783),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_881)
);

CKINVDCx11_ASAP7_75t_R g882 ( 
.A(n_794),
.Y(n_882)
);

INVx4_ASAP7_75t_L g883 ( 
.A(n_804),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_804),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_838),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_811),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_819),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_797),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_813),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_816),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_820),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_SL g892 ( 
.A1(n_839),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_839),
.Y(n_893)
);

INVx5_ASAP7_75t_L g894 ( 
.A(n_837),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_819),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_837),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_816),
.Y(n_897)
);

CKINVDCx6p67_ASAP7_75t_R g898 ( 
.A(n_818),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_799),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_816),
.Y(n_900)
);

OAI21x1_ASAP7_75t_L g901 ( 
.A1(n_893),
.A2(n_801),
.B(n_835),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_891),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_890),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_891),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_897),
.B(n_820),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_900),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_886),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_889),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_874),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_850),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_886),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_877),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_877),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_893),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_894),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_894),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_894),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_894),
.Y(n_918)
);

AO21x2_ASAP7_75t_L g919 ( 
.A1(n_888),
.A2(n_822),
.B(n_805),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_872),
.A2(n_801),
.B(n_835),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_899),
.B(n_822),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_899),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_840),
.B(n_805),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_852),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_867),
.Y(n_925)
);

OAI21x1_ASAP7_75t_L g926 ( 
.A1(n_872),
.A2(n_834),
.B(n_784),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_862),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_892),
.B(n_810),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_841),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_841),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_896),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_848),
.B(n_799),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_863),
.B(n_817),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_853),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_878),
.B(n_824),
.Y(n_935)
);

AO21x1_ASAP7_75t_L g936 ( 
.A1(n_870),
.A2(n_826),
.B(n_825),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_853),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_880),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_884),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_880),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_922),
.A2(n_881),
.B(n_895),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_923),
.B(n_848),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_925),
.B(n_860),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_909),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_932),
.A2(n_858),
.B(n_895),
.C(n_887),
.Y(n_945)
);

BUFx12f_ASAP7_75t_L g946 ( 
.A(n_910),
.Y(n_946)
);

AO32x2_ASAP7_75t_L g947 ( 
.A1(n_916),
.A2(n_883),
.A3(n_882),
.B1(n_847),
.B2(n_861),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_925),
.B(n_845),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_925),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_932),
.A2(n_858),
.B(n_887),
.C(n_881),
.Y(n_950)
);

OAI21x1_ASAP7_75t_SL g951 ( 
.A1(n_936),
.A2(n_842),
.B(n_869),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_922),
.A2(n_875),
.B(n_868),
.Y(n_952)
);

OA21x2_ASAP7_75t_L g953 ( 
.A1(n_901),
.A2(n_920),
.B(n_926),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_924),
.B(n_845),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_923),
.B(n_856),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_923),
.B(n_856),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_907),
.B(n_859),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_SL g958 ( 
.A1(n_910),
.A2(n_849),
.B1(n_855),
.B2(n_864),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_937),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_932),
.A2(n_898),
.B1(n_868),
.B2(n_865),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_925),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_932),
.A2(n_865),
.B(n_873),
.C(n_843),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_922),
.A2(n_885),
.B(n_871),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_909),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_923),
.B(n_857),
.Y(n_965)
);

NOR2x1_ASAP7_75t_R g966 ( 
.A(n_931),
.B(n_851),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_928),
.A2(n_859),
.B(n_878),
.C(n_863),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_924),
.B(n_883),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_907),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_931),
.B(n_925),
.Y(n_970)
);

CKINVDCx11_ASAP7_75t_R g971 ( 
.A(n_909),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_928),
.A2(n_871),
.B(n_859),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_931),
.B(n_863),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_928),
.A2(n_859),
.B(n_846),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_931),
.A2(n_879),
.B1(n_863),
.B2(n_866),
.Y(n_975)
);

AOI21xp33_ASAP7_75t_SL g976 ( 
.A1(n_924),
.A2(n_33),
.B(n_37),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_907),
.B(n_880),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_907),
.B(n_880),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_927),
.B(n_939),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_931),
.A2(n_876),
.B1(n_854),
.B2(n_844),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_921),
.B(n_876),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_970),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_949),
.B(n_916),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_950),
.A2(n_921),
.B1(n_928),
.B2(n_939),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_943),
.B(n_927),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_970),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_944),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_961),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_949),
.B(n_912),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_955),
.B(n_921),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_964),
.B(n_912),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_979),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_964),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_969),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_955),
.B(n_921),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_959),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_956),
.B(n_914),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_956),
.B(n_914),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_959),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_981),
.B(n_914),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_950),
.A2(n_939),
.B1(n_927),
.B2(n_876),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_948),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_953),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_954),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_965),
.B(n_912),
.Y(n_1005)
);

AND2x4_ASAP7_75t_SL g1006 ( 
.A(n_957),
.B(n_907),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_942),
.B(n_913),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_1007),
.B(n_942),
.Y(n_1008)
);

O2A1O1Ixp5_ASAP7_75t_L g1009 ( 
.A1(n_984),
.A2(n_945),
.B(n_960),
.C(n_941),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_1003),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_990),
.B(n_965),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_988),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1003),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_988),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_1006),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_1003),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_1007),
.B(n_913),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_990),
.B(n_981),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_996),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_995),
.B(n_997),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_996),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_996),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_991),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_992),
.B(n_913),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_982),
.B(n_973),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_994),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_991),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_995),
.B(n_953),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_984),
.A2(n_936),
.B1(n_951),
.B2(n_952),
.Y(n_1029)
);

AND2x2_ASAP7_75t_SL g1030 ( 
.A(n_1029),
.B(n_1006),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1010),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_1024),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1023),
.B(n_987),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1011),
.B(n_1006),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1012),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1023),
.B(n_1004),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_1016),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1012),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1014),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_1024),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_1015),
.B(n_983),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1035),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1031),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1032),
.B(n_1040),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1035),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_1033),
.B(n_1008),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1038),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1038),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1039),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1042),
.Y(n_1050)
);

NOR2xp67_ASAP7_75t_L g1051 ( 
.A(n_1046),
.B(n_1041),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_1046),
.B(n_1034),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_1044),
.B(n_1036),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1045),
.B(n_1034),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1050),
.Y(n_1055)
);

AOI221xp5_ASAP7_75t_L g1056 ( 
.A1(n_1053),
.A2(n_1009),
.B1(n_1048),
.B2(n_1047),
.C(n_1049),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1052),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1051),
.A2(n_1009),
.B(n_1030),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1052),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_1054),
.B(n_946),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_1054),
.B(n_946),
.Y(n_1061)
);

CKINVDCx16_ASAP7_75t_R g1062 ( 
.A(n_1053),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1050),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1052),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_1051),
.A2(n_1030),
.B(n_958),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1052),
.B(n_1030),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_1062),
.B(n_1041),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_1058),
.A2(n_945),
.B(n_962),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1057),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1059),
.Y(n_1070)
);

OAI21xp33_ASAP7_75t_L g1071 ( 
.A1(n_1056),
.A2(n_962),
.B(n_1037),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1055),
.Y(n_1072)
);

OAI21xp33_ASAP7_75t_SL g1073 ( 
.A1(n_1058),
.A2(n_1011),
.B(n_1020),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1063),
.Y(n_1074)
);

AOI32xp33_ASAP7_75t_L g1075 ( 
.A1(n_1066),
.A2(n_1001),
.A3(n_1037),
.B1(n_1028),
.B2(n_1043),
.Y(n_1075)
);

AND2x2_ASAP7_75t_SL g1076 ( 
.A(n_1060),
.B(n_975),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1065),
.A2(n_1043),
.B(n_1001),
.Y(n_1077)
);

OAI21xp33_ASAP7_75t_L g1078 ( 
.A1(n_1064),
.A2(n_1061),
.B(n_1037),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1058),
.A2(n_966),
.B(n_1039),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_1062),
.B(n_1017),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1057),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1064),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1064),
.B(n_1011),
.Y(n_1083)
);

AOI21xp33_ASAP7_75t_L g1084 ( 
.A1(n_1071),
.A2(n_976),
.B(n_37),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1080),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1082),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1068),
.B(n_1028),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1069),
.Y(n_1088)
);

OAI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_1077),
.A2(n_1016),
.B1(n_1037),
.B2(n_1013),
.Y(n_1089)
);

XOR2xp5_ASAP7_75t_L g1090 ( 
.A(n_1067),
.B(n_980),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1070),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1083),
.B(n_1028),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1076),
.B(n_1041),
.Y(n_1093)
);

XNOR2xp5_ASAP7_75t_L g1094 ( 
.A(n_1079),
.B(n_1041),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_1081),
.Y(n_1095)
);

OAI21xp33_ASAP7_75t_SL g1096 ( 
.A1(n_1075),
.A2(n_1020),
.B(n_1018),
.Y(n_1096)
);

AOI32xp33_ASAP7_75t_L g1097 ( 
.A1(n_1071),
.A2(n_1073),
.A3(n_1074),
.B1(n_1072),
.B2(n_1078),
.Y(n_1097)
);

INVxp67_ASAP7_75t_L g1098 ( 
.A(n_1078),
.Y(n_1098)
);

OAI21xp33_ASAP7_75t_L g1099 ( 
.A1(n_1071),
.A2(n_1005),
.B(n_1027),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1080),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1080),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1082),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1084),
.A2(n_1010),
.B(n_1013),
.C(n_1031),
.Y(n_1103)
);

NOR2x1_ASAP7_75t_L g1104 ( 
.A(n_1095),
.B(n_1026),
.Y(n_1104)
);

OAI32xp33_ASAP7_75t_L g1105 ( 
.A1(n_1087),
.A2(n_1008),
.A3(n_1017),
.B1(n_1015),
.B2(n_1025),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1084),
.A2(n_1027),
.B(n_1013),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_SL g1107 ( 
.A(n_1097),
.B(n_936),
.C(n_1026),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1102),
.B(n_1016),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1093),
.B(n_1016),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1085),
.B(n_1020),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1100),
.Y(n_1111)
);

NAND2xp33_ASAP7_75t_L g1112 ( 
.A(n_1101),
.B(n_1016),
.Y(n_1112)
);

XOR2x2_ASAP7_75t_L g1113 ( 
.A(n_1090),
.B(n_972),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1095),
.Y(n_1114)
);

AOI222xp33_ASAP7_75t_L g1115 ( 
.A1(n_1086),
.A2(n_1091),
.B1(n_1088),
.B2(n_1098),
.C1(n_1089),
.C2(n_1096),
.Y(n_1115)
);

AOI211xp5_ASAP7_75t_SL g1116 ( 
.A1(n_1099),
.A2(n_993),
.B(n_1014),
.C(n_969),
.Y(n_1116)
);

NAND4xp75_ASAP7_75t_L g1117 ( 
.A(n_1092),
.B(n_936),
.C(n_974),
.D(n_1010),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1094),
.Y(n_1118)
);

INVxp67_ASAP7_75t_L g1119 ( 
.A(n_1102),
.Y(n_1119)
);

NAND3xp33_ASAP7_75t_L g1120 ( 
.A(n_1119),
.B(n_1016),
.C(n_971),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1110),
.B(n_1016),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1114),
.B(n_1111),
.Y(n_1122)
);

AOI221xp5_ASAP7_75t_L g1123 ( 
.A1(n_1107),
.A2(n_992),
.B1(n_1022),
.B2(n_1021),
.C(n_1019),
.Y(n_1123)
);

NAND3xp33_ASAP7_75t_L g1124 ( 
.A(n_1118),
.B(n_971),
.C(n_993),
.Y(n_1124)
);

AOI221xp5_ASAP7_75t_L g1125 ( 
.A1(n_1103),
.A2(n_1022),
.B1(n_1021),
.B2(n_1019),
.C(n_1002),
.Y(n_1125)
);

INVxp67_ASAP7_75t_SL g1126 ( 
.A(n_1104),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1109),
.A2(n_1015),
.B1(n_1025),
.B2(n_1018),
.Y(n_1127)
);

AOI321xp33_ASAP7_75t_L g1128 ( 
.A1(n_1105),
.A2(n_967),
.A3(n_947),
.B1(n_1019),
.B2(n_1022),
.C(n_1021),
.Y(n_1128)
);

OAI21xp33_ASAP7_75t_L g1129 ( 
.A1(n_1115),
.A2(n_1018),
.B(n_985),
.Y(n_1129)
);

NOR3xp33_ASAP7_75t_L g1130 ( 
.A(n_1108),
.B(n_1112),
.C(n_1117),
.Y(n_1130)
);

NAND4xp75_ASAP7_75t_L g1131 ( 
.A(n_1106),
.B(n_963),
.C(n_998),
.D(n_997),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1115),
.A2(n_967),
.B(n_919),
.C(n_986),
.Y(n_1132)
);

AOI221xp5_ASAP7_75t_L g1133 ( 
.A1(n_1113),
.A2(n_1002),
.B1(n_919),
.B2(n_999),
.C(n_998),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_1116),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1110),
.Y(n_1135)
);

AOI21xp33_ASAP7_75t_L g1136 ( 
.A1(n_1111),
.A2(n_38),
.B(n_39),
.Y(n_1136)
);

AND3x1_ASAP7_75t_L g1137 ( 
.A(n_1114),
.B(n_969),
.C(n_968),
.Y(n_1137)
);

AOI211xp5_ASAP7_75t_L g1138 ( 
.A1(n_1107),
.A2(n_989),
.B(n_983),
.C(n_920),
.Y(n_1138)
);

AOI222xp33_ASAP7_75t_L g1139 ( 
.A1(n_1107),
.A2(n_947),
.B1(n_999),
.B2(n_915),
.C1(n_920),
.C2(n_917),
.Y(n_1139)
);

NAND4xp75_ASAP7_75t_SL g1140 ( 
.A(n_1109),
.B(n_953),
.C(n_1000),
.D(n_968),
.Y(n_1140)
);

AOI221xp5_ASAP7_75t_L g1141 ( 
.A1(n_1107),
.A2(n_919),
.B1(n_983),
.B2(n_989),
.C(n_908),
.Y(n_1141)
);

AO21x1_ASAP7_75t_L g1142 ( 
.A1(n_1114),
.A2(n_39),
.B(n_40),
.Y(n_1142)
);

AOI321xp33_ASAP7_75t_L g1143 ( 
.A1(n_1111),
.A2(n_947),
.A3(n_917),
.B1(n_918),
.B2(n_983),
.C(n_903),
.Y(n_1143)
);

OAI221xp5_ASAP7_75t_L g1144 ( 
.A1(n_1132),
.A2(n_844),
.B1(n_854),
.B2(n_916),
.C(n_907),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_1135),
.Y(n_1145)
);

OAI211xp5_ASAP7_75t_L g1146 ( 
.A1(n_1126),
.A2(n_994),
.B(n_43),
.C(n_44),
.Y(n_1146)
);

NOR3xp33_ASAP7_75t_L g1147 ( 
.A(n_1122),
.B(n_916),
.C(n_44),
.Y(n_1147)
);

AOI211xp5_ASAP7_75t_L g1148 ( 
.A1(n_1134),
.A2(n_41),
.B(n_45),
.C(n_920),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1142),
.Y(n_1149)
);

AO22x2_ASAP7_75t_L g1150 ( 
.A1(n_1124),
.A2(n_947),
.B1(n_45),
.B2(n_41),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_L g1151 ( 
.A(n_1136),
.B(n_911),
.C(n_917),
.Y(n_1151)
);

OAI311xp33_ASAP7_75t_L g1152 ( 
.A1(n_1129),
.A2(n_1123),
.A3(n_1141),
.B1(n_1139),
.C1(n_1133),
.Y(n_1152)
);

OAI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1121),
.A2(n_915),
.B1(n_844),
.B2(n_854),
.Y(n_1153)
);

NOR3xp33_ASAP7_75t_SL g1154 ( 
.A(n_1120),
.B(n_906),
.C(n_903),
.Y(n_1154)
);

OAI211xp5_ASAP7_75t_L g1155 ( 
.A1(n_1130),
.A2(n_908),
.B(n_1000),
.C(n_911),
.Y(n_1155)
);

AOI31xp33_ASAP7_75t_L g1156 ( 
.A1(n_1138),
.A2(n_978),
.A3(n_977),
.B(n_957),
.Y(n_1156)
);

AND3x4_ASAP7_75t_L g1157 ( 
.A(n_1140),
.B(n_978),
.C(n_977),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1131),
.A2(n_978),
.B1(n_977),
.B2(n_919),
.Y(n_1158)
);

AOI322xp5_ASAP7_75t_L g1159 ( 
.A1(n_1128),
.A2(n_918),
.A3(n_917),
.B1(n_915),
.B2(n_914),
.C1(n_905),
.C2(n_957),
.Y(n_1159)
);

NAND4xp25_ASAP7_75t_L g1160 ( 
.A(n_1127),
.B(n_908),
.C(n_911),
.D(n_940),
.Y(n_1160)
);

XNOR2x1_ASAP7_75t_L g1161 ( 
.A(n_1137),
.B(n_918),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1125),
.B(n_914),
.Y(n_1162)
);

OAI211xp5_ASAP7_75t_L g1163 ( 
.A1(n_1143),
.A2(n_908),
.B(n_911),
.C(n_940),
.Y(n_1163)
);

OAI221xp5_ASAP7_75t_SL g1164 ( 
.A1(n_1132),
.A2(n_911),
.B1(n_908),
.B2(n_918),
.C(n_933),
.Y(n_1164)
);

AOI211xp5_ASAP7_75t_L g1165 ( 
.A1(n_1126),
.A2(n_915),
.B(n_911),
.C(n_926),
.Y(n_1165)
);

AOI211xp5_ASAP7_75t_L g1166 ( 
.A1(n_1126),
.A2(n_915),
.B(n_926),
.C(n_935),
.Y(n_1166)
);

NOR2xp67_ASAP7_75t_L g1167 ( 
.A(n_1135),
.B(n_48),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1149),
.A2(n_919),
.B1(n_915),
.B2(n_938),
.Y(n_1168)
);

NAND4xp75_ASAP7_75t_L g1169 ( 
.A(n_1167),
.B(n_905),
.C(n_906),
.D(n_903),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1145),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1150),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1154),
.B(n_938),
.Y(n_1172)
);

OAI21xp33_ASAP7_75t_L g1173 ( 
.A1(n_1147),
.A2(n_940),
.B(n_938),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1146),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1150),
.A2(n_919),
.B1(n_915),
.B2(n_938),
.Y(n_1175)
);

NAND4xp75_ASAP7_75t_L g1176 ( 
.A(n_1158),
.B(n_905),
.C(n_906),
.D(n_52),
.Y(n_1176)
);

NAND4xp75_ASAP7_75t_L g1177 ( 
.A(n_1162),
.B(n_905),
.C(n_51),
.D(n_53),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1148),
.B(n_938),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1161),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1151),
.B(n_938),
.Y(n_1180)
);

NAND4xp75_ASAP7_75t_L g1181 ( 
.A(n_1152),
.B(n_50),
.C(n_63),
.D(n_64),
.Y(n_1181)
);

NOR2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1160),
.B(n_940),
.Y(n_1182)
);

NAND4xp75_ASAP7_75t_L g1183 ( 
.A(n_1159),
.B(n_65),
.C(n_68),
.D(n_70),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_1153),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1155),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1144),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_1156),
.Y(n_1187)
);

NAND4xp75_ASAP7_75t_L g1188 ( 
.A(n_1164),
.B(n_74),
.C(n_75),
.D(n_78),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1165),
.B(n_940),
.Y(n_1189)
);

NOR3xp33_ASAP7_75t_L g1190 ( 
.A(n_1170),
.B(n_1163),
.C(n_1166),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_1171),
.Y(n_1191)
);

NAND2xp33_ASAP7_75t_SL g1192 ( 
.A(n_1174),
.B(n_1157),
.Y(n_1192)
);

NOR2x1p5_ASAP7_75t_L g1193 ( 
.A(n_1181),
.B(n_940),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1179),
.Y(n_1194)
);

NOR2x1_ASAP7_75t_L g1195 ( 
.A(n_1185),
.B(n_935),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1178),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1187),
.A2(n_915),
.B1(n_935),
.B2(n_926),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1184),
.A2(n_935),
.B(n_901),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1175),
.A2(n_915),
.B1(n_935),
.B2(n_933),
.Y(n_1199)
);

AOI322xp5_ASAP7_75t_L g1200 ( 
.A1(n_1186),
.A2(n_915),
.A3(n_929),
.B1(n_934),
.B2(n_935),
.C1(n_937),
.C2(n_930),
.Y(n_1200)
);

OAI322xp33_ASAP7_75t_L g1201 ( 
.A1(n_1175),
.A2(n_934),
.A3(n_929),
.B1(n_937),
.B2(n_930),
.C1(n_904),
.C2(n_902),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1173),
.Y(n_1202)
);

NOR3xp33_ASAP7_75t_L g1203 ( 
.A(n_1177),
.B(n_79),
.C(n_87),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1172),
.B(n_901),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_1192),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1191),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1194),
.Y(n_1207)
);

OAI221xp5_ASAP7_75t_L g1208 ( 
.A1(n_1190),
.A2(n_1168),
.B1(n_1189),
.B2(n_1180),
.C(n_1176),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1202),
.A2(n_1168),
.B1(n_1182),
.B2(n_1183),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1195),
.A2(n_1188),
.B1(n_1169),
.B2(n_935),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1196),
.A2(n_901),
.B(n_933),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1193),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1204),
.A2(n_933),
.B1(n_934),
.B2(n_929),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1203),
.Y(n_1214)
);

NAND3xp33_ASAP7_75t_SL g1215 ( 
.A(n_1198),
.B(n_88),
.C(n_92),
.Y(n_1215)
);

NAND3xp33_ASAP7_75t_SL g1216 ( 
.A(n_1200),
.B(n_94),
.C(n_100),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1199),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1197),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1201),
.A2(n_933),
.B1(n_937),
.B2(n_930),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1205),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1207),
.Y(n_1221)
);

OA22x2_ASAP7_75t_L g1222 ( 
.A1(n_1206),
.A2(n_933),
.B1(n_937),
.B2(n_904),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1208),
.A2(n_933),
.B1(n_930),
.B2(n_904),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1212),
.A2(n_933),
.B1(n_904),
.B2(n_902),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1214),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_1218),
.Y(n_1226)
);

AO22x2_ASAP7_75t_L g1227 ( 
.A1(n_1209),
.A2(n_1216),
.B1(n_1215),
.B2(n_1213),
.Y(n_1227)
);

AO22x2_ASAP7_75t_L g1228 ( 
.A1(n_1217),
.A2(n_904),
.B1(n_902),
.B2(n_106),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1210),
.B(n_933),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1221),
.B(n_1211),
.Y(n_1230)
);

XOR2xp5_ASAP7_75t_L g1231 ( 
.A(n_1220),
.B(n_1219),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1228),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1226),
.Y(n_1233)
);

INVx2_ASAP7_75t_SL g1234 ( 
.A(n_1225),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1223),
.B(n_104),
.C(n_105),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1234),
.A2(n_1231),
.B1(n_1233),
.B2(n_1230),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1232),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1235),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_SL g1239 ( 
.A1(n_1231),
.A2(n_1227),
.B1(n_1224),
.B2(n_1229),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1236),
.A2(n_1222),
.B(n_110),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1240),
.B(n_1237),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1241),
.Y(n_1242)
);

XNOR2xp5_ASAP7_75t_L g1243 ( 
.A(n_1242),
.B(n_1239),
.Y(n_1243)
);

OAI221xp5_ASAP7_75t_R g1244 ( 
.A1(n_1243),
.A2(n_1238),
.B1(n_111),
.B2(n_117),
.C(n_118),
.Y(n_1244)
);

AOI211xp5_ASAP7_75t_L g1245 ( 
.A1(n_1244),
.A2(n_109),
.B(n_119),
.C(n_120),
.Y(n_1245)
);


endmodule