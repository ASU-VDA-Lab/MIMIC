module fake_jpeg_357_n_584 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_584);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_584;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_57),
.B(n_69),
.Y(n_136)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_59),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_60),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_62),
.B(n_63),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_64),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_65),
.B(n_68),
.Y(n_130)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_66),
.Y(n_199)
);

INVx11_ASAP7_75t_SL g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_67),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_1),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_70),
.B(n_88),
.Y(n_147)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_39),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_73),
.B(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_75),
.Y(n_208)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_80),
.Y(n_161)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_81),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_41),
.Y(n_83)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_84),
.Y(n_175)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_1),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_90),
.Y(n_172)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_93),
.Y(n_192)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_94),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_23),
.B(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_2),
.Y(n_166)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_96),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

INVx6_ASAP7_75t_SL g98 ( 
.A(n_20),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_114),
.Y(n_143)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_99),
.Y(n_205)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_100),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_102),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_104),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_107),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

BUFx4f_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

NAND2xp33_ASAP7_75t_SL g111 ( 
.A(n_31),
.B(n_29),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_34),
.Y(n_112)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_112),
.Y(n_215)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_113),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_38),
.B(n_26),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_48),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_123),
.Y(n_144)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_21),
.B(n_2),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_21),
.Y(n_124)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_125),
.A2(n_53),
.B(n_32),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_126),
.Y(n_214)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_54),
.B1(n_56),
.B2(n_26),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g273 ( 
.A1(n_137),
.A2(n_140),
.B1(n_142),
.B2(n_155),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_96),
.A2(n_56),
.B1(n_50),
.B2(n_49),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_76),
.A2(n_56),
.B1(n_50),
.B2(n_49),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_83),
.A2(n_22),
.B1(n_21),
.B2(n_50),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_84),
.A2(n_23),
.B1(n_52),
.B2(n_30),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_158),
.A2(n_180),
.B1(n_201),
.B2(n_219),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_73),
.B(n_36),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_163),
.A2(n_190),
.B(n_194),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_67),
.A2(n_22),
.B1(n_26),
.B2(n_49),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_164),
.A2(n_171),
.B1(n_183),
.B2(n_187),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_166),
.B(n_177),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_116),
.A2(n_22),
.B1(n_29),
.B2(n_35),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_114),
.B(n_123),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_107),
.A2(n_24),
.B1(n_29),
.B2(n_35),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_61),
.A2(n_24),
.B1(n_35),
.B2(n_46),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_100),
.A2(n_40),
.B1(n_52),
.B2(n_46),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_185),
.B(n_207),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_78),
.A2(n_45),
.B1(n_40),
.B2(n_36),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_86),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_189),
.B(n_195),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_75),
.B(n_45),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_64),
.B(n_30),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_59),
.B(n_24),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_197),
.B(n_206),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_109),
.B(n_3),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_12),
.C(n_13),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_87),
.A2(n_53),
.B1(n_6),
.B2(n_7),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_97),
.B(n_3),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_202),
.B(n_211),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_120),
.A2(n_53),
.B1(n_7),
.B2(n_8),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_203),
.A2(n_209),
.B1(n_216),
.B2(n_217),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_64),
.B(n_17),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_60),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_101),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_102),
.B(n_8),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_91),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_94),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_105),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_106),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_148),
.B(n_66),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_220),
.Y(n_318)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_134),
.Y(n_221)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_221),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_222),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_132),
.Y(n_223)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_223),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_147),
.B(n_126),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_224),
.B(n_230),
.Y(n_304)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_139),
.Y(n_226)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_226),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_148),
.A2(n_81),
.B(n_80),
.C(n_103),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g339 ( 
.A1(n_227),
.A2(n_236),
.B(n_228),
.C(n_285),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_163),
.B(n_93),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_228),
.B(n_240),
.Y(n_335)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_229),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_122),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_232),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_130),
.B(n_93),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_233),
.B(n_238),
.Y(n_329)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_234),
.Y(n_328)
);

A2O1A1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_136),
.A2(n_103),
.B(n_72),
.C(n_108),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_150),
.B(n_72),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_239),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_161),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_242),
.Y(n_332)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_135),
.Y(n_244)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_244),
.Y(n_346)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_133),
.Y(n_246)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_246),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_128),
.B(n_82),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_247),
.B(n_249),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_161),
.Y(n_248)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_248),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_143),
.B(n_79),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_117),
.B1(n_115),
.B2(n_99),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_250),
.A2(n_266),
.B1(n_268),
.B2(n_277),
.Y(n_343)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_251),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_149),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_252),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_144),
.B(n_154),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_253),
.B(n_258),
.Y(n_308)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_175),
.Y(n_254)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_254),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_190),
.A2(n_108),
.B1(n_15),
.B2(n_16),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_255),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_199),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_256),
.B(n_264),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_182),
.B(n_14),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_257),
.B(n_259),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_198),
.B(n_14),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_178),
.B(n_15),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_184),
.A2(n_16),
.B1(n_17),
.B2(n_167),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_260),
.B(n_262),
.Y(n_338)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_138),
.Y(n_261)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_261),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_151),
.B(n_17),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_152),
.B(n_162),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_146),
.C(n_160),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_219),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_133),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_271),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_135),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_267),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_183),
.A2(n_137),
.B1(n_203),
.B2(n_142),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_159),
.A2(n_167),
.B1(n_156),
.B2(n_210),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_269),
.A2(n_260),
.B1(n_241),
.B2(n_264),
.Y(n_324)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_213),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_270),
.Y(n_353)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_172),
.Y(n_271)
);

AO22x1_ASAP7_75t_SL g272 ( 
.A1(n_200),
.A2(n_156),
.B1(n_153),
.B2(n_146),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_272),
.B(n_286),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_149),
.B(n_208),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_274),
.B(n_275),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_131),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_173),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_279),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_155),
.A2(n_140),
.B1(n_171),
.B2(n_164),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_153),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_278),
.B(n_280),
.Y(n_310)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_141),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_169),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_173),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_281),
.B(n_284),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_169),
.A2(n_214),
.B1(n_188),
.B2(n_186),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_282),
.A2(n_222),
.B1(n_223),
.B2(n_267),
.Y(n_352)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_159),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_283),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_208),
.B(n_196),
.Y(n_284)
);

NAND2xp33_ASAP7_75t_SL g285 ( 
.A(n_131),
.B(n_129),
.Y(n_285)
);

NOR2x1_ASAP7_75t_R g340 ( 
.A(n_285),
.B(n_248),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_157),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_179),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_287),
.B(n_288),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_192),
.Y(n_288)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_145),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_145),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_181),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_170),
.A2(n_174),
.B1(n_205),
.B2(n_168),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_293),
.A2(n_269),
.B1(n_248),
.B2(n_291),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_181),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_294),
.B(n_297),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_179),
.B(n_214),
.Y(n_297)
);

AOI32xp33_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_205),
.A3(n_170),
.B1(n_186),
.B2(n_188),
.Y(n_299)
);

AOI32xp33_ASAP7_75t_L g383 ( 
.A1(n_299),
.A2(n_342),
.A3(n_312),
.B1(n_309),
.B2(n_322),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_300),
.B(n_339),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_220),
.B(n_204),
.C(n_168),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_307),
.B(n_299),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_224),
.B(n_174),
.CI(n_160),
.CON(n_309),
.SN(n_309)
);

MAJx2_ASAP7_75t_L g380 ( 
.A(n_309),
.B(n_279),
.C(n_289),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_235),
.A2(n_176),
.B1(n_204),
.B2(n_239),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_314),
.A2(n_345),
.B1(n_352),
.B2(n_270),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_225),
.A2(n_176),
.B1(n_266),
.B2(n_296),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_316),
.A2(n_321),
.B1(n_322),
.B2(n_325),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_296),
.A2(n_230),
.B1(n_236),
.B2(n_295),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_282),
.A2(n_245),
.B1(n_262),
.B2(n_227),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_324),
.A2(n_347),
.B1(n_283),
.B2(n_275),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_221),
.A2(n_226),
.B1(n_272),
.B2(n_287),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_272),
.A2(n_286),
.B1(n_258),
.B2(n_254),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_326),
.Y(n_357)
);

BUFx5_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_262),
.A2(n_228),
.B1(n_273),
.B2(n_263),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_308),
.B(n_237),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_354),
.B(n_364),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_243),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_361),
.Y(n_406)
);

NAND2x1p5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_220),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_358),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_359),
.Y(n_397)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_315),
.Y(n_360)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_351),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_263),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_362),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_273),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_363),
.B(n_367),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_308),
.B(n_253),
.Y(n_364)
);

OAI22xp33_ASAP7_75t_L g404 ( 
.A1(n_365),
.A2(n_373),
.B1(n_298),
.B2(n_352),
.Y(n_404)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_311),
.Y(n_366)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_366),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_309),
.B(n_273),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_311),
.Y(n_368)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_315),
.Y(n_369)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_369),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_343),
.A2(n_273),
.B1(n_280),
.B2(n_271),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_370),
.A2(n_371),
.B1(n_382),
.B2(n_365),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_314),
.A2(n_261),
.B1(n_229),
.B2(n_234),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_339),
.A2(n_242),
.B(n_251),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_372),
.A2(n_383),
.B(n_342),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_303),
.B(n_246),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_374),
.B(n_376),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_318),
.B(n_265),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_375),
.B(n_388),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_278),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_317),
.Y(n_377)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_377),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_321),
.B(n_276),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_378),
.B(n_380),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_332),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_379),
.B(n_384),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_316),
.A2(n_232),
.B1(n_244),
.B2(n_312),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_301),
.B(n_329),
.Y(n_384)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_385),
.B(n_386),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_303),
.B(n_338),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_338),
.B(n_344),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_387),
.B(n_390),
.Y(n_423)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_338),
.B(n_344),
.Y(n_391)
);

XOR2x2_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_396),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_323),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_392),
.Y(n_402)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_333),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_329),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_394),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_331),
.B(n_302),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_395),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_307),
.B(n_300),
.Y(n_396)
);

OAI21xp33_ASAP7_75t_SL g444 ( 
.A1(n_398),
.A2(n_362),
.B(n_381),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_396),
.B(n_319),
.C(n_330),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_403),
.B(n_375),
.C(n_358),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_404),
.A2(n_409),
.B1(n_412),
.B2(n_414),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_363),
.A2(n_320),
.B1(n_334),
.B2(n_335),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_370),
.A2(n_320),
.B1(n_334),
.B2(n_335),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_413),
.A2(n_368),
.B1(n_371),
.B2(n_385),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_367),
.A2(n_382),
.B1(n_355),
.B2(n_361),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_372),
.A2(n_335),
.B(n_353),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_420),
.A2(n_389),
.B(n_388),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_421),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_379),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_422),
.B(n_426),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_355),
.A2(n_310),
.B1(n_353),
.B2(n_346),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_355),
.A2(n_346),
.B1(n_341),
.B2(n_305),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_427),
.A2(n_369),
.B1(n_360),
.B2(n_359),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_356),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_391),
.Y(n_436)
);

AND2x4_ASAP7_75t_SL g431 ( 
.A(n_381),
.B(n_330),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_431),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g432 ( 
.A1(n_389),
.A2(n_349),
.B(n_337),
.Y(n_432)
);

O2A1O1Ixp33_ASAP7_75t_L g434 ( 
.A1(n_432),
.A2(n_357),
.B(n_393),
.C(n_387),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_429),
.A2(n_373),
.B1(n_357),
.B2(n_362),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_433),
.A2(n_458),
.B1(n_412),
.B2(n_409),
.Y(n_479)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_434),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_390),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_435),
.B(n_438),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_437),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_421),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_386),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_403),
.B(n_378),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_439),
.B(n_416),
.Y(n_489)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_407),
.Y(n_440)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_440),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_441),
.B(n_428),
.Y(n_476)
);

XNOR2x1_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_380),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_443),
.B(n_444),
.Y(n_472)
);

OA21x2_ASAP7_75t_SL g445 ( 
.A1(n_405),
.A2(n_375),
.B(n_358),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_445),
.B(n_405),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_456),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_408),
.B(n_377),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_448),
.B(n_452),
.C(n_460),
.Y(n_475)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_407),
.Y(n_449)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_449),
.Y(n_486)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_411),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_453),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_408),
.B(n_366),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_420),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_454),
.A2(n_455),
.B1(n_461),
.B2(n_463),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_427),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_411),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_457),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_406),
.A2(n_341),
.B1(n_350),
.B2(n_349),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_400),
.B(n_337),
.C(n_350),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_424),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_421),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_462),
.Y(n_473)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_424),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_398),
.A2(n_306),
.B(n_336),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_464),
.A2(n_430),
.B(n_422),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_446),
.A2(n_406),
.B1(n_414),
.B2(n_418),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_467),
.A2(n_471),
.B1(n_491),
.B2(n_442),
.Y(n_496)
);

AO21x1_ASAP7_75t_L g499 ( 
.A1(n_468),
.A2(n_478),
.B(n_453),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_446),
.A2(n_418),
.B1(n_400),
.B2(n_399),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_476),
.B(n_480),
.C(n_484),
.Y(n_497)
);

FAx1_ASAP7_75t_SL g478 ( 
.A(n_443),
.B(n_399),
.CI(n_428),
.CON(n_478),
.SN(n_478)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_479),
.A2(n_481),
.B1(n_493),
.B2(n_442),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_435),
.B(n_428),
.C(n_430),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_456),
.A2(n_413),
.B1(n_432),
.B2(n_426),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_458),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_483),
.B(n_463),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_438),
.B(n_416),
.C(n_425),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_439),
.B(n_431),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_490),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_441),
.B(n_416),
.C(n_425),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_488),
.C(n_451),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_448),
.B(n_416),
.C(n_432),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_489),
.B(n_451),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_452),
.B(n_431),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_447),
.A2(n_432),
.B1(n_410),
.B2(n_402),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_464),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_494),
.B(n_501),
.Y(n_532)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_469),
.Y(n_495)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_495),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_496),
.A2(n_498),
.B1(n_511),
.B2(n_512),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_499),
.A2(n_514),
.B(n_490),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_474),
.B(n_460),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_466),
.Y(n_502)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_502),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_503),
.B(n_505),
.C(n_510),
.Y(n_525)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_477),
.Y(n_504)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_504),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_491),
.B(n_465),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_506),
.B(n_485),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_481),
.A2(n_459),
.B1(n_434),
.B2(n_410),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_507),
.A2(n_514),
.B1(n_504),
.B2(n_502),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_470),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_509),
.Y(n_520)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_486),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_433),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_492),
.A2(n_419),
.B1(n_479),
.B2(n_417),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_482),
.A2(n_419),
.B1(n_417),
.B2(n_402),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_475),
.B(n_487),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_513),
.B(n_476),
.C(n_480),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_482),
.A2(n_459),
.B(n_431),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_515),
.A2(n_516),
.B1(n_440),
.B2(n_421),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_482),
.A2(n_461),
.B1(n_457),
.B2(n_450),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_506),
.A2(n_488),
.B(n_471),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_518),
.B(n_522),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_496),
.A2(n_467),
.B1(n_473),
.B2(n_478),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_516),
.Y(n_523)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_523),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_524),
.B(n_529),
.Y(n_544)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_526),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_533),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_472),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_499),
.A2(n_484),
.B(n_489),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_507),
.B(n_449),
.Y(n_530)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_530),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_532),
.B(n_513),
.C(n_503),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_535),
.B(n_536),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_532),
.B(n_497),
.C(n_501),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g538 ( 
.A(n_520),
.B(n_497),
.Y(n_538)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_538),
.Y(n_550)
);

OAI221xp5_ASAP7_75t_L g539 ( 
.A1(n_529),
.A2(n_510),
.B1(n_494),
.B2(n_505),
.C(n_478),
.Y(n_539)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_539),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_500),
.C(n_472),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_541),
.B(n_542),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_521),
.A2(n_500),
.B(n_415),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_545),
.A2(n_548),
.B(n_530),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_518),
.B(n_522),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_547),
.B(n_527),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_517),
.B(n_523),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_535),
.B(n_525),
.C(n_524),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_549),
.B(n_555),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_551),
.Y(n_569)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_552),
.Y(n_562)
);

AO21x1_ASAP7_75t_L g554 ( 
.A1(n_534),
.A2(n_526),
.B(n_519),
.Y(n_554)
);

AO21x1_ASAP7_75t_L g568 ( 
.A1(n_554),
.A2(n_543),
.B(n_541),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_546),
.A2(n_519),
.B1(n_517),
.B2(n_531),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_536),
.B(n_525),
.C(n_415),
.Y(n_556)
);

NOR2xp67_ASAP7_75t_L g563 ( 
.A(n_556),
.B(n_559),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_537),
.A2(n_531),
.B(n_401),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_557),
.A2(n_543),
.B(n_397),
.Y(n_566)
);

AOI21x1_ASAP7_75t_L g559 ( 
.A1(n_540),
.A2(n_401),
.B(n_397),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_553),
.A2(n_545),
.B(n_544),
.Y(n_561)
);

AOI21xp33_ASAP7_75t_L g574 ( 
.A1(n_561),
.A2(n_306),
.B(n_336),
.Y(n_574)
);

FAx1_ASAP7_75t_SL g564 ( 
.A(n_549),
.B(n_544),
.CI(n_547),
.CON(n_564),
.SN(n_564)
);

A2O1A1Ixp33_ASAP7_75t_SL g570 ( 
.A1(n_564),
.A2(n_556),
.B(n_550),
.C(n_551),
.Y(n_570)
);

INVx11_ASAP7_75t_L g565 ( 
.A(n_554),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_565),
.A2(n_566),
.B1(n_557),
.B2(n_555),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_568),
.B(n_327),
.Y(n_573)
);

AOI221xp5_ASAP7_75t_L g577 ( 
.A1(n_570),
.A2(n_571),
.B1(n_573),
.B2(n_574),
.C(n_575),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_567),
.B(n_558),
.C(n_560),
.Y(n_571)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_572),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_562),
.B(n_327),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_570),
.B(n_565),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_578),
.B(n_569),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_576),
.A2(n_563),
.B(n_568),
.Y(n_579)
);

OAI21xp33_ASAP7_75t_L g581 ( 
.A1(n_579),
.A2(n_580),
.B(n_569),
.Y(n_581)
);

AOI21x1_ASAP7_75t_L g582 ( 
.A1(n_581),
.A2(n_577),
.B(n_566),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_582),
.A2(n_328),
.B1(n_564),
.B2(n_577),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_583),
.B(n_564),
.Y(n_584)
);


endmodule