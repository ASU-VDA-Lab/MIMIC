module fake_jpeg_20927_n_322 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_32),
.B1(n_21),
.B2(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_60),
.B1(n_68),
.B2(n_24),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_62),
.Y(n_97)
);

CKINVDCx9p33_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_55),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_78),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_36),
.B1(n_32),
.B2(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_27),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_65),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_32),
.B1(n_19),
.B2(n_33),
.Y(n_68)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_71),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_75),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_18),
.B1(n_23),
.B2(n_33),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_79),
.B1(n_26),
.B2(n_23),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_77),
.B(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_19),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_18),
.B1(n_23),
.B2(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_38),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_90),
.B(n_96),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_59),
.A2(n_78),
.B(n_81),
.Y(n_91)
);

OAI21x1_ASAP7_75t_SL g153 ( 
.A1(n_91),
.A2(n_103),
.B(n_3),
.Y(n_153)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_26),
.B1(n_18),
.B2(n_28),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_106),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_28),
.B1(n_26),
.B2(n_70),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_102),
.Y(n_140)
);

NAND2xp33_ASAP7_75t_R g103 ( 
.A(n_55),
.B(n_36),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_108),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_28),
.B1(n_30),
.B2(n_35),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_116),
.B1(n_63),
.B2(n_72),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_30),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_54),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_113),
.B1(n_63),
.B2(n_2),
.Y(n_144)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_57),
.A2(n_22),
.B1(n_36),
.B2(n_37),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_54),
.B(n_61),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_119),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_60),
.B(n_31),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_72),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_37),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_67),
.B(n_31),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_121),
.A2(n_127),
.B(n_146),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_80),
.B1(n_69),
.B2(n_63),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_118),
.B1(n_113),
.B2(n_112),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_98),
.A2(n_31),
.B(n_80),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_72),
.A3(n_37),
.B1(n_17),
.B2(n_31),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_31),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_130),
.B(n_139),
.Y(n_163)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_17),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_63),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_141),
.B(n_145),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_90),
.B1(n_85),
.B2(n_119),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_72),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_1),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_148),
.B(n_150),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_1),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_85),
.B(n_2),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_117),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_101),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_3),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_6),
.Y(n_172)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_167),
.B1(n_149),
.B2(n_155),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_159),
.A2(n_129),
.B1(n_143),
.B2(n_137),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_160),
.A2(n_188),
.B(n_136),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_177),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_5),
.C(n_6),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_162),
.B(n_168),
.Y(n_203)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_176),
.Y(n_195)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_125),
.A2(n_111),
.B1(n_115),
.B2(n_84),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_131),
.B(n_5),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_170),
.B(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_172),
.B(n_178),
.Y(n_216)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_110),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_94),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_128),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_108),
.C(n_104),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_183),
.C(n_121),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_120),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_182),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_94),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_134),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_185),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_152),
.B(n_84),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_140),
.A2(n_92),
.B1(n_99),
.B2(n_110),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_125),
.A2(n_155),
.B(n_140),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_170),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_193),
.A2(n_211),
.B1(n_187),
.B2(n_184),
.Y(n_228)
);

OAI21x1_ASAP7_75t_R g198 ( 
.A1(n_179),
.A2(n_137),
.B(n_127),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_199),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_169),
.Y(n_199)
);

NAND2x1p5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_128),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_205),
.A2(n_202),
.B(n_196),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_156),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_207),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_166),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_142),
.Y(n_208)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_157),
.A2(n_153),
.B(n_144),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_157),
.B1(n_175),
.B2(n_164),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_138),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_215),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_160),
.B1(n_158),
.B2(n_167),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_161),
.B(n_143),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_151),
.C(n_123),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_181),
.C(n_188),
.Y(n_224)
);

INVx5_ASAP7_75t_SL g218 ( 
.A(n_180),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_133),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_222),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_217),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_220),
.B(n_223),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_228),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_160),
.B1(n_159),
.B2(n_173),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_189),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_225),
.C(n_231),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_205),
.B(n_163),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_168),
.B1(n_165),
.B2(n_132),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_232),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_215),
.B1(n_193),
.B2(n_213),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_190),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_238),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_186),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_236),
.C(n_200),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_192),
.B(n_87),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_176),
.B1(n_174),
.B2(n_151),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_192),
.B(n_87),
.C(n_123),
.Y(n_240)
);

OAI322xp33_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_206),
.A3(n_199),
.B1(n_207),
.B2(n_196),
.C1(n_212),
.C2(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_242),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_246),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_239),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_259),
.Y(n_265)
);

BUFx4f_ASAP7_75t_SL g253 ( 
.A(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_198),
.C(n_194),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_256),
.C(n_236),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_198),
.C(n_194),
.Y(n_256)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_260),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_234),
.B(n_216),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_253),
.C(n_8),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_257),
.Y(n_263)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_248),
.A2(n_223),
.B(n_225),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_264),
.A2(n_278),
.B1(n_252),
.B2(n_247),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_231),
.C(n_222),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_272),
.C(n_275),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_248),
.A2(n_235),
.B1(n_232),
.B2(n_242),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_258),
.B1(n_218),
.B2(n_210),
.Y(n_287)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_277),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_212),
.B1(n_203),
.B2(n_230),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_240),
.C(n_190),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_201),
.Y(n_273)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_209),
.C(n_197),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_261),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_244),
.A2(n_197),
.B(n_218),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_249),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_283),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_278),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_287),
.B1(n_265),
.B2(n_264),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_286),
.A2(n_268),
.B(n_270),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_174),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_291),
.Y(n_300)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_296),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_294),
.A2(n_295),
.B1(n_281),
.B2(n_289),
.Y(n_303)
);

NAND3xp33_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_269),
.C(n_265),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_290),
.A2(n_275),
.B(n_267),
.Y(n_296)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_272),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_280),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_7),
.C(n_8),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_284),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_303),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_307),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_279),
.A3(n_291),
.B1(n_285),
.B2(n_297),
.C1(n_253),
.C2(n_12),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_299),
.Y(n_307)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_306),
.A2(n_285),
.B(n_8),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_313),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_308),
.B1(n_305),
.B2(n_301),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_315),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_312),
.B(n_314),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_9),
.Y(n_319)
);

AOI211xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_318),
.B(n_10),
.C(n_11),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_320),
.B(n_9),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_9),
.Y(n_322)
);


endmodule