module fake_jpeg_28550_n_181 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_181);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx2_ASAP7_75t_R g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_7),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_78),
.Y(n_86)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_77),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_66),
.Y(n_78)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_80),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_0),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_60),
.B1(n_70),
.B2(n_68),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_88),
.B1(n_89),
.B2(n_93),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_71),
.B1(n_64),
.B2(n_65),
.Y(n_88)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_65),
.B1(n_71),
.B2(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_56),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_61),
.B1(n_51),
.B2(n_52),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_60),
.B1(n_68),
.B2(n_70),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_58),
.B1(n_53),
.B2(n_77),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_91),
.B(n_87),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_3),
.B(n_4),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_77),
.B1(n_60),
.B2(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_104),
.B1(n_4),
.B2(n_5),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_75),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_105),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_110),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_50),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_24),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_69),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_67),
.B1(n_55),
.B2(n_79),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_129),
.B1(n_131),
.B2(n_116),
.Y(n_138)
);

AO22x1_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_63),
.B1(n_18),
.B2(n_19),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_0),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_95),
.B(n_63),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_5),
.C(n_6),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_1),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_1),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_2),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_128),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_2),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_129),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_3),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_27),
.B1(n_47),
.B2(n_46),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_124),
.B(n_127),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_135),
.Y(n_164)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_137),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_138),
.A2(n_148),
.B1(n_150),
.B2(n_13),
.Y(n_163)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_143),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

NOR2x1p5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_29),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_144),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_149),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_48),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_116),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_152),
.C(n_12),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_34),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_42),
.A3(n_32),
.B1(n_35),
.B2(n_15),
.C1(n_17),
.C2(n_41),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_140),
.C(n_153),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_161),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_164),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_147),
.B1(n_158),
.B2(n_157),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_169),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_172),
.B1(n_171),
.B2(n_165),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_171),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_160),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_156),
.C(n_149),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_178),
.A2(n_154),
.B1(n_152),
.B2(n_155),
.Y(n_179)
);

AO21x1_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_146),
.B(n_162),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_162),
.Y(n_181)
);


endmodule