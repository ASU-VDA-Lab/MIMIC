module real_jpeg_29830_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_336, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_336;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_286;
wire n_166;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_0),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_SL g108 ( 
.A1(n_0),
.A2(n_29),
.B(n_33),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_0),
.B(n_31),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_0),
.A2(n_55),
.B(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_0),
.B(n_55),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_0),
.B(n_68),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_0),
.A2(n_130),
.B1(n_132),
.B2(n_198),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_0),
.A2(n_32),
.B(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_1),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_1),
.A2(n_45),
.B1(n_55),
.B2(n_56),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_45),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_90),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_2),
.A2(n_50),
.B1(n_52),
.B2(n_90),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_90),
.Y(n_218)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_3),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_5),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_95),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_5),
.A2(n_50),
.B1(n_52),
.B2(n_95),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_95),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_36),
.B1(n_55),
.B2(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_7),
.A2(n_36),
.B1(n_50),
.B2(n_52),
.Y(n_151)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_9),
.A2(n_55),
.B1(n_56),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_9),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_9),
.A2(n_50),
.B1(n_52),
.B2(n_98),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_98),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_98),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_10),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_10),
.A2(n_27),
.B1(n_50),
.B2(n_52),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_10),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_88),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_11),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_88),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_88),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_11),
.A2(n_50),
.B1(n_52),
.B2(n_88),
.Y(n_191)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_13),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_105),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_105),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_13),
.A2(n_50),
.B1(n_52),
.B2(n_105),
.Y(n_198)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_15),
.A2(n_55),
.B1(n_56),
.B2(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_16),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_17),
.A2(n_43),
.B1(n_50),
.B2(n_52),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_17),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_255)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_328),
.B(n_331),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_76),
.B(n_327),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_21),
.B(n_37),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_21),
.B(n_329),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_21),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_23),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_25),
.A2(n_34),
.B(n_102),
.C(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_31),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_28),
.A2(n_31),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_28),
.A2(n_31),
.B1(n_139),
.B2(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_28),
.A2(n_31),
.B1(n_158),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_28),
.A2(n_31),
.B(n_35),
.Y(n_330)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_31),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_32),
.A2(n_62),
.B(n_64),
.C(n_65),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_62),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_32),
.A2(n_56),
.A3(n_62),
.B1(n_215),
.B2(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_33),
.B(n_102),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_69),
.C(n_71),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_38),
.A2(n_39),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_58),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_40),
.B(n_312),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_42),
.A2(n_73),
.B1(n_75),
.B2(n_280),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_46),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_46),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_46),
.A2(n_58),
.B1(n_306),
.B2(n_313),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_53),
.B(n_57),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_47),
.A2(n_53),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_47),
.A2(n_53),
.B1(n_128),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_47),
.A2(n_53),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_47),
.A2(n_53),
.B1(n_172),
.B2(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_47),
.B(n_102),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_47),
.A2(n_53),
.B1(n_94),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_47),
.A2(n_53),
.B1(n_57),
.B2(n_262),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_48),
.A2(n_52),
.A3(n_55),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_49),
.B(n_50),
.Y(n_176)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_50),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_50),
.B(n_204),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_55),
.B(n_66),
.Y(n_223)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_58),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_59),
.A2(n_60),
.B1(n_68),
.B2(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_60),
.A2(n_68),
.B1(n_87),
.B2(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_60),
.A2(n_68),
.B1(n_142),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_60),
.A2(n_68),
.B1(n_160),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_65),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_65),
.B1(n_86),
.B2(n_89),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_61),
.A2(n_65),
.B1(n_89),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_61),
.A2(n_65),
.B1(n_119),
.B2(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_61),
.A2(n_65),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_325),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_69),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_73),
.A2(n_75),
.B1(n_104),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_73),
.A2(n_75),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_320),
.B(n_326),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_297),
.A3(n_316),
.B1(n_318),
.B2(n_319),
.C(n_336),
.Y(n_77)
);

AOI321xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_249),
.A3(n_286),
.B1(n_291),
.B2(n_296),
.C(n_337),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_144),
.C(n_162),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_123),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_81),
.B(n_123),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_106),
.C(n_115),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_82),
.B(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_100),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_91),
.B2(n_92),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_92),
.C(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_96),
.A2(n_99),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_96),
.A2(n_99),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_97),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_102),
.B(n_132),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_106),
.A2(n_115),
.B1(n_116),
.B2(n_247),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_106),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_109),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_110),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx5_ASAP7_75t_SL g199 ( 
.A(n_111),
.Y(n_199)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_122),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_117),
.B(n_234),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_120),
.B(n_122),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_121),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_135),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_134),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_134),
.C(n_135),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_129),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_132),
.B1(n_133),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_130),
.A2(n_132),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_130),
.A2(n_191),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_130),
.A2(n_132),
.B1(n_186),
.B2(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_130),
.A2(n_132),
.B(n_151),
.Y(n_264)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_143),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_140),
.C(n_143),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g292 ( 
.A1(n_145),
.A2(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_146),
.B(n_147),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_161),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_149),
.B(n_154),
.C(n_161),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_150),
.B(n_152),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_153),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_155),
.B(n_157),
.C(n_159),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_243),
.B(n_248),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_229),
.B(n_242),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_208),
.B(n_228),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_187),
.B(n_207),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_177),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_167),
.B(n_177),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_173),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_171),
.Y(n_175)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_182),
.C(n_184),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_183),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_195),
.B(n_206),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_189),
.B(n_194),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_201),
.B(n_205),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_197),
.B(n_200),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_209),
.B(n_210),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_221),
.B1(n_226),
.B2(n_227),
.Y(n_210)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_212),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_220),
.C(n_227),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_218),
.Y(n_239)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_224),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_230),
.B(n_231),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_238),
.C(n_240),
.Y(n_244)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_266),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_266),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_257),
.C(n_265),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_257),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_251),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_254),
.CI(n_256),
.CON(n_251),
.SN(n_251)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_254),
.C(n_256),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_253),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_255),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_263),
.B2(n_264),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_258),
.B(n_264),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_264),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_263),
.A2(n_278),
.B(n_281),
.Y(n_308)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_284),
.B2(n_285),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_275),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_269),
.B(n_275),
.C(n_285),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_273),
.B(n_274),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_273),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_272),
.Y(n_304)
);

FAx1_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_299),
.CI(n_308),
.CON(n_298),
.SN(n_298)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_275)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_276),
.Y(n_283)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_284),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_287),
.A2(n_292),
.B(n_295),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_289),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_309),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_298),
.B(n_317),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_309),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_302),
.B2(n_307),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_301),
.B1(n_311),
.B2(n_314),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_303),
.C(n_306),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_314),
.C(n_315),
.Y(n_321)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_302),
.Y(n_307)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_315),
.Y(n_309)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_311),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_330),
.B(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_332),
.Y(n_331)
);


endmodule