module fake_jpeg_13690_n_480 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_480);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_480;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_47),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_7),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_48),
.B(n_69),
.Y(n_124)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_53),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_57),
.Y(n_141)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_83),
.Y(n_100)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_7),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_35),
.B(n_7),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_93),
.Y(n_127)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_92),
.Y(n_101)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_21),
.B1(n_28),
.B2(n_26),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_94),
.A2(n_45),
.B1(n_66),
.B2(n_137),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_48),
.B(n_35),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_118),
.B(n_122),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_SL g120 ( 
.A(n_69),
.B(n_39),
.C(n_24),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_52),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_37),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_57),
.A2(n_18),
.B1(n_41),
.B2(n_32),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_138),
.B1(n_146),
.B2(n_42),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_68),
.B(n_37),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_47),
.B(n_39),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_65),
.A2(n_18),
.B1(n_41),
.B2(n_32),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_61),
.A2(n_21),
.B1(n_39),
.B2(n_24),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_143),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_149),
.Y(n_204)
);

AOI32xp33_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_26),
.A3(n_28),
.B1(n_53),
.B2(n_76),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_150),
.A2(n_191),
.B(n_192),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_37),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_171),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_95),
.C(n_99),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_185),
.C(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_156),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_101),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_158),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_37),
.Y(n_158)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

BUFx2_ASAP7_75t_SL g219 ( 
.A(n_159),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_160),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_100),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_161),
.B(n_178),
.Y(n_228)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_137),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_168),
.B(n_179),
.Y(n_227)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_120),
.A2(n_93),
.B1(n_91),
.B2(n_89),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_170),
.A2(n_175),
.B1(n_94),
.B2(n_59),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_116),
.A2(n_17),
.B(n_41),
.C(n_32),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_24),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_183),
.Y(n_211)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_107),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_175)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_125),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_97),
.B(n_26),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_111),
.B(n_26),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_186),
.Y(n_206)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_182),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_42),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_184),
.A2(n_187),
.B1(n_189),
.B2(n_147),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_98),
.B(n_28),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_128),
.B(n_42),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_188),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_144),
.B(n_19),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_108),
.B(n_19),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_128),
.B(n_19),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_148),
.B1(n_185),
.B2(n_142),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_178),
.A2(n_113),
.B1(n_129),
.B2(n_104),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_157),
.A2(n_113),
.B1(n_142),
.B2(n_147),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_152),
.A2(n_135),
.B1(n_21),
.B2(n_140),
.Y(n_213)
);

OAI211xp5_ASAP7_75t_L g238 ( 
.A1(n_213),
.A2(n_192),
.B(n_186),
.C(n_155),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_160),
.A2(n_80),
.B1(n_70),
.B2(n_67),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_183),
.B1(n_139),
.B2(n_176),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_230),
.A2(n_231),
.B1(n_237),
.B2(n_250),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_171),
.B(n_154),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_232),
.A2(n_233),
.B(n_159),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_205),
.A2(n_173),
.B1(n_149),
.B2(n_177),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_203),
.A2(n_228),
.B(n_221),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_235),
.A2(n_258),
.B(n_216),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_249),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_104),
.B1(n_139),
.B2(n_112),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_238),
.B(n_242),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_153),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_251),
.C(n_252),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_210),
.A2(n_175),
.B1(n_181),
.B2(n_182),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_240),
.A2(n_201),
.B1(n_166),
.B2(n_194),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_215),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_204),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_193),
.Y(n_242)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

NOR2x1p5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_185),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_247),
.B(n_217),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_161),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_172),
.B1(n_165),
.B2(n_162),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_163),
.C(n_156),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_123),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_174),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_255),
.Y(n_276)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_221),
.B(n_164),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_103),
.B1(n_112),
.B2(n_115),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_237),
.B1(n_231),
.B2(n_233),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_209),
.A2(n_213),
.B(n_227),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_249),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_259),
.B(n_272),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_232),
.A2(n_209),
.B(n_200),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_265),
.A2(n_283),
.B(n_284),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_253),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_274),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_268),
.A2(n_287),
.B1(n_246),
.B2(n_245),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_220),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_270),
.B(n_247),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_204),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_241),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_230),
.A2(n_220),
.B1(n_217),
.B2(n_130),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_275),
.A2(n_219),
.B1(n_194),
.B2(n_197),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_229),
.A2(n_201),
.B1(n_187),
.B2(n_189),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_277),
.A2(n_219),
.B1(n_202),
.B2(n_223),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_239),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_197),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_258),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_282),
.B(n_286),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_235),
.A2(n_216),
.B(n_214),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_236),
.B(n_214),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_248),
.A2(n_198),
.B(n_215),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_240),
.A2(n_202),
.B1(n_198),
.B2(n_130),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_288),
.A2(n_257),
.B1(n_250),
.B2(n_243),
.Y(n_301)
);

OAI32xp33_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_255),
.A3(n_247),
.B1(n_238),
.B2(n_254),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_293),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_234),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_252),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_297),
.C(n_300),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_264),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_299),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_284),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_251),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_260),
.Y(n_298)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_251),
.C(n_239),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_301),
.A2(n_309),
.B1(n_312),
.B2(n_195),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_303),
.A2(n_311),
.B1(n_317),
.B2(n_277),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_269),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_310),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_261),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_247),
.C(n_199),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_319),
.C(n_265),
.Y(n_330)
);

OAI22x1_ASAP7_75t_L g307 ( 
.A1(n_265),
.A2(n_198),
.B1(n_167),
.B2(n_169),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_307),
.A2(n_313),
.B1(n_315),
.B2(n_267),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_282),
.A2(n_202),
.B1(n_244),
.B2(n_256),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_223),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_272),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_274),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_260),
.Y(n_316)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_262),
.B(n_199),
.Y(n_318)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_318),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_270),
.B(n_106),
.Y(n_319)
);

NAND2xp33_ASAP7_75t_SL g349 ( 
.A(n_320),
.B(n_324),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_322),
.B(n_327),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_302),
.A2(n_275),
.B1(n_263),
.B2(n_259),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_323),
.A2(n_325),
.B1(n_331),
.B2(n_340),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_302),
.A2(n_263),
.B1(n_268),
.B2(n_278),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_313),
.A2(n_266),
.B1(n_317),
.B2(n_314),
.Y(n_328)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_328),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_305),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_290),
.A2(n_261),
.B1(n_276),
.B2(n_283),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_292),
.A2(n_266),
.B1(n_290),
.B2(n_295),
.Y(n_332)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_332),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_297),
.B(n_261),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_335),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_294),
.B(n_280),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_280),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_342),
.C(n_347),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_301),
.A2(n_279),
.B1(n_273),
.B2(n_285),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_308),
.A2(n_273),
.B1(n_279),
.B2(n_287),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_341),
.A2(n_315),
.B(n_307),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_296),
.B(n_281),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_289),
.Y(n_343)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_343),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_308),
.A2(n_285),
.B1(n_288),
.B2(n_195),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_344),
.A2(n_345),
.B1(n_311),
.B2(n_316),
.Y(n_362)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_298),
.Y(n_346)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_346),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_306),
.B(n_168),
.C(n_106),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_123),
.C(n_141),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_72),
.C(n_71),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_353),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_337),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_354),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_329),
.B(n_293),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_309),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_358),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_338),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_347),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_291),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_361),
.B(n_363),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_312),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_336),
.A2(n_304),
.B1(n_299),
.B2(n_103),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_366),
.A2(n_369),
.B1(n_26),
.B2(n_28),
.Y(n_389)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_340),
.Y(n_367)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_367),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_331),
.Y(n_368)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_368),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_323),
.A2(n_84),
.B1(n_81),
.B2(n_73),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_321),
.B(n_14),
.Y(n_370)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_370),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_374),
.C(n_375),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_326),
.B(n_13),
.Y(n_372)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_372),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_43),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_43),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_355),
.B(n_342),
.C(n_334),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_382),
.C(n_393),
.Y(n_400)
);

NAND3xp33_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_396),
.C(n_0),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_327),
.C(n_348),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_373),
.A2(n_325),
.B1(n_322),
.B2(n_341),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_383),
.A2(n_394),
.B1(n_369),
.B2(n_371),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_366),
.Y(n_385)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_385),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_357),
.B(n_344),
.Y(n_386)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_389),
.A2(n_392),
.B1(n_399),
.B2(n_36),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_356),
.A2(n_43),
.B1(n_29),
.B2(n_27),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_390),
.A2(n_8),
.B1(n_15),
.B2(n_2),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_364),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_29),
.C(n_27),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_373),
.A2(n_29),
.B1(n_27),
.B2(n_18),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_359),
.B(n_17),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_17),
.C(n_28),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_352),
.C(n_374),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_349),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_365),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_401),
.B(n_404),
.Y(n_436)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_384),
.Y(n_402)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_402),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_387),
.A2(n_349),
.B(n_350),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_414),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_376),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_410),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_363),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_380),
.C(n_382),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_388),
.B(n_395),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_408),
.B(n_379),
.Y(n_424)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_397),
.Y(n_411)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_411),
.Y(n_426)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_391),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_415),
.Y(n_432)
);

AOI21x1_ASAP7_75t_L g414 ( 
.A1(n_386),
.A2(n_352),
.B(n_353),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_375),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_416),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_383),
.A2(n_28),
.B1(n_9),
.B2(n_3),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_417),
.A2(n_389),
.B1(n_390),
.B2(n_394),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_385),
.A2(n_7),
.B(n_15),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_418),
.A2(n_419),
.B1(n_36),
.B2(n_9),
.Y(n_433)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_420),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_428),
.Y(n_440)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_424),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_427),
.A2(n_6),
.B1(n_14),
.B2(n_3),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_378),
.C(n_379),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_429),
.Y(n_439)
);

FAx1_ASAP7_75t_SL g429 ( 
.A(n_414),
.B(n_393),
.CI(n_398),
.CON(n_429),
.SN(n_429)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_400),
.B(n_36),
.C(n_1),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_431),
.B(n_434),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_433),
.B(n_435),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_407),
.A2(n_409),
.B1(n_411),
.B2(n_412),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_36),
.C(n_1),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_440),
.B(n_446),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_420),
.Y(n_441)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_441),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_421),
.A2(n_403),
.B(n_402),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_442),
.B(n_444),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_423),
.B(n_415),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_443),
.B(n_445),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_421),
.A2(n_418),
.B1(n_413),
.B2(n_417),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_432),
.B(n_406),
.Y(n_445)
);

NOR3xp33_ASAP7_75t_L g446 ( 
.A(n_425),
.B(n_416),
.C(n_6),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_422),
.B(n_6),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_447),
.A2(n_429),
.B(n_6),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_430),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_439),
.A2(n_426),
.B(n_431),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_451),
.A2(n_454),
.B(n_458),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_440),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_457),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_448),
.A2(n_434),
.B(n_436),
.Y(n_454)
);

A2O1A1Ixp33_ASAP7_75t_L g458 ( 
.A1(n_441),
.A2(n_429),
.B(n_435),
.C(n_436),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_450),
.B(n_430),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_460),
.B(n_461),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_459),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_464),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_455),
.B(n_437),
.C(n_442),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_465),
.B(n_468),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_456),
.A2(n_444),
.B(n_438),
.Y(n_466)
);

A2O1A1O1Ixp25_ASAP7_75t_L g474 ( 
.A1(n_466),
.A2(n_4),
.B(n_10),
.C(n_13),
.D(n_14),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_456),
.B(n_5),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_15),
.C(n_5),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_469),
.B(n_0),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_472),
.C(n_474),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_462),
.A2(n_3),
.B(n_4),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_470),
.B(n_463),
.C(n_464),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_476),
.B(n_473),
.Y(n_477)
);

OAI221xp5_ASAP7_75t_L g478 ( 
.A1(n_477),
.A2(n_467),
.B1(n_475),
.B2(n_10),
.C(n_1),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_478),
.B(n_10),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_479),
.B(n_10),
.Y(n_480)
);


endmodule