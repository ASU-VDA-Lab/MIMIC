module fake_jpeg_20418_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_60),
.Y(n_65)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_59),
.B(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_74),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_52),
.B1(n_48),
.B2(n_42),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_68),
.B1(n_71),
.B2(n_50),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_52),
.B1(n_41),
.B2(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_4),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_45),
.B1(n_51),
.B2(n_43),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_25),
.B1(n_30),
.B2(n_29),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_50),
.B1(n_49),
.B2(n_51),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_80),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_74),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_85),
.Y(n_98)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_89),
.B1(n_5),
.B2(n_6),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_88),
.B1(n_6),
.B2(n_7),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_1),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_69),
.B(n_20),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_5),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_87),
.B1(n_83),
.B2(n_10),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_21),
.B1(n_38),
.B2(n_36),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_84),
.B1(n_95),
.B2(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_99),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_102),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_98),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_104),
.B(n_105),
.Y(n_106)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

AOI221xp5_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_97),
.B1(n_98),
.B2(n_90),
.C(n_83),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_103),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_110),
.A3(n_108),
.B1(n_9),
.B2(n_8),
.C1(n_15),
.C2(n_16),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_105),
.B1(n_97),
.B2(n_10),
.Y(n_110)
);

AOI31xp67_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_109),
.A3(n_18),
.B(n_26),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_13),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_28),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_31),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_32),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_34),
.Y(n_118)
);


endmodule