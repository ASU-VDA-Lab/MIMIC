module fake_netlist_1_7583_n_32 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_32);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_7;
wire n_27;
BUFx3_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
BUFx10_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
CKINVDCx20_ASAP7_75t_R g9 ( .A(n_6), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_1), .Y(n_10) );
AND2x6_ASAP7_75t_L g11 ( .A(n_3), .B(n_2), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_9), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_10), .B(n_0), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_12), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_7), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
INVx4_ASAP7_75t_SL g18 ( .A(n_15), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_13), .B(n_8), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_18), .B(n_14), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
AOI221xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_19), .B1(n_13), .B2(n_22), .C(n_21), .Y(n_25) );
NOR2xp33_ASAP7_75t_R g26 ( .A(n_23), .B(n_11), .Y(n_26) );
CKINVDCx16_ASAP7_75t_R g27 ( .A(n_26), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_8), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_25), .B(n_11), .Y(n_29) );
HB1xp67_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
AOI22xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_29), .B1(n_30), .B2(n_11), .Y(n_32) );
endmodule