module fake_jpeg_23023_n_48 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_7),
.A2(n_0),
.B(n_3),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_8),
.A2(n_14),
.B1(n_15),
.B2(n_11),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_17),
.A2(n_10),
.B1(n_9),
.B2(n_12),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_7),
.B(n_6),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_18),
.B(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_22),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_23),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_5),
.C(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_17),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_21),
.Y(n_33)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_33),
.C(n_26),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_41),
.C(n_29),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_40),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_30),
.C(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_28),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_28),
.C(n_42),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_10),
.C(n_12),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_13),
.B(n_32),
.C(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_47),
.B(n_13),
.Y(n_48)
);


endmodule