module fake_jpeg_17560_n_159 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_159);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_37),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_36),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_SL g37 ( 
.A1(n_14),
.A2(n_6),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_44),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_10),
.B1(n_26),
.B2(n_16),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_45),
.B1(n_18),
.B2(n_23),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_14),
.A2(n_20),
.B1(n_24),
.B2(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_47),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_23),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_18),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_47),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_31),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_73),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_70),
.B1(n_55),
.B2(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_75),
.Y(n_88)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_37),
.B(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_81),
.Y(n_92)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_81),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_93),
.Y(n_113)
);

OR2x4_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_56),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_92),
.B(n_87),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_95),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_65),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_100),
.C(n_102),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_101),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_57),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_59),
.B(n_74),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_71),
.B1(n_76),
.B2(n_73),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_58),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_105),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_58),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g107 ( 
.A(n_94),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

XOR2x2_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_69),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_117),
.C(n_118),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_71),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_113),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_98),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_117),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_83),
.B(n_98),
.C(n_100),
.D(n_113),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_127),
.A2(n_112),
.B(n_107),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_131),
.Y(n_133)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_136),
.B1(n_139),
.B2(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_127),
.B(n_110),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_138),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_110),
.B(n_103),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_140),
.B(n_128),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_126),
.A2(n_107),
.B1(n_116),
.B2(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_139),
.B(n_128),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_131),
.B1(n_121),
.B2(n_120),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_137),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_134),
.C(n_133),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_145),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_147),
.B(n_143),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_133),
.C(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_152),
.Y(n_155)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_148),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_141),
.C(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_153),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_150),
.B1(n_155),
.B2(n_157),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_158),
.Y(n_159)
);


endmodule