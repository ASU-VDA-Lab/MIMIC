module fake_jpeg_21237_n_225 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx11_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_40),
.Y(n_42)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_47),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_22),
.B1(n_25),
.B2(n_16),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_45),
.A2(n_34),
.B1(n_35),
.B2(n_17),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_29),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_25),
.B1(n_22),
.B2(n_17),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_34),
.B1(n_39),
.B2(n_25),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_16),
.B1(n_23),
.B2(n_26),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_26),
.B1(n_21),
.B2(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_53),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_20),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_49),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_64),
.Y(n_108)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_65),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_28),
.B(n_18),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_67),
.B1(n_75),
.B2(n_78),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_27),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_34),
.B1(n_39),
.B2(n_22),
.Y(n_67)
);

BUFx24_ASAP7_75t_SL g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_82),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_58),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_19),
.C(n_37),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_41),
.C(n_38),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_33),
.Y(n_109)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_34),
.B1(n_39),
.B2(n_23),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_77),
.B(n_81),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_42),
.B1(n_46),
.B2(n_44),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_43),
.B(n_23),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_46),
.B(n_24),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_85),
.Y(n_105)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_90),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_34),
.B1(n_39),
.B2(n_35),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_35),
.B1(n_18),
.B2(n_32),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_89),
.B1(n_33),
.B2(n_32),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_35),
.B1(n_41),
.B2(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_0),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_100),
.B1(n_102),
.B2(n_107),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_38),
.B1(n_37),
.B2(n_32),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_19),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_109),
.B(n_112),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_62),
.B1(n_76),
.B2(n_78),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_72),
.B1(n_83),
.B2(n_80),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_38),
.B1(n_37),
.B2(n_18),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_33),
.B(n_1),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_87),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_70),
.B(n_74),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_86),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_63),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_96),
.B(n_95),
.C(n_97),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_108),
.B(n_85),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_120),
.B(n_123),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_126),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_90),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_125),
.C(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_60),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_101),
.C(n_93),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_127),
.A2(n_130),
.B(n_6),
.Y(n_158)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_0),
.B1(n_6),
.B2(n_7),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_79),
.B1(n_38),
.B2(n_3),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_138),
.B1(n_97),
.B2(n_5),
.Y(n_151)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_84),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_94),
.B(n_15),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_137),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_138)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_146),
.C(n_150),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_104),
.B(n_112),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_158),
.B(n_159),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_100),
.C(n_107),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_149),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_99),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_103),
.C(n_84),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_157),
.B1(n_132),
.B2(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_154),
.B(n_138),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_31),
.B(n_7),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_155),
.A2(n_127),
.B(n_132),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_9),
.B(n_10),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_163),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_164),
.B1(n_169),
.B2(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_131),
.B(n_124),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_170),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_124),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_136),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_157),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_133),
.C(n_137),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_146),
.C(n_149),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_148),
.B1(n_151),
.B2(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_182),
.C(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_142),
.C(n_141),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_142),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_190),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_145),
.B1(n_154),
.B2(n_158),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_187),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_145),
.B1(n_159),
.B2(n_155),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_168),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_172),
.B(n_161),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_186),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_189),
.A2(n_168),
.B1(n_167),
.B2(n_164),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_165),
.B1(n_182),
.B2(n_171),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_197),
.C(n_134),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_162),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_163),
.C(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_152),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_185),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_203),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_188),
.B(n_183),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_205),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_128),
.B(n_152),
.C(n_139),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_195),
.A3(n_152),
.B1(n_197),
.B2(n_194),
.C1(n_200),
.C2(n_9),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_207),
.B(n_208),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_201),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_212),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_202),
.B(n_198),
.Y(n_212)
);

OAI21x1_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_11),
.B(n_13),
.Y(n_218)
);

OAI21x1_ASAP7_75t_L g216 ( 
.A1(n_214),
.A2(n_206),
.B(n_200),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_218),
.B(n_213),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_206),
.B(n_12),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_13),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_221),
.C(n_14),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_210),
.C(n_14),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_222),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_223),
.Y(n_225)
);


endmodule