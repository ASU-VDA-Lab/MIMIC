module real_jpeg_5563_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_1),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_2),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_2),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_2),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_2),
.B(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_2),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_2),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_2),
.B(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_3),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_3),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_3),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_3),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_4),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_4),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_4),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_4),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_4),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_4),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_4),
.B(n_465),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_5),
.B(n_91),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_5),
.A2(n_116),
.B(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_5),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_5),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_5),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_5),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_5),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_5),
.B(n_368),
.Y(n_395)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_7),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_7),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_7),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g368 ( 
.A(n_7),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_8),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_8),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_8),
.B(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_8),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_8),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_8),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_8),
.B(n_467),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_9),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_9),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_9),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_9),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_9),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_9),
.B(n_357),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_9),
.B(n_392),
.Y(n_391)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_10),
.Y(n_117)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_10),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g299 ( 
.A(n_10),
.Y(n_299)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_12),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_12),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_12),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_12),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_12),
.B(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_12),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_12),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_12),
.B(n_409),
.Y(n_408)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_13),
.Y(n_122)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_13),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_13),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_14),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_14),
.Y(n_357)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_14),
.Y(n_412)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_15),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_15),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_15),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_15),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_15),
.B(n_86),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_15),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_447),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_203),
.B(n_445),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_170),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_20),
.B(n_170),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_98),
.C(n_126),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_21),
.B(n_98),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_60),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_42),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_23),
.B(n_42),
.C(n_60),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.C(n_40),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_24),
.B(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.C(n_32),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_52),
.C(n_56),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_25),
.A2(n_56),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_25),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_25),
.A2(n_32),
.B1(n_94),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_25),
.A2(n_94),
.B1(n_370),
.B2(n_372),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_25),
.B(n_372),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_27),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_27),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_27),
.A2(n_129),
.B1(n_198),
.B2(n_202),
.Y(n_197)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_31),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_31),
.Y(n_228)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_31),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_32),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_32),
.B(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_32),
.A2(n_132),
.B1(n_264),
.B2(n_265),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_33),
.Y(n_364)
);

INVx8_ASAP7_75t_L g386 ( 
.A(n_33),
.Y(n_386)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_34),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_35),
.A2(n_40),
.B1(n_50),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_35),
.Y(n_169)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_39),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_44),
.B1(n_45),
.B2(n_50),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_51),
.B1(n_58),
.B2(n_59),
.Y(n_42)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_45),
.B(n_50),
.C(n_59),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_48),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_48),
.Y(n_218)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_49),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_49),
.Y(n_311)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_52),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_52),
.B(n_226),
.C(n_229),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_52),
.A2(n_96),
.B1(n_226),
.B2(n_294),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_80),
.C(n_92),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_61),
.B(n_80),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_67),
.B2(n_68),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_70),
.C(n_75),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_62),
.A2(n_63),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_62),
.B(n_121),
.C(n_125),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_62),
.A2(n_63),
.B1(n_147),
.B2(n_148),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_63),
.B(n_148),
.Y(n_302)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_75),
.B2(n_79),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_72),
.Y(n_161)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_73),
.Y(n_330)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_74),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_74),
.Y(n_354)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_75),
.A2(n_79),
.B1(n_459),
.B2(n_460),
.Y(n_458)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.C(n_88),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_85),
.B(n_88),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_87),
.Y(n_242)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_92),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_118),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_100),
.B(n_101),
.C(n_118),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_112),
.B2(n_113),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_106),
.B1(n_110),
.B2(n_111),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_106),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_106),
.B(n_110),
.C(n_113),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_106),
.B(n_135),
.Y(n_212)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_134),
.C(n_139),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_117),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_124),
.B2(n_125),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_121),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_124),
.A2(n_125),
.B1(n_182),
.B2(n_185),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_124),
.B(n_256),
.C(n_260),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_124),
.A2(n_125),
.B1(n_260),
.B2(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_125),
.B(n_178),
.C(n_182),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_126),
.B(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_145),
.C(n_167),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_127),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.C(n_143),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_128),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_129),
.B(n_193),
.C(n_198),
.Y(n_457)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_133),
.B(n_143),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_139),
.B(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_145),
.B(n_167),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_160),
.C(n_162),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_146),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.C(n_159),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_147),
.A2(n_148),
.B1(n_159),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_152),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_153),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_153),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_153),
.A2(n_177),
.B1(n_178),
.B2(n_269),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_158),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_159),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_160),
.A2(n_162),
.B1(n_163),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_166),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g471 ( 
.A(n_170),
.Y(n_471)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.CI(n_186),
.CON(n_170),
.SN(n_170)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_171),
.B(n_172),
.C(n_186),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_174),
.B(n_175),
.C(n_176),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_214),
.C(n_219),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_177),
.A2(n_178),
.B1(n_214),
.B2(n_215),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_182),
.Y(n_185)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_184),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_187),
.B(n_189),
.C(n_192),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_195),
.Y(n_465)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AOI221xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_343),
.B1(n_438),
.B2(n_443),
.C(n_444),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_282),
.C(n_286),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_206),
.A2(n_439),
.B(n_442),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_275),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_207),
.B(n_275),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_248),
.C(n_251),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_208),
.B(n_248),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_233),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_209),
.B(n_234),
.C(n_245),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.C(n_224),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_211),
.B(n_225),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_213),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_219),
.B(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g371 ( 
.A(n_223),
.Y(n_371)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_226),
.Y(n_294)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_229),
.B(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_245),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_240),
.C(n_243),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_274),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_235),
.A2(n_236),
.B(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_243),
.Y(n_274)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_242),
.B(n_297),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_251),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_268),
.C(n_273),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.C(n_262),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_253),
.B(n_339),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_255),
.A2(n_262),
.B1(n_263),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_255),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_256),
.B(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_260),
.Y(n_323)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_273),
.Y(n_290)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_279),
.C(n_281),
.Y(n_283)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_282),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_283),
.B(n_284),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_316),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_287),
.A2(n_440),
.B(n_441),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_314),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_288),
.B(n_314),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.C(n_312),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_289),
.B(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_291),
.B(n_312),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.C(n_300),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_295),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.C(n_306),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_301),
.A2(n_302),
.B1(n_426),
.B2(n_427),
.Y(n_425)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_303),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_311),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_341),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_317),
.B(n_341),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.C(n_338),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_318),
.B(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_320),
.B(n_338),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.C(n_336),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_321),
.B(n_429),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_324),
.A2(n_336),
.B1(n_337),
.B2(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_324),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_328),
.C(n_331),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_325),
.A2(n_326),
.B1(n_331),
.B2(n_332),
.Y(n_418)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_328),
.B(n_418),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_330),
.Y(n_379)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_433),
.B(n_437),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_420),
.B(n_432),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_404),
.B(n_419),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_380),
.B(n_403),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_373),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_348),
.B(n_373),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_360),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_349),
.B(n_361),
.C(n_369),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_355),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_350),
.B(n_356),
.C(n_358),
.Y(n_416)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_369),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_365),
.Y(n_374)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_370),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.C(n_376),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_375),
.A2(n_376),
.B1(n_377),
.B2(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_375),
.Y(n_401)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_397),
.B(n_402),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_390),
.B(n_396),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_389),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_389),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_387),
.Y(n_398)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_395),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_399),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_406),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_415),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_407),
.A2(n_423),
.B1(n_424),
.B2(n_425),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_407),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_416),
.C(n_417),
.Y(n_431)
);

FAx1_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_413),
.CI(n_414),
.CON(n_407),
.SN(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_431),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_431),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_428),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_423),
.B(n_425),
.C(n_428),
.Y(n_434)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_426),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_434),
.B(n_435),
.Y(n_437)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_470),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_450),
.B(n_451),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_461),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_464),
.A2(n_466),
.B1(n_468),
.B2(n_469),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_464),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_466),
.Y(n_469)
);


endmodule